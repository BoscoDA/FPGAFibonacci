-- Copyright (C) 2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, the Intel Quartus Prime License Agreement, the Intel
-- MegaCore Function License Agreement, or other applicable 
-- license agreement, including, without limitation, that your
-- use is for the sole purpose of simulating designs for use 
-- exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- Quartus Prime 17.0.1 Build 598 06/07/2017
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_atx_pll	is
	generic (
		-- Entity parameters
		analog_mode	:	string	:=	"user_custom";
		bandwidth_range_high	:	string	:=	"0 hz";
		bandwidth_range_low	:	string	:=	"0 hz";
		bonding	:	string	:=	"pll_bonding";
		bw_sel	:	string	:=	"low";
		cal_status	:	string	:=	"cal_done";
		calibration_mode	:	string	:=	"cal_off";
		cascadeclk_test	:	string	:=	"cascadetest_off";
		cgb_div	:	integer	:=	1;
		clk_high_perf_voltage	:	bit_vector	:=	B"000000000000";
		clk_low_power_voltage	:	bit_vector	:=	B"000000000000";
		clk_mid_power_voltage	:	bit_vector	:=	B"000000000000";
		cp_compensation_enable	:	string	:=	"true";
		cp_current_setting	:	string	:=	"cp_current_setting0";
		cp_lf_3rd_pole_freq	:	string	:=	"lf_3rd_pole_setting0";
		cp_lf_order	:	string	:=	"lf_2nd_order";
		cp_testmode	:	string	:=	"cp_normal";
		d2a_voltage	:	string	:=	"d2a_disable";
		datarate	:	string	:=	"0 bps";
		device_variant	:	string	:=	"device1";
		dprio_clk_vreg_boost_expected_voltage	:	bit_vector	:=	B"000000000000";
		dprio_clk_vreg_boost_scratch	:	bit_vector	:=	B"000";
		dprio_clk_vreg_boost_step_size	:	bit_vector	:=	B"00000";
		dprio_lc_vreg1_boost_expected_voltage	:	bit_vector	:=	B"000000000000";
		dprio_lc_vreg1_boost_scratch	:	bit_vector	:=	B"000";
		dprio_lc_vreg_boost_expected_voltage	:	bit_vector	:=	B"000000000000";
		dprio_lc_vreg_boost_scratch	:	bit_vector	:=	B"000";
		dprio_mcgb_vreg_boost_expected_voltage	:	bit_vector	:=	B"000000000000";
		dprio_mcgb_vreg_boost_scratch	:	bit_vector	:=	B"000";
		dprio_mcgb_vreg_boost_step_size	:	bit_vector	:=	B"00000";
		dprio_vreg1_boost_step_size	:	bit_vector	:=	B"00000";
		dprio_vreg_boost_step_size	:	bit_vector	:=	B"00000";
		dsm_ecn_bypass	:	string	:=	"false";
		dsm_ecn_test_en	:	string	:=	"false";
		dsm_fractional_division	:	string	:=	"00000000000000000000000000000000";
		dsm_fractional_value_ready	:	string	:=	"pll_k_ready";
		dsm_mode	:	string	:=	"dsm_mode_integer";
		dsm_out_sel	:	string	:=	"pll_dsm_disable";
		enable_hclk	:	string	:=	"hclk_disabled";
		enable_idle_atx_pll_support	:	string	:=	"idle_none";
		enable_lc_calibration	:	string	:=	"false";
		enable_lc_vreg_calibration	:	string	:=	"false";
		expected_lc_boost_voltage	:	bit_vector	:=	B"000000000000";
		f_max_lcnt_fpll_cascading	:	string	:=	"000000000000000000000000000000000001";
		f_max_pfd	:	string	:=	"0 hz";
		f_max_pfd_fractional	:	string	:=	"0 hz";
		f_max_ref	:	string	:=	"0 hz";
		f_max_tank_0	:	string	:=	"0 hz";
		f_max_tank_1	:	string	:=	"0 hz";
		f_max_tank_2	:	string	:=	"0 hz";
		f_max_vco	:	string	:=	"0 hz";
		f_max_vco_fractional	:	string	:=	"0 hz";
		f_max_x1	:	string	:=	"0 hz";
		f_min_pfd	:	string	:=	"0 hz";
		f_min_ref	:	string	:=	"0 hz";
		f_min_tank_0	:	string	:=	"0 hz";
		f_min_tank_1	:	string	:=	"0 hz";
		f_min_tank_2	:	string	:=	"0 hz";
		f_min_vco	:	string	:=	"0 hz";
		fb_select	:	string	:=	"direct_fb";
		fpll_refclk_selection	:	string	:=	"select_div_by_2";
		hclk_divide	:	integer	:=	1;
		initial_settings	:	string	:=	"false";
		iqclk_mux_sel	:	string	:=	"power_down";
		is_cascaded_pll	:	string	:=	"false";
		is_otn	:	string	:=	"false";
		is_sdi	:	string	:=	"false";
		l_counter	:	integer	:=	1;
		l_counter_enable	:	string	:=	"false";
		l_counter_scratch	:	bit_vector	:=	B"00001";
		lc_atb	:	string	:=	"atb_selectdisable";
		lc_mode	:	string	:=	"lccmu_pd";
		lc_to_fpll_l_counter	:	string	:=	"lcounter_setting0";
		lc_to_fpll_l_counter_scratch	:	bit_vector	:=	B"00001";
		lf_cbig_size	:	string	:=	"lf_cbig_setting0";
		lf_resistance	:	string	:=	"lf_setting0";
		lf_ripplecap	:	string	:=	"lf_ripple_cap_0";
		m_counter	:	integer	:=	8;
		max_fractional_percentage	:	bit_vector	:=	B"0000000";
		min_fractional_percentage	:	bit_vector	:=	B"0000000";
		n_counter_scratch	:	bit_vector	:=	B"0001";
		output_clock_frequency	:	string	:=	"0 hz";
		output_regulator_supply	:	string	:=	"vreg1v_setting3";
		overrange_voltage	:	string	:=	"over_setting5";
		pfd_delay_compensation	:	string	:=	"normal_delay";
		pfd_pulse_width	:	string	:=	"pulse_width_setting0";
		pm_speed_grade	:	string	:=	"e2";
		pma_width	:	integer	:=	8;
		power_mode	:	string	:=	"low_power";
		power_rail_et	:	integer	:=	0;
		powerdown_mode	:	string	:=	"powerup";
		primary_use	:	string	:=	"hssi_x1";
		prot_mode	:	string	:=	"basic_tx";
		ref_clk_div	:	integer	:=	1;
		reference_clock_frequency	:	string	:=	"0 hz";
		regulator_bypass	:	string	:=	"reg_enable";
		side	:	string	:=	"side_unknown";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode";
		tank_band	:	string	:=	"lc_band0";
		tank_sel	:	string	:=	"lctank0";
		tank_voltage_coarse	:	string	:=	"vreg_setting_coarse0";
		tank_voltage_fine	:	string	:=	"vreg_setting5";
		top_or_bottom	:	string	:=	"tb_unknown";
		underrange_voltage	:	string	:=	"under_setting4";
		vccdreg_clk	:	string	:=	"vreg_clk0";
		vccdreg_fb	:	string	:=	"vreg_fb0";
		vccdreg_fw	:	string	:=	"vreg_fw0";
		vco_bypass_enable	:	string	:=	"false";
		vco_freq	:	string	:=	"0 hz";
		xcpvco_xchgpmplf_cp_current_boost	:	string	:=	"normal_setting"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		core_clk	:	in	std_logic	:=	'0';
		iqtxrxclk	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		lf_rst_n	:	in	std_logic	:=	'0';
		refclk	:	in	std_logic	:=	'0';
		rst_n	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		clk0_16g	:	out	std_logic	:=	'0';
		clk0_8g	:	out	std_logic	:=	'0';
		clk180_16g	:	out	std_logic	:=	'0';
		clk180_8g	:	out	std_logic	:=	'0';
		clklow_buf	:	out	std_logic	:=	'0';
		fref_buf	:	out	std_logic	:=	'0';
		hclk_out	:	out	std_logic	:=	'0';
		iqtxrxclk_out	:	out	std_logic	:=	'0';
		lc_to_fpll_refclk	:	out	std_logic	:=	'0';
		lock	:	out	std_logic	:=	'0';
		m_cnt_int	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		overrange	:	out	std_logic	:=	'0';
		underrange	:	out	std_logic	:=	'0'
	);
end twentynm_atx_pll;

architecture behavior of twentynm_atx_pll	is

constant clk_high_perf_voltage_int	:	integer	:=	bin2int(clk_high_perf_voltage);
constant clk_low_power_voltage_int	:	integer	:=	bin2int(clk_low_power_voltage);
constant clk_mid_power_voltage_int	:	integer	:=	bin2int(clk_mid_power_voltage);
constant dprio_clk_vreg_boost_expected_voltage_int	:	integer	:=	bin2int(dprio_clk_vreg_boost_expected_voltage);
constant dprio_clk_vreg_boost_scratch_int	:	integer	:=	bin2int(dprio_clk_vreg_boost_scratch);
constant dprio_clk_vreg_boost_step_size_int	:	integer	:=	bin2int(dprio_clk_vreg_boost_step_size);
constant dprio_lc_vreg1_boost_expected_voltage_int	:	integer	:=	bin2int(dprio_lc_vreg1_boost_expected_voltage);
constant dprio_lc_vreg1_boost_scratch_int	:	integer	:=	bin2int(dprio_lc_vreg1_boost_scratch);
constant dprio_lc_vreg_boost_expected_voltage_int	:	integer	:=	bin2int(dprio_lc_vreg_boost_expected_voltage);
constant dprio_lc_vreg_boost_scratch_int	:	integer	:=	bin2int(dprio_lc_vreg_boost_scratch);
constant dprio_mcgb_vreg_boost_expected_voltage_int	:	integer	:=	bin2int(dprio_mcgb_vreg_boost_expected_voltage);
constant dprio_mcgb_vreg_boost_scratch_int	:	integer	:=	bin2int(dprio_mcgb_vreg_boost_scratch);
constant dprio_mcgb_vreg_boost_step_size_int	:	integer	:=	bin2int(dprio_mcgb_vreg_boost_step_size);
constant dprio_vreg1_boost_step_size_int	:	integer	:=	bin2int(dprio_vreg1_boost_step_size);
constant dprio_vreg_boost_step_size_int	:	integer	:=	bin2int(dprio_vreg_boost_step_size);
constant expected_lc_boost_voltage_int	:	integer	:=	bin2int(expected_lc_boost_voltage);
constant l_counter_scratch_int	:	integer	:=	bin2int(l_counter_scratch);
constant lc_to_fpll_l_counter_scratch_int	:	integer	:=	bin2int(lc_to_fpll_l_counter_scratch);
constant max_fractional_percentage_int	:	integer	:=	bin2int(max_fractional_percentage);
constant min_fractional_percentage_int	:	integer	:=	bin2int(min_fractional_percentage);
constant n_counter_scratch_int	:	integer	:=	bin2int(n_counter_scratch);



component	twentynm_atx_pll_encrypted
	generic (
		-- Architecture parameters
		analog_mode	:	string	:=	"user_custom";
		bandwidth_range_high	:	string	:=	"0 hz";
		bandwidth_range_low	:	string	:=	"0 hz";
		bonding	:	string	:=	"pll_bonding";
		bw_sel	:	string	:=	"low";
		cal_status	:	string	:=	"cal_done";
		calibration_mode	:	string	:=	"cal_off";
		cascadeclk_test	:	string	:=	"cascadetest_off";
		cgb_div	:	integer	:=	1;
		clk_high_perf_voltage	:	integer	:=	0;
		clk_low_power_voltage	:	integer	:=	0;
		clk_mid_power_voltage	:	integer	:=	0;
		cp_compensation_enable	:	string	:=	"true";
		cp_current_setting	:	string	:=	"cp_current_setting0";
		cp_lf_3rd_pole_freq	:	string	:=	"lf_3rd_pole_setting0";
		cp_lf_order	:	string	:=	"lf_2nd_order";
		cp_testmode	:	string	:=	"cp_normal";
		d2a_voltage	:	string	:=	"d2a_disable";
		datarate	:	string	:=	"0 bps";
		device_variant	:	string	:=	"device1";
		dprio_clk_vreg_boost_expected_voltage	:	integer	:=	0;
		dprio_clk_vreg_boost_scratch	:	integer	:=	0;
		dprio_clk_vreg_boost_step_size	:	integer	:=	0;
		dprio_lc_vreg1_boost_expected_voltage	:	integer	:=	0;
		dprio_lc_vreg1_boost_scratch	:	integer	:=	0;
		dprio_lc_vreg_boost_expected_voltage	:	integer	:=	0;
		dprio_lc_vreg_boost_scratch	:	integer	:=	0;
		dprio_mcgb_vreg_boost_expected_voltage	:	integer	:=	0;
		dprio_mcgb_vreg_boost_scratch	:	integer	:=	0;
		dprio_mcgb_vreg_boost_step_size	:	integer	:=	0;
		dprio_vreg1_boost_step_size	:	integer	:=	0;
		dprio_vreg_boost_step_size	:	integer	:=	0;
		dsm_ecn_bypass	:	string	:=	"false";
		dsm_ecn_test_en	:	string	:=	"false";
		dsm_fractional_division	:	string	:=	"00000000000000000000000000000000";
		dsm_fractional_value_ready	:	string	:=	"pll_k_ready";
		dsm_mode	:	string	:=	"dsm_mode_integer";
		dsm_out_sel	:	string	:=	"pll_dsm_disable";
		enable_hclk	:	string	:=	"hclk_disabled";
		enable_idle_atx_pll_support	:	string	:=	"idle_none";
		enable_lc_calibration	:	string	:=	"false";
		enable_lc_vreg_calibration	:	string	:=	"false";
		expected_lc_boost_voltage	:	integer	:=	0;
		f_max_lcnt_fpll_cascading	:	string	:=	"000000000000000000000000000000000001";
		f_max_pfd	:	string	:=	"0 hz";
		f_max_pfd_fractional	:	string	:=	"0 hz";
		f_max_ref	:	string	:=	"0 hz";
		f_max_tank_0	:	string	:=	"0 hz";
		f_max_tank_1	:	string	:=	"0 hz";
		f_max_tank_2	:	string	:=	"0 hz";
		f_max_vco	:	string	:=	"0 hz";
		f_max_vco_fractional	:	string	:=	"0 hz";
		f_max_x1	:	string	:=	"0 hz";
		f_min_pfd	:	string	:=	"0 hz";
		f_min_ref	:	string	:=	"0 hz";
		f_min_tank_0	:	string	:=	"0 hz";
		f_min_tank_1	:	string	:=	"0 hz";
		f_min_tank_2	:	string	:=	"0 hz";
		f_min_vco	:	string	:=	"0 hz";
		fb_select	:	string	:=	"direct_fb";
		fpll_refclk_selection	:	string	:=	"select_div_by_2";
		hclk_divide	:	integer	:=	1;
		initial_settings	:	string	:=	"false";
		iqclk_mux_sel	:	string	:=	"power_down";
		is_cascaded_pll	:	string	:=	"false";
		is_otn	:	string	:=	"false";
		is_sdi	:	string	:=	"false";
		l_counter	:	integer	:=	1;
		l_counter_enable	:	string	:=	"false";
		l_counter_scratch	:	integer	:=	1;
		lc_atb	:	string	:=	"atb_selectdisable";
		lc_mode	:	string	:=	"lccmu_pd";
		lc_to_fpll_l_counter	:	string	:=	"lcounter_setting0";
		lc_to_fpll_l_counter_scratch	:	integer	:=	1;
		lf_cbig_size	:	string	:=	"lf_cbig_setting0";
		lf_resistance	:	string	:=	"lf_setting0";
		lf_ripplecap	:	string	:=	"lf_ripple_cap_0";
		m_counter	:	integer	:=	8;
		max_fractional_percentage	:	integer	:=	0;
		min_fractional_percentage	:	integer	:=	0;
		n_counter_scratch	:	integer	:=	1;
		output_clock_frequency	:	string	:=	"0 hz";
		output_regulator_supply	:	string	:=	"vreg1v_setting3";
		overrange_voltage	:	string	:=	"over_setting5";
		pfd_delay_compensation	:	string	:=	"normal_delay";
		pfd_pulse_width	:	string	:=	"pulse_width_setting0";
		pm_speed_grade	:	string	:=	"e2";
		pma_width	:	integer	:=	8;
		power_mode	:	string	:=	"low_power";
		power_rail_et	:	integer	:=	0;
		powerdown_mode	:	string	:=	"powerup";
		primary_use	:	string	:=	"hssi_x1";
		prot_mode	:	string	:=	"basic_tx";
		ref_clk_div	:	integer	:=	1;
		reference_clock_frequency	:	string	:=	"0 hz";
		regulator_bypass	:	string	:=	"reg_enable";
		side	:	string	:=	"side_unknown";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode";
		tank_band	:	string	:=	"lc_band0";
		tank_sel	:	string	:=	"lctank0";
		tank_voltage_coarse	:	string	:=	"vreg_setting_coarse0";
		tank_voltage_fine	:	string	:=	"vreg_setting5";
		top_or_bottom	:	string	:=	"tb_unknown";
		underrange_voltage	:	string	:=	"under_setting4";
		vccdreg_clk	:	string	:=	"vreg_clk0";
		vccdreg_fb	:	string	:=	"vreg_fb0";
		vccdreg_fw	:	string	:=	"vreg_fw0";
		vco_bypass_enable	:	string	:=	"false";
		vco_freq	:	string	:=	"0 hz";
		xcpvco_xchgpmplf_cp_current_boost	:	string	:=	"normal_setting"
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		core_clk	:	in	std_logic	:=	'0';
		iqtxrxclk	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		lf_rst_n	:	in	std_logic	:=	'0';
		refclk	:	in	std_logic	:=	'0';
		rst_n	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		clk0_16g	:	out	std_logic	:=	'0';
		clk0_8g	:	out	std_logic	:=	'0';
		clk180_16g	:	out	std_logic	:=	'0';
		clk180_8g	:	out	std_logic	:=	'0';
		clklow_buf	:	out	std_logic	:=	'0';
		fref_buf	:	out	std_logic	:=	'0';
		hclk_out	:	out	std_logic	:=	'0';
		iqtxrxclk_out	:	out	std_logic	:=	'0';
		lc_to_fpll_refclk	:	out	std_logic	:=	'0';
		lock	:	out	std_logic	:=	'0';
		m_cnt_int	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		overrange	:	out	std_logic	:=	'0';
		underrange	:	out	std_logic	:=	'0'
	);
end component;

begin



inst : twentynm_atx_pll_encrypted
	generic map (
		-- Instance parameters
		analog_mode	=>	analog_mode,
		bandwidth_range_high	=>	bandwidth_range_high,
		bandwidth_range_low	=>	bandwidth_range_low,
		bonding	=>	bonding,
		bw_sel	=>	bw_sel,
		cal_status	=>	cal_status,
		calibration_mode	=>	calibration_mode,
		cascadeclk_test	=>	cascadeclk_test,
		cgb_div	=>	cgb_div,
		clk_high_perf_voltage	=>	clk_high_perf_voltage_int,
		clk_low_power_voltage	=>	clk_low_power_voltage_int,
		clk_mid_power_voltage	=>	clk_mid_power_voltage_int,
		cp_compensation_enable	=>	cp_compensation_enable,
		cp_current_setting	=>	cp_current_setting,
		cp_lf_3rd_pole_freq	=>	cp_lf_3rd_pole_freq,
		cp_lf_order	=>	cp_lf_order,
		cp_testmode	=>	cp_testmode,
		d2a_voltage	=>	d2a_voltage,
		datarate	=>	datarate,
		device_variant	=>	device_variant,
		dprio_clk_vreg_boost_expected_voltage	=>	dprio_clk_vreg_boost_expected_voltage_int,
		dprio_clk_vreg_boost_scratch	=>	dprio_clk_vreg_boost_scratch_int,
		dprio_clk_vreg_boost_step_size	=>	dprio_clk_vreg_boost_step_size_int,
		dprio_lc_vreg1_boost_expected_voltage	=>	dprio_lc_vreg1_boost_expected_voltage_int,
		dprio_lc_vreg1_boost_scratch	=>	dprio_lc_vreg1_boost_scratch_int,
		dprio_lc_vreg_boost_expected_voltage	=>	dprio_lc_vreg_boost_expected_voltage_int,
		dprio_lc_vreg_boost_scratch	=>	dprio_lc_vreg_boost_scratch_int,
		dprio_mcgb_vreg_boost_expected_voltage	=>	dprio_mcgb_vreg_boost_expected_voltage_int,
		dprio_mcgb_vreg_boost_scratch	=>	dprio_mcgb_vreg_boost_scratch_int,
		dprio_mcgb_vreg_boost_step_size	=>	dprio_mcgb_vreg_boost_step_size_int,
		dprio_vreg1_boost_step_size	=>	dprio_vreg1_boost_step_size_int,
		dprio_vreg_boost_step_size	=>	dprio_vreg_boost_step_size_int,
		dsm_ecn_bypass	=>	dsm_ecn_bypass,
		dsm_ecn_test_en	=>	dsm_ecn_test_en,
		dsm_fractional_division	=>	dsm_fractional_division,
		dsm_fractional_value_ready	=>	dsm_fractional_value_ready,
		dsm_mode	=>	dsm_mode,
		dsm_out_sel	=>	dsm_out_sel,
		enable_hclk	=>	enable_hclk,
		enable_idle_atx_pll_support	=>	enable_idle_atx_pll_support,
		enable_lc_calibration	=>	enable_lc_calibration,
		enable_lc_vreg_calibration	=>	enable_lc_vreg_calibration,
		expected_lc_boost_voltage	=>	expected_lc_boost_voltage_int,
		f_max_lcnt_fpll_cascading	=>	f_max_lcnt_fpll_cascading,
		f_max_pfd	=>	f_max_pfd,
		f_max_pfd_fractional	=>	f_max_pfd_fractional,
		f_max_ref	=>	f_max_ref,
		f_max_tank_0	=>	f_max_tank_0,
		f_max_tank_1	=>	f_max_tank_1,
		f_max_tank_2	=>	f_max_tank_2,
		f_max_vco	=>	f_max_vco,
		f_max_vco_fractional	=>	f_max_vco_fractional,
		f_max_x1	=>	f_max_x1,
		f_min_pfd	=>	f_min_pfd,
		f_min_ref	=>	f_min_ref,
		f_min_tank_0	=>	f_min_tank_0,
		f_min_tank_1	=>	f_min_tank_1,
		f_min_tank_2	=>	f_min_tank_2,
		f_min_vco	=>	f_min_vco,
		fb_select	=>	fb_select,
		fpll_refclk_selection	=>	fpll_refclk_selection,
		hclk_divide	=>	hclk_divide,
		initial_settings	=>	initial_settings,
		iqclk_mux_sel	=>	iqclk_mux_sel,
		is_cascaded_pll	=>	is_cascaded_pll,
		is_otn	=>	is_otn,
		is_sdi	=>	is_sdi,
		l_counter	=>	l_counter,
		l_counter_enable	=>	l_counter_enable,
		l_counter_scratch	=>	l_counter_scratch_int,
		lc_atb	=>	lc_atb,
		lc_mode	=>	lc_mode,
		lc_to_fpll_l_counter	=>	lc_to_fpll_l_counter,
		lc_to_fpll_l_counter_scratch	=>	lc_to_fpll_l_counter_scratch_int,
		lf_cbig_size	=>	lf_cbig_size,
		lf_resistance	=>	lf_resistance,
		lf_ripplecap	=>	lf_ripplecap,
		m_counter	=>	m_counter,
		max_fractional_percentage	=>	max_fractional_percentage_int,
		min_fractional_percentage	=>	min_fractional_percentage_int,
		n_counter_scratch	=>	n_counter_scratch_int,
		output_clock_frequency	=>	output_clock_frequency,
		output_regulator_supply	=>	output_regulator_supply,
		overrange_voltage	=>	overrange_voltage,
		pfd_delay_compensation	=>	pfd_delay_compensation,
		pfd_pulse_width	=>	pfd_pulse_width,
		pm_speed_grade	=>	pm_speed_grade,
		pma_width	=>	pma_width,
		power_mode	=>	power_mode,
		power_rail_et	=>	power_rail_et,
		powerdown_mode	=>	powerdown_mode,
		primary_use	=>	primary_use,
		prot_mode	=>	prot_mode,
		ref_clk_div	=>	ref_clk_div,
		reference_clock_frequency	=>	reference_clock_frequency,
		regulator_bypass	=>	regulator_bypass,
		side	=>	side,
		silicon_rev	=>	silicon_rev,
		sup_mode	=>	sup_mode,
		tank_band	=>	tank_band,
		tank_sel	=>	tank_sel,
		tank_voltage_coarse	=>	tank_voltage_coarse,
		tank_voltage_fine	=>	tank_voltage_fine,
		top_or_bottom	=>	top_or_bottom,
		underrange_voltage	=>	underrange_voltage,
		vccdreg_clk	=>	vccdreg_clk,
		vccdreg_fb	=>	vccdreg_fb,
		vccdreg_fw	=>	vccdreg_fw,
		vco_bypass_enable	=>	vco_bypass_enable,
		vco_freq	=>	vco_freq,
		xcpvco_xchgpmplf_cp_current_boost	=>	xcpvco_xchgpmplf_cp_current_boost
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		core_clk	=>	core_clk,
		iqtxrxclk	=>	iqtxrxclk,
		lf_rst_n	=>	lf_rst_n,
		refclk	=>	refclk,
		rst_n	=>	rst_n,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		clk0_16g	=>	clk0_16g,
		clk0_8g	=>	clk0_8g,
		clk180_16g	=>	clk180_16g,
		clk180_8g	=>	clk180_8g,
		clklow_buf	=>	clklow_buf,
		fref_buf	=>	fref_buf,
		hclk_out	=>	hclk_out,
		iqtxrxclk_out	=>	iqtxrxclk_out,
		lc_to_fpll_refclk	=>	lc_to_fpll_refclk,
		lock	=>	lock,
		m_cnt_int	=>	m_cnt_int,
		overrange	=>	overrange,
		underrange	=>	underrange
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_cmu_fpll_refclk_select	is
	generic (
		-- Entity parameters
		mux0_inclk0_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		mux0_inclk1_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		mux0_inclk2_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		mux0_inclk3_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		mux0_inclk4_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		mux1_inclk0_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		mux1_inclk1_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		mux1_inclk2_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		mux1_inclk3_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		mux1_inclk4_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		pll_auto_clk_sw_en	:	string	:=	"false";
		pll_clk_loss_edge	:	string	:=	"pll_clk_loss_both_edges";
		pll_clk_loss_sw_en	:	string	:=	"false";
		pll_clk_sel_override	:	string	:=	"normal";
		pll_clk_sel_override_value	:	string	:=	"select_clk0";
		pll_clk_sw_dly	:	integer	:=	0;
		pll_clkin_0_scratch0_src	:	string	:=	"pll_clkin_0_scratch0_src_vss";
		pll_clkin_0_scratch1_src	:	string	:=	"pll_clkin_0_scratch1_src_vss";
		pll_clkin_0_scratch2_src	:	string	:=	"pll_clkin_0_scratch2_src_vss";
		pll_clkin_0_scratch3_src	:	string	:=	"pll_clkin_0_scratch3_src_vss";
		pll_clkin_0_scratch4_src	:	string	:=	"pll_clkin_0_scratch4_src_vss";
		pll_clkin_0_src	:	string	:=	"pll_clkin_0_src_vss";
		pll_clkin_1_scratch0_src	:	string	:=	"pll_clkin_1_scratch0_src_vss";
		pll_clkin_1_scratch1_src	:	string	:=	"pll_clkin_1_scratch1_src_vss";
		pll_clkin_1_scratch2_src	:	string	:=	"pll_clkin_1_scratch2_src_vss";
		pll_clkin_1_scratch3_src	:	string	:=	"pll_clkin_1_scratch3_src_vss";
		pll_clkin_1_scratch4_src	:	string	:=	"pll_clkin_1_scratch4_src_vss";
		pll_clkin_1_src	:	string	:=	"pll_clkin_1_src_vss";
		pll_manu_clk_sw_en	:	string	:=	"false";
		pll_powerdown_mode	:	string	:=	"false";
		pll_sup_mode	:	string	:=	"user_mode";
		pll_sw_refclk_src	:	string	:=	"pll_sw_refclk_src_clk_0";
		refclk_select0	:	string	:=	"ref_iqclk0";
		refclk_select1	:	string	:=	"ref_iqclk0";
		silicon_rev	:	string	:=	"20nm5es";
		xpm_iqref_mux0_iqclk_sel	:	string	:=	"power_down";
		xpm_iqref_mux0_scratch0_src	:	string	:=	"scratch0_power_down";
		xpm_iqref_mux0_scratch1_src	:	string	:=	"scratch1_power_down";
		xpm_iqref_mux0_scratch2_src	:	string	:=	"scratch2_power_down";
		xpm_iqref_mux0_scratch3_src	:	string	:=	"scratch3_power_down";
		xpm_iqref_mux0_scratch4_src	:	string	:=	"scratch4_power_down";
		xpm_iqref_mux1_iqclk_sel	:	string	:=	"power_down";
		xpm_iqref_mux1_scratch0_src	:	string	:=	"scratch0_power_down";
		xpm_iqref_mux1_scratch1_src	:	string	:=	"scratch1_power_down";
		xpm_iqref_mux1_scratch2_src	:	string	:=	"scratch2_power_down";
		xpm_iqref_mux1_scratch3_src	:	string	:=	"scratch3_power_down";
		xpm_iqref_mux1_scratch4_src	:	string	:=	"scratch4_power_down"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		core_refclk	:	in	std_logic	:=	'0';
		extswitch	:	in	std_logic	:=	'0';
		fpll_cr_pllen	:	in	std_logic	:=	'0';
		iqtxrxclk	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		refclk	:	in	std_logic	:=	'0';
		pll_cascade_in	:	in	std_logic	:=	'0';
		ref_iqclk	:	in	std_logic_vector(11 downto 0)	:=	"000000000000";
		tx_rx_core_refclk	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		clk_src	:	out	std_logic_vector(1 downto 0)	:=	"00";
		clk0bad	:	out	std_logic	:=	'0';
		clk1bad	:	out	std_logic	:=	'0';
		outclk	:	out	std_logic	:=	'0';
		extswitch_buf	:	out	std_logic	:=	'0';
		pllclksel	:	out	std_logic	:=	'0'
	);
end twentynm_cmu_fpll_refclk_select;

architecture behavior of twentynm_cmu_fpll_refclk_select	is




component	twentynm_cmu_fpll_refclk_select_encrypted
	generic (
		-- Architecture parameters
		mux0_inclk0_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		mux0_inclk1_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		mux0_inclk2_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		mux0_inclk3_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		mux0_inclk4_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		mux1_inclk0_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		mux1_inclk1_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		mux1_inclk2_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		mux1_inclk3_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		mux1_inclk4_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		pll_auto_clk_sw_en	:	string	:=	"false";
		pll_clk_loss_edge	:	string	:=	"pll_clk_loss_both_edges";
		pll_clk_loss_sw_en	:	string	:=	"false";
		pll_clk_sel_override	:	string	:=	"normal";
		pll_clk_sel_override_value	:	string	:=	"select_clk0";
		pll_clk_sw_dly	:	integer	:=	0;
		pll_clkin_0_scratch0_src	:	string	:=	"pll_clkin_0_scratch0_src_vss";
		pll_clkin_0_scratch1_src	:	string	:=	"pll_clkin_0_scratch1_src_vss";
		pll_clkin_0_scratch2_src	:	string	:=	"pll_clkin_0_scratch2_src_vss";
		pll_clkin_0_scratch3_src	:	string	:=	"pll_clkin_0_scratch3_src_vss";
		pll_clkin_0_scratch4_src	:	string	:=	"pll_clkin_0_scratch4_src_vss";
		pll_clkin_0_src	:	string	:=	"pll_clkin_0_src_vss";
		pll_clkin_1_scratch0_src	:	string	:=	"pll_clkin_1_scratch0_src_vss";
		pll_clkin_1_scratch1_src	:	string	:=	"pll_clkin_1_scratch1_src_vss";
		pll_clkin_1_scratch2_src	:	string	:=	"pll_clkin_1_scratch2_src_vss";
		pll_clkin_1_scratch3_src	:	string	:=	"pll_clkin_1_scratch3_src_vss";
		pll_clkin_1_scratch4_src	:	string	:=	"pll_clkin_1_scratch4_src_vss";
		pll_clkin_1_src	:	string	:=	"pll_clkin_1_src_vss";
		pll_manu_clk_sw_en	:	string	:=	"false";
		pll_powerdown_mode	:	string	:=	"false";
		pll_sup_mode	:	string	:=	"user_mode";
		pll_sw_refclk_src	:	string	:=	"pll_sw_refclk_src_clk_0";
		refclk_select0	:	string	:=	"ref_iqclk0";
		refclk_select1	:	string	:=	"ref_iqclk0";
		silicon_rev	:	string	:=	"20nm5es";
		xpm_iqref_mux0_iqclk_sel	:	string	:=	"power_down";
		xpm_iqref_mux0_scratch0_src	:	string	:=	"scratch0_power_down";
		xpm_iqref_mux0_scratch1_src	:	string	:=	"scratch1_power_down";
		xpm_iqref_mux0_scratch2_src	:	string	:=	"scratch2_power_down";
		xpm_iqref_mux0_scratch3_src	:	string	:=	"scratch3_power_down";
		xpm_iqref_mux0_scratch4_src	:	string	:=	"scratch4_power_down";
		xpm_iqref_mux1_iqclk_sel	:	string	:=	"power_down";
		xpm_iqref_mux1_scratch0_src	:	string	:=	"scratch0_power_down";
		xpm_iqref_mux1_scratch1_src	:	string	:=	"scratch1_power_down";
		xpm_iqref_mux1_scratch2_src	:	string	:=	"scratch2_power_down";
		xpm_iqref_mux1_scratch3_src	:	string	:=	"scratch3_power_down";
		xpm_iqref_mux1_scratch4_src	:	string	:=	"scratch4_power_down"
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		core_refclk	:	in	std_logic	:=	'0';
		extswitch	:	in	std_logic	:=	'0';
		fpll_cr_pllen	:	in	std_logic	:=	'0';
		iqtxrxclk	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		refclk	:	in	std_logic	:=	'0';
		pll_cascade_in	:	in	std_logic	:=	'0';
		ref_iqclk	:	in	std_logic_vector(11 downto 0)	:=	"000000000000";
		tx_rx_core_refclk	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		clk_src	:	out	std_logic_vector(1 downto 0)	:=	"00";
		clk0bad	:	out	std_logic	:=	'0';
		clk1bad	:	out	std_logic	:=	'0';
		outclk	:	out	std_logic	:=	'0';
		extswitch_buf	:	out	std_logic	:=	'0';
		pllclksel	:	out	std_logic	:=	'0'
	);
end component;

begin



inst : twentynm_cmu_fpll_refclk_select_encrypted
	generic map (
		-- Instance parameters
		mux0_inclk0_logical_to_physical_mapping	=>	mux0_inclk0_logical_to_physical_mapping,
		mux0_inclk1_logical_to_physical_mapping	=>	mux0_inclk1_logical_to_physical_mapping,
		mux0_inclk2_logical_to_physical_mapping	=>	mux0_inclk2_logical_to_physical_mapping,
		mux0_inclk3_logical_to_physical_mapping	=>	mux0_inclk3_logical_to_physical_mapping,
		mux0_inclk4_logical_to_physical_mapping	=>	mux0_inclk4_logical_to_physical_mapping,
		mux1_inclk0_logical_to_physical_mapping	=>	mux1_inclk0_logical_to_physical_mapping,
		mux1_inclk1_logical_to_physical_mapping	=>	mux1_inclk1_logical_to_physical_mapping,
		mux1_inclk2_logical_to_physical_mapping	=>	mux1_inclk2_logical_to_physical_mapping,
		mux1_inclk3_logical_to_physical_mapping	=>	mux1_inclk3_logical_to_physical_mapping,
		mux1_inclk4_logical_to_physical_mapping	=>	mux1_inclk4_logical_to_physical_mapping,
		pll_auto_clk_sw_en	=>	pll_auto_clk_sw_en,
		pll_clk_loss_edge	=>	pll_clk_loss_edge,
		pll_clk_loss_sw_en	=>	pll_clk_loss_sw_en,
		pll_clk_sel_override	=>	pll_clk_sel_override,
		pll_clk_sel_override_value	=>	pll_clk_sel_override_value,
		pll_clk_sw_dly	=>	pll_clk_sw_dly,
		pll_clkin_0_scratch0_src	=>	pll_clkin_0_scratch0_src,
		pll_clkin_0_scratch1_src	=>	pll_clkin_0_scratch1_src,
		pll_clkin_0_scratch2_src	=>	pll_clkin_0_scratch2_src,
		pll_clkin_0_scratch3_src	=>	pll_clkin_0_scratch3_src,
		pll_clkin_0_scratch4_src	=>	pll_clkin_0_scratch4_src,
		pll_clkin_0_src	=>	pll_clkin_0_src,
		pll_clkin_1_scratch0_src	=>	pll_clkin_1_scratch0_src,
		pll_clkin_1_scratch1_src	=>	pll_clkin_1_scratch1_src,
		pll_clkin_1_scratch2_src	=>	pll_clkin_1_scratch2_src,
		pll_clkin_1_scratch3_src	=>	pll_clkin_1_scratch3_src,
		pll_clkin_1_scratch4_src	=>	pll_clkin_1_scratch4_src,
		pll_clkin_1_src	=>	pll_clkin_1_src,
		pll_manu_clk_sw_en	=>	pll_manu_clk_sw_en,
		pll_powerdown_mode	=>	pll_powerdown_mode,
		pll_sup_mode	=>	pll_sup_mode,
		pll_sw_refclk_src	=>	pll_sw_refclk_src,
		refclk_select0	=>	refclk_select0,
		refclk_select1	=>	refclk_select1,
		silicon_rev	=>	silicon_rev,
		xpm_iqref_mux0_iqclk_sel	=>	xpm_iqref_mux0_iqclk_sel,
		xpm_iqref_mux0_scratch0_src	=>	xpm_iqref_mux0_scratch0_src,
		xpm_iqref_mux0_scratch1_src	=>	xpm_iqref_mux0_scratch1_src,
		xpm_iqref_mux0_scratch2_src	=>	xpm_iqref_mux0_scratch2_src,
		xpm_iqref_mux0_scratch3_src	=>	xpm_iqref_mux0_scratch3_src,
		xpm_iqref_mux0_scratch4_src	=>	xpm_iqref_mux0_scratch4_src,
		xpm_iqref_mux1_iqclk_sel	=>	xpm_iqref_mux1_iqclk_sel,
		xpm_iqref_mux1_scratch0_src	=>	xpm_iqref_mux1_scratch0_src,
		xpm_iqref_mux1_scratch1_src	=>	xpm_iqref_mux1_scratch1_src,
		xpm_iqref_mux1_scratch2_src	=>	xpm_iqref_mux1_scratch2_src,
		xpm_iqref_mux1_scratch3_src	=>	xpm_iqref_mux1_scratch3_src,
		xpm_iqref_mux1_scratch4_src	=>	xpm_iqref_mux1_scratch4_src
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		core_refclk	=>	core_refclk,
		extswitch	=>	extswitch,
		fpll_cr_pllen	=>	fpll_cr_pllen,
		iqtxrxclk	=>	iqtxrxclk,
		refclk	=>	refclk,
		pll_cascade_in	=>	pll_cascade_in,
		ref_iqclk	=>	ref_iqclk,
		tx_rx_core_refclk	=>	tx_rx_core_refclk,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		clk_src	=>	clk_src,
		clk0bad	=>	clk0bad,
		clk1bad	=>	clk1bad,
		outclk	=>	outclk,
		extswitch_buf	=>	extswitch_buf,
		pllclksel	=>	pllclksel
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_cmu_fpll	is
	generic (
		-- Entity parameters
		analog_mode	:	string	:=	"user_custom";
		bandwidth_range_high	:	string	:=	"000000000000000000000000000000000001";
		bandwidth_range_low	:	string	:=	"000000000000000000000000000000000001";
		bonding	:	string	:=	"pll_bonding";
		bw_sel	:	string	:=	"auto";
		cgb_div	:	integer	:=	1;
		compensation_mode	:	string	:=	"direct";
		datarate	:	string	:=	"0 bps";
		duty_cycle_0	:	integer	:=	50;
		duty_cycle_1	:	integer	:=	50;
		duty_cycle_2	:	integer	:=	50;
		duty_cycle_3	:	integer	:=	50;
		enable_idle_fpll_support	:	string	:=	"idle_none";
		f_max_band_0	:	string	:=	"000000000000000000000000000000000001";
		f_max_band_1	:	string	:=	"000000000000000000000000000000000001";
		f_max_band_2	:	string	:=	"000000000000000000000000000000000001";
		f_max_band_3	:	string	:=	"000000000000000000000000000000000001";
		f_max_band_4	:	string	:=	"000000000000000000000000000000000001";
		f_max_band_5	:	string	:=	"000000000000000000000000000000000001";
		f_max_band_6	:	string	:=	"000000000000000000000000000000000001";
		f_max_band_7	:	string	:=	"000000000000000000000000000000000001";
		f_max_band_8	:	string	:=	"000000000000000000000000000000000001";
		f_max_band_9	:	string	:=	"000000000000000000000000000000000001";
		f_max_div_two_bypass	:	string	:=	"000000000000000000000000000000000001";
		f_max_pfd	:	string	:=	"000000000000000000000000000000000001";
		f_max_pfd_bonded	:	string	:=	"000000000000000000000000000000000001";
		f_max_pfd_fractional	:	string	:=	"000000000000000000000000000001011111";
		f_max_pfd_integer	:	string	:=	"000000000000000000000000000000000001";
		f_max_vco	:	string	:=	"000000000000000000000000000000000001";
		f_max_vco_fractional	:	string	:=	"000000000000000000000000000000000101";
		f_min_band_0	:	string	:=	"000000000000000000000000000000000001";
		f_min_band_1	:	string	:=	"000000000000000000000000000000000001";
		f_min_band_2	:	string	:=	"000000000000000000000000000000000001";
		f_min_band_3	:	string	:=	"000000000000000000000000000000000001";
		f_min_band_4	:	string	:=	"000000000000000000000000000000000001";
		f_min_band_5	:	string	:=	"000000000000000000000000000000000001";
		f_min_band_6	:	string	:=	"000000000000000000000000000000000001";
		f_min_band_7	:	string	:=	"000000000000000000000000000000000001";
		f_min_band_8	:	string	:=	"000000000000000000000000000000000001";
		f_min_band_9	:	string	:=	"000000000000000000000000000000000001";
		f_min_pfd	:	string	:=	"000000000000000000000000000000000001";
		f_min_vco	:	string	:=	"000000000000000000000000000000000001";
		f_out_c0	:	string	:=	"000000000000000000000000000000000001";
		f_out_c0_hz	:	string	:=	"0 hz";
		f_out_c1	:	string	:=	"000000000000000000000000000000000001";
		f_out_c1_hz	:	string	:=	"0 hz";
		f_out_c2	:	string	:=	"000000000000000000000000000000000001";
		f_out_c2_hz	:	string	:=	"0 hz";
		f_out_c3	:	string	:=	"000000000000000000000000000000000001";
		f_out_c3_hz	:	string	:=	"0 hz";
		feedback	:	string	:=	"normal";
		fpll_cal_test_sel	:	string	:=	"sel_cal_out_7_to_0";
		fpll_cas_out_enable	:	string	:=	"fpll_cas_out_disable";
		fpll_hclk_out_enable	:	string	:=	"fpll_hclk_out_disable";
		fpll_iqtxrxclk_out_enable	:	string	:=	"fpll_iqtxrxclk_out_disable";
		hssi_output_clock_frequency	:	string	:=	"0 ps";
		initial_settings	:	string	:=	"true";
		input_tolerance	:	bit_vector	:=	B"00000000";
		is_cascaded_pll	:	string	:=	"false";
		is_otn	:	string	:=	"false";
		is_pa_core	:	string	:=	"false";
		is_sdi	:	string	:=	"false";
		l_counter	:	bit_vector	:=	B"000001";
		m_counter	:	bit_vector	:=	B"00000001";
		m_counter_c0	:	bit_vector	:=	B"000000000";
		m_counter_c1	:	bit_vector	:=	B"000000000";
		m_counter_c2	:	bit_vector	:=	B"000000000";
		m_counter_c3	:	bit_vector	:=	B"000000000";
		max_fractional_percentage	:	bit_vector	:=	B"0000000";
		min_fractional_percentage	:	bit_vector	:=	B"0000000";
		n_counter	:	bit_vector	:=	B"000001";
		out_freq	:	string	:=	"000000000000000000000000000000000001";
		out_freq_hz	:	string	:=	"0 hz";
		output_clock_frequency_0	:	string	:=	"0 ps";
		output_clock_frequency_1	:	string	:=	"0 ps";
		output_clock_frequency_2	:	string	:=	"0 ps";
		output_clock_frequency_3	:	string	:=	"0 ps";
		output_tolerance	:	bit_vector	:=	B"00000000";
		pfd_freq	:	string	:=	"000000000000000000000000000000000001";
		phase_shift_0	:	string	:=	"0 ps";
		phase_shift_1	:	string	:=	"0 ps";
		phase_shift_2	:	string	:=	"0 ps";
		phase_shift_3	:	string	:=	"0 ps";
		pll_atb	:	string	:=	"atb_selectdisable";
		pll_bw_mode	:	string	:=	"low_bw";
		pll_c0_pllcout_enable	:	string	:=	"false";
		pll_c1_pllcout_enable	:	string	:=	"false";
		pll_c2_pllcout_enable	:	string	:=	"false";
		pll_c3_pllcout_enable	:	string	:=	"false";
		pll_c_counter_0	:	integer	:=	1;
		pll_c_counter_0_coarse_dly	:	string	:=	"0 ps";
		pll_c_counter_0_fine_dly	:	string	:=	"0 ps";
		pll_c_counter_0_in_src	:	string	:=	"m_cnt_in_src_test_clk";
		pll_c_counter_0_min_tco_enable	:	string	:=	"true";
		pll_c_counter_0_ph_mux_prst	:	integer	:=	0;
		pll_c_counter_0_prst	:	integer	:=	1;
		pll_c_counter_1	:	integer	:=	1;
		pll_c_counter_1_coarse_dly	:	string	:=	"0 ps";
		pll_c_counter_1_fine_dly	:	string	:=	"0 ps";
		pll_c_counter_1_in_src	:	string	:=	"m_cnt_in_src_test_clk";
		pll_c_counter_1_min_tco_enable	:	string	:=	"true";
		pll_c_counter_1_ph_mux_prst	:	integer	:=	0;
		pll_c_counter_1_prst	:	integer	:=	1;
		pll_c_counter_2	:	integer	:=	1;
		pll_c_counter_2_coarse_dly	:	string	:=	"0 ps";
		pll_c_counter_2_fine_dly	:	string	:=	"0 ps";
		pll_c_counter_2_in_src	:	string	:=	"m_cnt_in_src_test_clk";
		pll_c_counter_2_min_tco_enable	:	string	:=	"true";
		pll_c_counter_2_ph_mux_prst	:	integer	:=	0;
		pll_c_counter_2_prst	:	integer	:=	1;
		pll_c_counter_3	:	integer	:=	1;
		pll_c_counter_3_coarse_dly	:	string	:=	"0 ps";
		pll_c_counter_3_fine_dly	:	string	:=	"0 ps";
		pll_c_counter_3_in_src	:	string	:=	"m_cnt_in_src_test_clk";
		pll_c_counter_3_min_tco_enable	:	string	:=	"true";
		pll_c_counter_3_ph_mux_prst	:	integer	:=	0;
		pll_c_counter_3_prst	:	integer	:=	1;
		pll_cal_status	:	string	:=	"true";
		pll_calibration	:	string	:=	"false";
		pll_cmp_buf_dly	:	string	:=	"0 ps";
		pll_cmu_rstn_value	:	string	:=	"true";
		pll_core_cali_ref_off	:	string	:=	"true";
		pll_core_cali_vco_off	:	string	:=	"true";
		pll_core_vccdreg_fb	:	string	:=	"vreg_fb0";
		pll_core_vccdreg_fw	:	string	:=	"vreg_fw0";
		pll_core_vreg0_atbsel	:	string	:=	"atb_disabled";
		pll_core_vreg1_atbsel	:	string	:=	"atb_disabled1";
		pll_cp_compensation	:	string	:=	"true";
		pll_cp_current_setting	:	string	:=	"cp_current_setting0";
		pll_cp_lf_3rd_pole_freq	:	string	:=	"lf_3rd_pole_setting0";
		pll_cp_lf_order	:	string	:=	"lf_2nd_order";
		pll_cp_testmode	:	string	:=	"cp_normal";
		pll_ctrl_override_setting	:	string	:=	"true";
		pll_ctrl_plniotri_override	:	string	:=	"false";
		pll_device_variant	:	string	:=	"device1";
		pll_dprio_base_addr	:	integer	:=	256;
		pll_dprio_broadcast_en	:	string	:=	"false";
		pll_dprio_clk_vreg_boost	:	string	:=	"clk_fpll_vreg_no_voltage_boost";
		pll_dprio_cvp_inter_sel	:	string	:=	"true";
		pll_dprio_force_inter_sel	:	string	:=	"false";
		pll_dprio_fpll_vreg1_boost	:	string	:=	"fpll_vreg1_no_voltage_boost";
		pll_dprio_fpll_vreg_boost	:	string	:=	"fpll_vreg_no_voltage_boost";
		pll_dprio_power_iso_en	:	string	:=	"true";
		pll_dprio_status_select	:	string	:=	"dprio_normal_status";
		pll_dsm_ecn_bypass	:	string	:=	"false";
		pll_dsm_ecn_test_en	:	string	:=	"false";
		pll_dsm_fractional_division	:	string	:=	"00000000000000000000000000000000";
		pll_dsm_fractional_value_ready	:	string	:=	"pll_k_ready";
		pll_dsm_mode	:	string	:=	"dsm_mode_integer";
		pll_dsm_out_sel	:	string	:=	"pll_dsm_disable";
		pll_enable	:	string	:=	"false";
		pll_extra_csr	:	integer	:=	0;
		pll_fbclk_mux_1	:	string	:=	"pll_fbclk_mux_1_glb";
		pll_fbclk_mux_2	:	string	:=	"pll_fbclk_mux_2_fb_1";
		pll_iqclk_mux_sel	:	string	:=	"power_down";
		pll_l_counter	:	integer	:=	1;
		pll_l_counter_bypass	:	string	:=	"false";
		pll_l_counter_enable	:	string	:=	"true";
		pll_lf_cbig	:	string	:=	"lf_cbig_setting0";
		pll_lf_resistance	:	string	:=	"lf_res_setting0";
		pll_lf_ripplecap	:	string	:=	"lf_ripple_enabled_0";
		pll_lock_fltr_cfg	:	integer	:=	1;
		pll_lock_fltr_test	:	string	:=	"pll_lock_fltr_nrm";
		pll_lpf_rstn_value	:	string	:=	"lpf_normal";
		pll_m_counter	:	integer	:=	1;
		pll_m_counter_coarse_dly	:	string	:=	"0 ps";
		pll_m_counter_fine_dly	:	string	:=	"0 ps";
		pll_m_counter_in_src	:	string	:=	"m_cnt_in_src_test_clk";
		pll_m_counter_min_tco_enable	:	string	:=	"true";
		pll_m_counter_ph_mux_prst	:	integer	:=	0;
		pll_m_counter_prst	:	integer	:=	1;
		pll_n_counter	:	integer	:=	1;
		pll_n_counter_coarse_dly	:	string	:=	"0 ps";
		pll_n_counter_fine_dly	:	string	:=	"0 ps";
		pll_nreset_invert	:	string	:=	"false";
		pll_op_mode	:	string	:=	"false";
		pll_optimal	:	string	:=	"true";
		pll_powerdown_mode	:	string	:=	"false";
		pll_ppm_clk0_src	:	string	:=	"ppm_clk0_vss";
		pll_ppm_clk1_src	:	string	:=	"ppm_clk1_vss";
		pll_ref_buf_dly	:	string	:=	"0 ps";
		pll_rstn_override	:	string	:=	"false";
		pll_self_reset	:	string	:=	"false";
		pll_sup_mode	:	string	:=	"user_mode";
		pll_tclk_mux_en	:	string	:=	"false";
		pll_tclk_sel	:	string	:=	"pll_tclk_m_src";
		pll_test_enable	:	string	:=	"false";
		pll_unlock_fltr_cfg	:	integer	:=	0;
		pll_vccr_pd_en	:	string	:=	"false";
		pll_vco_freq_band_0	:	string	:=	"pll_freq_band0";
		pll_vco_freq_band_0_dyn_high_bits	:	bit_vector	:=	B"00";
		pll_vco_freq_band_0_dyn_low_bits	:	bit_vector	:=	B"000";
		pll_vco_freq_band_0_fix	:	bit_vector	:=	B"00001";
		pll_vco_freq_band_0_fix_high	:	string	:=	"pll_vco_freq_band_0_fix_high_0";
		pll_vco_freq_band_1	:	string	:=	"pll_freq_band0_1";
		pll_vco_freq_band_1_dyn_high_bits	:	bit_vector	:=	B"00";
		pll_vco_freq_band_1_dyn_low_bits	:	bit_vector	:=	B"000";
		pll_vco_freq_band_1_fix	:	bit_vector	:=	B"00001";
		pll_vco_freq_band_1_fix_high	:	string	:=	"pll_vco_freq_band_1_fix_high_0";
		pll_vco_ph0_en	:	string	:=	"false";
		pll_vco_ph0_value	:	string	:=	"pll_vco_ph0_vss";
		pll_vco_ph1_en	:	string	:=	"false";
		pll_vco_ph1_value	:	string	:=	"pll_vco_ph1_vss";
		pll_vco_ph2_en	:	string	:=	"false";
		pll_vco_ph2_value	:	string	:=	"pll_vco_ph2_vss";
		pll_vco_ph3_en	:	string	:=	"false";
		pll_vco_ph3_value	:	string	:=	"pll_vco_ph3_vss";
		pm_speed_grade	:	string	:=	"e2";
		pma_width	:	integer	:=	8;
		power_mode	:	string	:=	"low_power";
		power_rail_et	:	integer	:=	0;
		primary_use	:	string	:=	"tx";
		prot_mode	:	string	:=	"basic_tx";
		reference_clock_frequency	:	string	:=	"0 ps";
		reference_clock_frequency_scratch	:	string	:=	"0 hz";
		set_fpll_input_freq_range	:	bit_vector	:=	B"00000000";
		side	:	string	:=	"side_unknown";
		silicon_rev	:	string	:=	"20nm5es";
		top_or_bottom	:	string	:=	"tb_unknown";
		vco_freq	:	string	:=	"000000000000000000000000000000000001";
		vco_freq_hz	:	string	:=	"0 hz";
		vco_frequency	:	string	:=	"0 ps";
		xpm_cmu_fpll_core_cal_vco_count_length	:	string	:=	"sel_8b_count";
		xpm_cmu_fpll_core_fpll_refclk_source	:	string	:=	"normal_refclk";
		xpm_cmu_fpll_core_fpll_vco_div_by_2_sel	:	string	:=	"bypass_divide_by_2";
		xpm_cmu_fpll_core_pfd_delay_compensation	:	string	:=	"normal_delay";
		xpm_cmu_fpll_core_pfd_pulse_width	:	string	:=	"pulse_width_setting0";
		xpm_cmu_fpll_core_xpm_cpvco_fpll_xpm_chgpmplf_fpll_cp_current_boost	:	string	:=	"normal_setting"
	);
	port (
		-- Entity ports
		clk0bad_in	:	in	std_logic	:=	'0';
		clk1bad_in	:	in	std_logic	:=	'0';
		cnt_sel	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		core_refclk	:	in	std_logic	:=	'0';
		csr_bufin	:	in	std_logic	:=	'0';
		csr_clk	:	in	std_logic	:=	'0';
		csr_en	:	in	std_logic	:=	'0';
		csr_en_dly	:	in	std_logic	:=	'0';
		csr_in	:	in	std_logic	:=	'0';
		avmmclk	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		dps_rst_n	:	in	std_logic	:=	'0';
		extswitch_buf	:	in	std_logic	:=	'0';
		fbclk_in	:	in	std_logic	:=	'0';
		fpll_ppm_clk	:	in	std_logic_vector(1 downto 0)	:=	"00";
		iqtxrxclk	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		lc_to_fpll_refclk	:	in	std_logic	:=	'0';
		mdio_dis	:	in	std_logic	:=	'0';
		nfrzdrv	:	in	std_logic	:=	'0';
		nrpi_freeze	:	in	std_logic	:=	'0';
		num_phase_shifts	:	in	std_logic_vector(2 downto 0)	:=	"000";
		pfden	:	in	std_logic	:=	'0';
		phase_en	:	in	std_logic	:=	'0';
		pllclksel	:	in	std_logic	:=	'0';
		pma_atpg_los_en_n	:	in	std_logic	:=	'0';
		pma_csr_test_dis	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		refclk	:	in	std_logic	:=	'0';
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		rst_n	:	in	std_logic	:=	'0';
		scan_mode_n	:	in	std_logic	:=	'0';
		scan_shift_n	:	in	std_logic	:=	'0';
		up_dn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		block_select	:	out	std_logic	:=	'0';
		clk0	:	out	std_logic	:=	'0';
		clk0bad	:	out	std_logic	:=	'0';
		clk180	:	out	std_logic	:=	'0';
		clk1bad	:	out	std_logic	:=	'0';
		clklow	:	out	std_logic	:=	'0';
		csr_bufout	:	out	std_logic	:=	'0';
		csr_out	:	out	std_logic	:=	'0';
		fbclk_out	:	out	std_logic	:=	'0';
		clk_sel_override	:	out	std_logic	:=	'0';
		clk_sel_override_value	:	out	std_logic	:=	'0';
		fref	:	out	std_logic	:=	'0';
		hclk_out	:	out	std_logic	:=	'0';
		iqtxrxclk_out	:	out	std_logic	:=	'0';
		lock	:	out	std_logic	:=	'0';
		phase_done	:	out	std_logic	:=	'0';
		pll_cascade_out	:	out	std_logic	:=	'0';
		outclk	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		ppm_clk	:	out	std_logic_vector(1 downto 0)	:=	"00";
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000"
	);
end twentynm_cmu_fpll;

architecture behavior of twentynm_cmu_fpll	is

constant input_tolerance_int	:	integer	:=	bin2int(input_tolerance);
constant l_counter_int	:	integer	:=	bin2int(l_counter);
constant m_counter_int	:	integer	:=	bin2int(m_counter);
constant m_counter_c0_int	:	integer	:=	bin2int(m_counter_c0);
constant m_counter_c1_int	:	integer	:=	bin2int(m_counter_c1);
constant m_counter_c2_int	:	integer	:=	bin2int(m_counter_c2);
constant m_counter_c3_int	:	integer	:=	bin2int(m_counter_c3);
constant max_fractional_percentage_int	:	integer	:=	bin2int(max_fractional_percentage);
constant min_fractional_percentage_int	:	integer	:=	bin2int(min_fractional_percentage);
constant n_counter_int	:	integer	:=	bin2int(n_counter);
constant output_tolerance_int	:	integer	:=	bin2int(output_tolerance);
constant pll_vco_freq_band_0_dyn_high_bits_int	:	integer	:=	bin2int(pll_vco_freq_band_0_dyn_high_bits);
constant pll_vco_freq_band_0_dyn_low_bits_int	:	integer	:=	bin2int(pll_vco_freq_band_0_dyn_low_bits);
constant pll_vco_freq_band_0_fix_int	:	integer	:=	bin2int(pll_vco_freq_band_0_fix);
constant pll_vco_freq_band_1_dyn_high_bits_int	:	integer	:=	bin2int(pll_vco_freq_band_1_dyn_high_bits);
constant pll_vco_freq_band_1_dyn_low_bits_int	:	integer	:=	bin2int(pll_vco_freq_band_1_dyn_low_bits);
constant pll_vco_freq_band_1_fix_int	:	integer	:=	bin2int(pll_vco_freq_band_1_fix);
constant set_fpll_input_freq_range_int	:	integer	:=	bin2int(set_fpll_input_freq_range);



component	twentynm_cmu_fpll_encrypted
	generic (
		-- Architecture parameters
		analog_mode	:	string	:=	"user_custom";
		bandwidth_range_high	:	string	:=	"000000000000000000000000000000000001";
		bandwidth_range_low	:	string	:=	"000000000000000000000000000000000001";
		bonding	:	string	:=	"pll_bonding";
		bw_sel	:	string	:=	"auto";
		cgb_div	:	integer	:=	1;
		compensation_mode	:	string	:=	"direct";
		datarate	:	string	:=	"0 bps";
		duty_cycle_0	:	integer	:=	50;
		duty_cycle_1	:	integer	:=	50;
		duty_cycle_2	:	integer	:=	50;
		duty_cycle_3	:	integer	:=	50;
		enable_idle_fpll_support	:	string	:=	"idle_none";
		f_max_band_0	:	string	:=	"000000000000000000000000000000000001";
		f_max_band_1	:	string	:=	"000000000000000000000000000000000001";
		f_max_band_2	:	string	:=	"000000000000000000000000000000000001";
		f_max_band_3	:	string	:=	"000000000000000000000000000000000001";
		f_max_band_4	:	string	:=	"000000000000000000000000000000000001";
		f_max_band_5	:	string	:=	"000000000000000000000000000000000001";
		f_max_band_6	:	string	:=	"000000000000000000000000000000000001";
		f_max_band_7	:	string	:=	"000000000000000000000000000000000001";
		f_max_band_8	:	string	:=	"000000000000000000000000000000000001";
		f_max_band_9	:	string	:=	"000000000000000000000000000000000001";
		f_max_div_two_bypass	:	string	:=	"000000000000000000000000000000000001";
		f_max_pfd	:	string	:=	"000000000000000000000000000000000001";
		f_max_pfd_bonded	:	string	:=	"000000000000000000000000000000000001";
		f_max_pfd_fractional	:	string	:=	"000000000000000000000000000001011111";
		f_max_pfd_integer	:	string	:=	"000000000000000000000000000000000001";
		f_max_vco	:	string	:=	"000000000000000000000000000000000001";
		f_max_vco_fractional	:	string	:=	"000000000000000000000000000000000101";
		f_min_band_0	:	string	:=	"000000000000000000000000000000000001";
		f_min_band_1	:	string	:=	"000000000000000000000000000000000001";
		f_min_band_2	:	string	:=	"000000000000000000000000000000000001";
		f_min_band_3	:	string	:=	"000000000000000000000000000000000001";
		f_min_band_4	:	string	:=	"000000000000000000000000000000000001";
		f_min_band_5	:	string	:=	"000000000000000000000000000000000001";
		f_min_band_6	:	string	:=	"000000000000000000000000000000000001";
		f_min_band_7	:	string	:=	"000000000000000000000000000000000001";
		f_min_band_8	:	string	:=	"000000000000000000000000000000000001";
		f_min_band_9	:	string	:=	"000000000000000000000000000000000001";
		f_min_pfd	:	string	:=	"000000000000000000000000000000000001";
		f_min_vco	:	string	:=	"000000000000000000000000000000000001";
		f_out_c0	:	string	:=	"000000000000000000000000000000000001";
		f_out_c0_hz	:	string	:=	"0 hz";
		f_out_c1	:	string	:=	"000000000000000000000000000000000001";
		f_out_c1_hz	:	string	:=	"0 hz";
		f_out_c2	:	string	:=	"000000000000000000000000000000000001";
		f_out_c2_hz	:	string	:=	"0 hz";
		f_out_c3	:	string	:=	"000000000000000000000000000000000001";
		f_out_c3_hz	:	string	:=	"0 hz";
		feedback	:	string	:=	"normal";
		fpll_cal_test_sel	:	string	:=	"sel_cal_out_7_to_0";
		fpll_cas_out_enable	:	string	:=	"fpll_cas_out_disable";
		fpll_hclk_out_enable	:	string	:=	"fpll_hclk_out_disable";
		fpll_iqtxrxclk_out_enable	:	string	:=	"fpll_iqtxrxclk_out_disable";
		hssi_output_clock_frequency	:	string	:=	"0 ps";
		initial_settings	:	string	:=	"true";
		input_tolerance	:	integer	:=	0;
		is_cascaded_pll	:	string	:=	"false";
		is_otn	:	string	:=	"false";
		is_pa_core	:	string	:=	"false";
		is_sdi	:	string	:=	"false";
		l_counter	:	integer	:=	1;
		m_counter	:	integer	:=	1;
		m_counter_c0	:	integer	:=	0;
		m_counter_c1	:	integer	:=	0;
		m_counter_c2	:	integer	:=	0;
		m_counter_c3	:	integer	:=	0;
		max_fractional_percentage	:	integer	:=	0;
		min_fractional_percentage	:	integer	:=	0;
		n_counter	:	integer	:=	1;
		out_freq	:	string	:=	"000000000000000000000000000000000001";
		out_freq_hz	:	string	:=	"0 hz";
		output_clock_frequency_0	:	string	:=	"0 ps";
		output_clock_frequency_1	:	string	:=	"0 ps";
		output_clock_frequency_2	:	string	:=	"0 ps";
		output_clock_frequency_3	:	string	:=	"0 ps";
		output_tolerance	:	integer	:=	0;
		pfd_freq	:	string	:=	"000000000000000000000000000000000001";
		phase_shift_0	:	string	:=	"0 ps";
		phase_shift_1	:	string	:=	"0 ps";
		phase_shift_2	:	string	:=	"0 ps";
		phase_shift_3	:	string	:=	"0 ps";
		pll_atb	:	string	:=	"atb_selectdisable";
		pll_bw_mode	:	string	:=	"low_bw";
		pll_c0_pllcout_enable	:	string	:=	"false";
		pll_c1_pllcout_enable	:	string	:=	"false";
		pll_c2_pllcout_enable	:	string	:=	"false";
		pll_c3_pllcout_enable	:	string	:=	"false";
		pll_c_counter_0	:	integer	:=	1;
		pll_c_counter_0_coarse_dly	:	string	:=	"0 ps";
		pll_c_counter_0_fine_dly	:	string	:=	"0 ps";
		pll_c_counter_0_in_src	:	string	:=	"m_cnt_in_src_test_clk";
		pll_c_counter_0_min_tco_enable	:	string	:=	"true";
		pll_c_counter_0_ph_mux_prst	:	integer	:=	0;
		pll_c_counter_0_prst	:	integer	:=	1;
		pll_c_counter_1	:	integer	:=	1;
		pll_c_counter_1_coarse_dly	:	string	:=	"0 ps";
		pll_c_counter_1_fine_dly	:	string	:=	"0 ps";
		pll_c_counter_1_in_src	:	string	:=	"m_cnt_in_src_test_clk";
		pll_c_counter_1_min_tco_enable	:	string	:=	"true";
		pll_c_counter_1_ph_mux_prst	:	integer	:=	0;
		pll_c_counter_1_prst	:	integer	:=	1;
		pll_c_counter_2	:	integer	:=	1;
		pll_c_counter_2_coarse_dly	:	string	:=	"0 ps";
		pll_c_counter_2_fine_dly	:	string	:=	"0 ps";
		pll_c_counter_2_in_src	:	string	:=	"m_cnt_in_src_test_clk";
		pll_c_counter_2_min_tco_enable	:	string	:=	"true";
		pll_c_counter_2_ph_mux_prst	:	integer	:=	0;
		pll_c_counter_2_prst	:	integer	:=	1;
		pll_c_counter_3	:	integer	:=	1;
		pll_c_counter_3_coarse_dly	:	string	:=	"0 ps";
		pll_c_counter_3_fine_dly	:	string	:=	"0 ps";
		pll_c_counter_3_in_src	:	string	:=	"m_cnt_in_src_test_clk";
		pll_c_counter_3_min_tco_enable	:	string	:=	"true";
		pll_c_counter_3_ph_mux_prst	:	integer	:=	0;
		pll_c_counter_3_prst	:	integer	:=	1;
		pll_cal_status	:	string	:=	"true";
		pll_calibration	:	string	:=	"false";
		pll_cmp_buf_dly	:	string	:=	"0 ps";
		pll_cmu_rstn_value	:	string	:=	"true";
		pll_core_cali_ref_off	:	string	:=	"true";
		pll_core_cali_vco_off	:	string	:=	"true";
		pll_core_vccdreg_fb	:	string	:=	"vreg_fb0";
		pll_core_vccdreg_fw	:	string	:=	"vreg_fw0";
		pll_core_vreg0_atbsel	:	string	:=	"atb_disabled";
		pll_core_vreg1_atbsel	:	string	:=	"atb_disabled1";
		pll_cp_compensation	:	string	:=	"true";
		pll_cp_current_setting	:	string	:=	"cp_current_setting0";
		pll_cp_lf_3rd_pole_freq	:	string	:=	"lf_3rd_pole_setting0";
		pll_cp_lf_order	:	string	:=	"lf_2nd_order";
		pll_cp_testmode	:	string	:=	"cp_normal";
		pll_ctrl_override_setting	:	string	:=	"true";
		pll_ctrl_plniotri_override	:	string	:=	"false";
		pll_device_variant	:	string	:=	"device1";
		pll_dprio_base_addr	:	integer	:=	256;
		pll_dprio_broadcast_en	:	string	:=	"false";
		pll_dprio_clk_vreg_boost	:	string	:=	"clk_fpll_vreg_no_voltage_boost";
		pll_dprio_cvp_inter_sel	:	string	:=	"true";
		pll_dprio_force_inter_sel	:	string	:=	"false";
		pll_dprio_fpll_vreg1_boost	:	string	:=	"fpll_vreg1_no_voltage_boost";
		pll_dprio_fpll_vreg_boost	:	string	:=	"fpll_vreg_no_voltage_boost";
		pll_dprio_power_iso_en	:	string	:=	"true";
		pll_dprio_status_select	:	string	:=	"dprio_normal_status";
		pll_dsm_ecn_bypass	:	string	:=	"false";
		pll_dsm_ecn_test_en	:	string	:=	"false";
		pll_dsm_fractional_division	:	string	:=	"00000000000000000000000000000000";
		pll_dsm_fractional_value_ready	:	string	:=	"pll_k_ready";
		pll_dsm_mode	:	string	:=	"dsm_mode_integer";
		pll_dsm_out_sel	:	string	:=	"pll_dsm_disable";
		pll_enable	:	string	:=	"false";
		pll_extra_csr	:	integer	:=	0;
		pll_fbclk_mux_1	:	string	:=	"pll_fbclk_mux_1_glb";
		pll_fbclk_mux_2	:	string	:=	"pll_fbclk_mux_2_fb_1";
		pll_iqclk_mux_sel	:	string	:=	"power_down";
		pll_l_counter	:	integer	:=	1;
		pll_l_counter_bypass	:	string	:=	"false";
		pll_l_counter_enable	:	string	:=	"true";
		pll_lf_cbig	:	string	:=	"lf_cbig_setting0";
		pll_lf_resistance	:	string	:=	"lf_res_setting0";
		pll_lf_ripplecap	:	string	:=	"lf_ripple_enabled_0";
		pll_lock_fltr_cfg	:	integer	:=	1;
		pll_lock_fltr_test	:	string	:=	"pll_lock_fltr_nrm";
		pll_lpf_rstn_value	:	string	:=	"lpf_normal";
		pll_m_counter	:	integer	:=	1;
		pll_m_counter_coarse_dly	:	string	:=	"0 ps";
		pll_m_counter_fine_dly	:	string	:=	"0 ps";
		pll_m_counter_in_src	:	string	:=	"m_cnt_in_src_test_clk";
		pll_m_counter_min_tco_enable	:	string	:=	"true";
		pll_m_counter_ph_mux_prst	:	integer	:=	0;
		pll_m_counter_prst	:	integer	:=	1;
		pll_n_counter	:	integer	:=	1;
		pll_n_counter_coarse_dly	:	string	:=	"0 ps";
		pll_n_counter_fine_dly	:	string	:=	"0 ps";
		pll_nreset_invert	:	string	:=	"false";
		pll_op_mode	:	string	:=	"false";
		pll_optimal	:	string	:=	"true";
		pll_powerdown_mode	:	string	:=	"false";
		pll_ppm_clk0_src	:	string	:=	"ppm_clk0_vss";
		pll_ppm_clk1_src	:	string	:=	"ppm_clk1_vss";
		pll_ref_buf_dly	:	string	:=	"0 ps";
		pll_rstn_override	:	string	:=	"false";
		pll_self_reset	:	string	:=	"false";
		pll_sup_mode	:	string	:=	"user_mode";
		pll_tclk_mux_en	:	string	:=	"false";
		pll_tclk_sel	:	string	:=	"pll_tclk_m_src";
		pll_test_enable	:	string	:=	"false";
		pll_unlock_fltr_cfg	:	integer	:=	0;
		pll_vccr_pd_en	:	string	:=	"false";
		pll_vco_freq_band_0	:	string	:=	"pll_freq_band0";
		pll_vco_freq_band_0_dyn_high_bits	:	integer	:=	0;
		pll_vco_freq_band_0_dyn_low_bits	:	integer	:=	0;
		pll_vco_freq_band_0_fix	:	integer	:=	1;
		pll_vco_freq_band_0_fix_high	:	string	:=	"pll_vco_freq_band_0_fix_high_0";
		pll_vco_freq_band_1	:	string	:=	"pll_freq_band0_1";
		pll_vco_freq_band_1_dyn_high_bits	:	integer	:=	0;
		pll_vco_freq_band_1_dyn_low_bits	:	integer	:=	0;
		pll_vco_freq_band_1_fix	:	integer	:=	1;
		pll_vco_freq_band_1_fix_high	:	string	:=	"pll_vco_freq_band_1_fix_high_0";
		pll_vco_ph0_en	:	string	:=	"false";
		pll_vco_ph0_value	:	string	:=	"pll_vco_ph0_vss";
		pll_vco_ph1_en	:	string	:=	"false";
		pll_vco_ph1_value	:	string	:=	"pll_vco_ph1_vss";
		pll_vco_ph2_en	:	string	:=	"false";
		pll_vco_ph2_value	:	string	:=	"pll_vco_ph2_vss";
		pll_vco_ph3_en	:	string	:=	"false";
		pll_vco_ph3_value	:	string	:=	"pll_vco_ph3_vss";
		pm_speed_grade	:	string	:=	"e2";
		pma_width	:	integer	:=	8;
		power_mode	:	string	:=	"low_power";
		power_rail_et	:	integer	:=	0;
		primary_use	:	string	:=	"tx";
		prot_mode	:	string	:=	"basic_tx";
		reference_clock_frequency	:	string	:=	"0 ps";
		reference_clock_frequency_scratch	:	string	:=	"0 hz";
		set_fpll_input_freq_range	:	integer	:=	0;
		side	:	string	:=	"side_unknown";
		silicon_rev	:	string	:=	"20nm5es";
		top_or_bottom	:	string	:=	"tb_unknown";
		vco_freq	:	string	:=	"000000000000000000000000000000000001";
		vco_freq_hz	:	string	:=	"0 hz";
		vco_frequency	:	string	:=	"0 ps";
		xpm_cmu_fpll_core_cal_vco_count_length	:	string	:=	"sel_8b_count";
		xpm_cmu_fpll_core_fpll_refclk_source	:	string	:=	"normal_refclk";
		xpm_cmu_fpll_core_fpll_vco_div_by_2_sel	:	string	:=	"bypass_divide_by_2";
		xpm_cmu_fpll_core_pfd_delay_compensation	:	string	:=	"normal_delay";
		xpm_cmu_fpll_core_pfd_pulse_width	:	string	:=	"pulse_width_setting0";
		xpm_cmu_fpll_core_xpm_cpvco_fpll_xpm_chgpmplf_fpll_cp_current_boost	:	string	:=	"normal_setting"
	);
	port (
		-- Architecture ports
		clk0bad_in	:	in	std_logic	:=	'0';
		clk1bad_in	:	in	std_logic	:=	'0';
		cnt_sel	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		core_refclk	:	in	std_logic	:=	'0';
		csr_bufin	:	in	std_logic	:=	'0';
		csr_clk	:	in	std_logic	:=	'0';
		csr_en	:	in	std_logic	:=	'0';
		csr_en_dly	:	in	std_logic	:=	'0';
		csr_in	:	in	std_logic	:=	'0';
		avmmclk	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		dps_rst_n	:	in	std_logic	:=	'0';
		extswitch_buf	:	in	std_logic	:=	'0';
		fbclk_in	:	in	std_logic	:=	'0';
		fpll_ppm_clk	:	in	std_logic_vector(1 downto 0)	:=	"00";
		iqtxrxclk	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		lc_to_fpll_refclk	:	in	std_logic	:=	'0';
		mdio_dis	:	in	std_logic	:=	'0';
		nfrzdrv	:	in	std_logic	:=	'0';
		nrpi_freeze	:	in	std_logic	:=	'0';
		num_phase_shifts	:	in	std_logic_vector(2 downto 0)	:=	"000";
		pfden	:	in	std_logic	:=	'0';
		phase_en	:	in	std_logic	:=	'0';
		pllclksel	:	in	std_logic	:=	'0';
		pma_atpg_los_en_n	:	in	std_logic	:=	'0';
		pma_csr_test_dis	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		refclk	:	in	std_logic	:=	'0';
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		rst_n	:	in	std_logic	:=	'0';
		scan_mode_n	:	in	std_logic	:=	'0';
		scan_shift_n	:	in	std_logic	:=	'0';
		up_dn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		block_select	:	out	std_logic	:=	'0';
		clk0	:	out	std_logic	:=	'0';
		clk0bad	:	out	std_logic	:=	'0';
		clk180	:	out	std_logic	:=	'0';
		clk1bad	:	out	std_logic	:=	'0';
		clklow	:	out	std_logic	:=	'0';
		csr_bufout	:	out	std_logic	:=	'0';
		csr_out	:	out	std_logic	:=	'0';
		fbclk_out	:	out	std_logic	:=	'0';
		clk_sel_override	:	out	std_logic	:=	'0';
		clk_sel_override_value	:	out	std_logic	:=	'0';
		fref	:	out	std_logic	:=	'0';
		hclk_out	:	out	std_logic	:=	'0';
		iqtxrxclk_out	:	out	std_logic	:=	'0';
		lock	:	out	std_logic	:=	'0';
		phase_done	:	out	std_logic	:=	'0';
		pll_cascade_out	:	out	std_logic	:=	'0';
		outclk	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		ppm_clk	:	out	std_logic_vector(1 downto 0)	:=	"00";
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000"
	);
end component;

begin



inst : twentynm_cmu_fpll_encrypted
	generic map (
		-- Instance parameters
		analog_mode	=>	analog_mode,
		bandwidth_range_high	=>	bandwidth_range_high,
		bandwidth_range_low	=>	bandwidth_range_low,
		bonding	=>	bonding,
		bw_sel	=>	bw_sel,
		cgb_div	=>	cgb_div,
		compensation_mode	=>	compensation_mode,
		datarate	=>	datarate,
		duty_cycle_0	=>	duty_cycle_0,
		duty_cycle_1	=>	duty_cycle_1,
		duty_cycle_2	=>	duty_cycle_2,
		duty_cycle_3	=>	duty_cycle_3,
		enable_idle_fpll_support	=>	enable_idle_fpll_support,
		f_max_band_0	=>	f_max_band_0,
		f_max_band_1	=>	f_max_band_1,
		f_max_band_2	=>	f_max_band_2,
		f_max_band_3	=>	f_max_band_3,
		f_max_band_4	=>	f_max_band_4,
		f_max_band_5	=>	f_max_band_5,
		f_max_band_6	=>	f_max_band_6,
		f_max_band_7	=>	f_max_band_7,
		f_max_band_8	=>	f_max_band_8,
		f_max_band_9	=>	f_max_band_9,
		f_max_div_two_bypass	=>	f_max_div_two_bypass,
		f_max_pfd	=>	f_max_pfd,
		f_max_pfd_bonded	=>	f_max_pfd_bonded,
		f_max_pfd_fractional	=>	f_max_pfd_fractional,
		f_max_pfd_integer	=>	f_max_pfd_integer,
		f_max_vco	=>	f_max_vco,
		f_max_vco_fractional	=>	f_max_vco_fractional,
		f_min_band_0	=>	f_min_band_0,
		f_min_band_1	=>	f_min_band_1,
		f_min_band_2	=>	f_min_band_2,
		f_min_band_3	=>	f_min_band_3,
		f_min_band_4	=>	f_min_band_4,
		f_min_band_5	=>	f_min_band_5,
		f_min_band_6	=>	f_min_band_6,
		f_min_band_7	=>	f_min_band_7,
		f_min_band_8	=>	f_min_band_8,
		f_min_band_9	=>	f_min_band_9,
		f_min_pfd	=>	f_min_pfd,
		f_min_vco	=>	f_min_vco,
		f_out_c0	=>	f_out_c0,
		f_out_c0_hz	=>	f_out_c0_hz,
		f_out_c1	=>	f_out_c1,
		f_out_c1_hz	=>	f_out_c1_hz,
		f_out_c2	=>	f_out_c2,
		f_out_c2_hz	=>	f_out_c2_hz,
		f_out_c3	=>	f_out_c3,
		f_out_c3_hz	=>	f_out_c3_hz,
		feedback	=>	feedback,
		fpll_cal_test_sel	=>	fpll_cal_test_sel,
		fpll_cas_out_enable	=>	fpll_cas_out_enable,
		fpll_hclk_out_enable	=>	fpll_hclk_out_enable,
		fpll_iqtxrxclk_out_enable	=>	fpll_iqtxrxclk_out_enable,
		hssi_output_clock_frequency	=>	hssi_output_clock_frequency,
		initial_settings	=>	initial_settings,
		input_tolerance	=>	input_tolerance_int,
		is_cascaded_pll	=>	is_cascaded_pll,
		is_otn	=>	is_otn,
		is_pa_core	=>	is_pa_core,
		is_sdi	=>	is_sdi,
		l_counter	=>	l_counter_int,
		m_counter	=>	m_counter_int,
		m_counter_c0	=>	m_counter_c0_int,
		m_counter_c1	=>	m_counter_c1_int,
		m_counter_c2	=>	m_counter_c2_int,
		m_counter_c3	=>	m_counter_c3_int,
		max_fractional_percentage	=>	max_fractional_percentage_int,
		min_fractional_percentage	=>	min_fractional_percentage_int,
		n_counter	=>	n_counter_int,
		out_freq	=>	out_freq,
		out_freq_hz	=>	out_freq_hz,
		output_clock_frequency_0	=>	output_clock_frequency_0,
		output_clock_frequency_1	=>	output_clock_frequency_1,
		output_clock_frequency_2	=>	output_clock_frequency_2,
		output_clock_frequency_3	=>	output_clock_frequency_3,
		output_tolerance	=>	output_tolerance_int,
		pfd_freq	=>	pfd_freq,
		phase_shift_0	=>	phase_shift_0,
		phase_shift_1	=>	phase_shift_1,
		phase_shift_2	=>	phase_shift_2,
		phase_shift_3	=>	phase_shift_3,
		pll_atb	=>	pll_atb,
		pll_bw_mode	=>	pll_bw_mode,
		pll_c0_pllcout_enable	=>	pll_c0_pllcout_enable,
		pll_c1_pllcout_enable	=>	pll_c1_pllcout_enable,
		pll_c2_pllcout_enable	=>	pll_c2_pllcout_enable,
		pll_c3_pllcout_enable	=>	pll_c3_pllcout_enable,
		pll_c_counter_0	=>	pll_c_counter_0,
		pll_c_counter_0_coarse_dly	=>	pll_c_counter_0_coarse_dly,
		pll_c_counter_0_fine_dly	=>	pll_c_counter_0_fine_dly,
		pll_c_counter_0_in_src	=>	pll_c_counter_0_in_src,
		pll_c_counter_0_min_tco_enable	=>	pll_c_counter_0_min_tco_enable,
		pll_c_counter_0_ph_mux_prst	=>	pll_c_counter_0_ph_mux_prst,
		pll_c_counter_0_prst	=>	pll_c_counter_0_prst,
		pll_c_counter_1	=>	pll_c_counter_1,
		pll_c_counter_1_coarse_dly	=>	pll_c_counter_1_coarse_dly,
		pll_c_counter_1_fine_dly	=>	pll_c_counter_1_fine_dly,
		pll_c_counter_1_in_src	=>	pll_c_counter_1_in_src,
		pll_c_counter_1_min_tco_enable	=>	pll_c_counter_1_min_tco_enable,
		pll_c_counter_1_ph_mux_prst	=>	pll_c_counter_1_ph_mux_prst,
		pll_c_counter_1_prst	=>	pll_c_counter_1_prst,
		pll_c_counter_2	=>	pll_c_counter_2,
		pll_c_counter_2_coarse_dly	=>	pll_c_counter_2_coarse_dly,
		pll_c_counter_2_fine_dly	=>	pll_c_counter_2_fine_dly,
		pll_c_counter_2_in_src	=>	pll_c_counter_2_in_src,
		pll_c_counter_2_min_tco_enable	=>	pll_c_counter_2_min_tco_enable,
		pll_c_counter_2_ph_mux_prst	=>	pll_c_counter_2_ph_mux_prst,
		pll_c_counter_2_prst	=>	pll_c_counter_2_prst,
		pll_c_counter_3	=>	pll_c_counter_3,
		pll_c_counter_3_coarse_dly	=>	pll_c_counter_3_coarse_dly,
		pll_c_counter_3_fine_dly	=>	pll_c_counter_3_fine_dly,
		pll_c_counter_3_in_src	=>	pll_c_counter_3_in_src,
		pll_c_counter_3_min_tco_enable	=>	pll_c_counter_3_min_tco_enable,
		pll_c_counter_3_ph_mux_prst	=>	pll_c_counter_3_ph_mux_prst,
		pll_c_counter_3_prst	=>	pll_c_counter_3_prst,
		pll_cal_status	=>	pll_cal_status,
		pll_calibration	=>	pll_calibration,
		pll_cmp_buf_dly	=>	pll_cmp_buf_dly,
		pll_cmu_rstn_value	=>	pll_cmu_rstn_value,
		pll_core_cali_ref_off	=>	pll_core_cali_ref_off,
		pll_core_cali_vco_off	=>	pll_core_cali_vco_off,
		pll_core_vccdreg_fb	=>	pll_core_vccdreg_fb,
		pll_core_vccdreg_fw	=>	pll_core_vccdreg_fw,
		pll_core_vreg0_atbsel	=>	pll_core_vreg0_atbsel,
		pll_core_vreg1_atbsel	=>	pll_core_vreg1_atbsel,
		pll_cp_compensation	=>	pll_cp_compensation,
		pll_cp_current_setting	=>	pll_cp_current_setting,
		pll_cp_lf_3rd_pole_freq	=>	pll_cp_lf_3rd_pole_freq,
		pll_cp_lf_order	=>	pll_cp_lf_order,
		pll_cp_testmode	=>	pll_cp_testmode,
		pll_ctrl_override_setting	=>	pll_ctrl_override_setting,
		pll_ctrl_plniotri_override	=>	pll_ctrl_plniotri_override,
		pll_device_variant	=>	pll_device_variant,
		pll_dprio_base_addr	=>	pll_dprio_base_addr,
		pll_dprio_broadcast_en	=>	pll_dprio_broadcast_en,
		pll_dprio_clk_vreg_boost	=>	pll_dprio_clk_vreg_boost,
		pll_dprio_cvp_inter_sel	=>	pll_dprio_cvp_inter_sel,
		pll_dprio_force_inter_sel	=>	pll_dprio_force_inter_sel,
		pll_dprio_fpll_vreg1_boost	=>	pll_dprio_fpll_vreg1_boost,
		pll_dprio_fpll_vreg_boost	=>	pll_dprio_fpll_vreg_boost,
		pll_dprio_power_iso_en	=>	pll_dprio_power_iso_en,
		pll_dprio_status_select	=>	pll_dprio_status_select,
		pll_dsm_ecn_bypass	=>	pll_dsm_ecn_bypass,
		pll_dsm_ecn_test_en	=>	pll_dsm_ecn_test_en,
		pll_dsm_fractional_division	=>	pll_dsm_fractional_division,
		pll_dsm_fractional_value_ready	=>	pll_dsm_fractional_value_ready,
		pll_dsm_mode	=>	pll_dsm_mode,
		pll_dsm_out_sel	=>	pll_dsm_out_sel,
		pll_enable	=>	pll_enable,
		pll_extra_csr	=>	pll_extra_csr,
		pll_fbclk_mux_1	=>	pll_fbclk_mux_1,
		pll_fbclk_mux_2	=>	pll_fbclk_mux_2,
		pll_iqclk_mux_sel	=>	pll_iqclk_mux_sel,
		pll_l_counter	=>	pll_l_counter,
		pll_l_counter_bypass	=>	pll_l_counter_bypass,
		pll_l_counter_enable	=>	pll_l_counter_enable,
		pll_lf_cbig	=>	pll_lf_cbig,
		pll_lf_resistance	=>	pll_lf_resistance,
		pll_lf_ripplecap	=>	pll_lf_ripplecap,
		pll_lock_fltr_cfg	=>	pll_lock_fltr_cfg,
		pll_lock_fltr_test	=>	pll_lock_fltr_test,
		pll_lpf_rstn_value	=>	pll_lpf_rstn_value,
		pll_m_counter	=>	pll_m_counter,
		pll_m_counter_coarse_dly	=>	pll_m_counter_coarse_dly,
		pll_m_counter_fine_dly	=>	pll_m_counter_fine_dly,
		pll_m_counter_in_src	=>	pll_m_counter_in_src,
		pll_m_counter_min_tco_enable	=>	pll_m_counter_min_tco_enable,
		pll_m_counter_ph_mux_prst	=>	pll_m_counter_ph_mux_prst,
		pll_m_counter_prst	=>	pll_m_counter_prst,
		pll_n_counter	=>	pll_n_counter,
		pll_n_counter_coarse_dly	=>	pll_n_counter_coarse_dly,
		pll_n_counter_fine_dly	=>	pll_n_counter_fine_dly,
		pll_nreset_invert	=>	pll_nreset_invert,
		pll_op_mode	=>	pll_op_mode,
		pll_optimal	=>	pll_optimal,
		pll_powerdown_mode	=>	pll_powerdown_mode,
		pll_ppm_clk0_src	=>	pll_ppm_clk0_src,
		pll_ppm_clk1_src	=>	pll_ppm_clk1_src,
		pll_ref_buf_dly	=>	pll_ref_buf_dly,
		pll_rstn_override	=>	pll_rstn_override,
		pll_self_reset	=>	pll_self_reset,
		pll_sup_mode	=>	pll_sup_mode,
		pll_tclk_mux_en	=>	pll_tclk_mux_en,
		pll_tclk_sel	=>	pll_tclk_sel,
		pll_test_enable	=>	pll_test_enable,
		pll_unlock_fltr_cfg	=>	pll_unlock_fltr_cfg,
		pll_vccr_pd_en	=>	pll_vccr_pd_en,
		pll_vco_freq_band_0	=>	pll_vco_freq_band_0,
		pll_vco_freq_band_0_dyn_high_bits	=>	pll_vco_freq_band_0_dyn_high_bits_int,
		pll_vco_freq_band_0_dyn_low_bits	=>	pll_vco_freq_band_0_dyn_low_bits_int,
		pll_vco_freq_band_0_fix	=>	pll_vco_freq_band_0_fix_int,
		pll_vco_freq_band_0_fix_high	=>	pll_vco_freq_band_0_fix_high,
		pll_vco_freq_band_1	=>	pll_vco_freq_band_1,
		pll_vco_freq_band_1_dyn_high_bits	=>	pll_vco_freq_band_1_dyn_high_bits_int,
		pll_vco_freq_band_1_dyn_low_bits	=>	pll_vco_freq_band_1_dyn_low_bits_int,
		pll_vco_freq_band_1_fix	=>	pll_vco_freq_band_1_fix_int,
		pll_vco_freq_band_1_fix_high	=>	pll_vco_freq_band_1_fix_high,
		pll_vco_ph0_en	=>	pll_vco_ph0_en,
		pll_vco_ph0_value	=>	pll_vco_ph0_value,
		pll_vco_ph1_en	=>	pll_vco_ph1_en,
		pll_vco_ph1_value	=>	pll_vco_ph1_value,
		pll_vco_ph2_en	=>	pll_vco_ph2_en,
		pll_vco_ph2_value	=>	pll_vco_ph2_value,
		pll_vco_ph3_en	=>	pll_vco_ph3_en,
		pll_vco_ph3_value	=>	pll_vco_ph3_value,
		pm_speed_grade	=>	pm_speed_grade,
		pma_width	=>	pma_width,
		power_mode	=>	power_mode,
		power_rail_et	=>	power_rail_et,
		primary_use	=>	primary_use,
		prot_mode	=>	prot_mode,
		reference_clock_frequency	=>	reference_clock_frequency,
		reference_clock_frequency_scratch	=>	reference_clock_frequency_scratch,
		set_fpll_input_freq_range	=>	set_fpll_input_freq_range_int,
		side	=>	side,
		silicon_rev	=>	silicon_rev,
		top_or_bottom	=>	top_or_bottom,
		vco_freq	=>	vco_freq,
		vco_freq_hz	=>	vco_freq_hz,
		vco_frequency	=>	vco_frequency,
		xpm_cmu_fpll_core_cal_vco_count_length	=>	xpm_cmu_fpll_core_cal_vco_count_length,
		xpm_cmu_fpll_core_fpll_refclk_source	=>	xpm_cmu_fpll_core_fpll_refclk_source,
		xpm_cmu_fpll_core_fpll_vco_div_by_2_sel	=>	xpm_cmu_fpll_core_fpll_vco_div_by_2_sel,
		xpm_cmu_fpll_core_pfd_delay_compensation	=>	xpm_cmu_fpll_core_pfd_delay_compensation,
		xpm_cmu_fpll_core_pfd_pulse_width	=>	xpm_cmu_fpll_core_pfd_pulse_width,
		xpm_cmu_fpll_core_xpm_cpvco_fpll_xpm_chgpmplf_fpll_cp_current_boost	=>	xpm_cmu_fpll_core_xpm_cpvco_fpll_xpm_chgpmplf_fpll_cp_current_boost
	)
	port map (
		-- Instance ports
		clk0bad_in	=>	clk0bad_in,
		clk1bad_in	=>	clk1bad_in,
		cnt_sel	=>	cnt_sel,
		core_refclk	=>	core_refclk,
		csr_bufin	=>	csr_bufin,
		csr_clk	=>	csr_clk,
		csr_en	=>	csr_en,
		csr_en_dly	=>	csr_en_dly,
		csr_in	=>	csr_in,
		avmmclk	=>	avmmclk,
		avmmrstn	=>	avmmrstn,
		dps_rst_n	=>	dps_rst_n,
		extswitch_buf	=>	extswitch_buf,
		fbclk_in	=>	fbclk_in,
		fpll_ppm_clk	=>	fpll_ppm_clk,
		iqtxrxclk	=>	iqtxrxclk,
		lc_to_fpll_refclk	=>	lc_to_fpll_refclk,
		mdio_dis	=>	mdio_dis,
		nfrzdrv	=>	nfrzdrv,
		nrpi_freeze	=>	nrpi_freeze,
		num_phase_shifts	=>	num_phase_shifts,
		pfden	=>	pfden,
		phase_en	=>	phase_en,
		pllclksel	=>	pllclksel,
		pma_atpg_los_en_n	=>	pma_atpg_los_en_n,
		pma_csr_test_dis	=>	pma_csr_test_dis,
		avmmread	=>	avmmread,
		refclk	=>	refclk,
		avmmaddress	=>	avmmaddress,
		rst_n	=>	rst_n,
		scan_mode_n	=>	scan_mode_n,
		scan_shift_n	=>	scan_shift_n,
		up_dn	=>	up_dn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		block_select	=>	block_select,
		clk0	=>	clk0,
		clk0bad	=>	clk0bad,
		clk180	=>	clk180,
		clk1bad	=>	clk1bad,
		clklow	=>	clklow,
		csr_bufout	=>	csr_bufout,
		csr_out	=>	csr_out,
		fbclk_out	=>	fbclk_out,
		clk_sel_override	=>	clk_sel_override,
		clk_sel_override_value	=>	clk_sel_override_value,
		fref	=>	fref,
		hclk_out	=>	hclk_out,
		iqtxrxclk_out	=>	iqtxrxclk_out,
		lock	=>	lock,
		phase_done	=>	phase_done,
		pll_cascade_out	=>	pll_cascade_out,
		outclk	=>	outclk,
		ppm_clk	=>	ppm_clk,
		avmmreaddata	=>	avmmreaddata
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_10g_rx_pcs	is
	generic (
		-- Entity parameters
		advanced_user_mode	:	string	:=	"disable";
		align_del	:	string	:=	"align_del_en";
		ber_bit_err_total_cnt	:	string	:=	"bit_err_total_cnt_10g";
		ber_clken	:	string	:=	"ber_clk_dis";
		ber_xus_timer_window	:	bit_vector	:=	B"000000100110001001010";
		bitslip_mode	:	string	:=	"bitslip_dis";
		blksync_bitslip_type	:	string	:=	"bitslip_comb";
		blksync_bitslip_wait_cnt	:	bit_vector	:=	B"001";
		blksync_bitslip_wait_type	:	string	:=	"bitslip_match";
		blksync_bypass	:	string	:=	"blksync_bypass_dis";
		blksync_clken	:	string	:=	"blksync_clk_dis";
		blksync_enum_invalid_sh_cnt	:	string	:=	"enum_invalid_sh_cnt_10g";
		blksync_knum_sh_cnt_postlock	:	string	:=	"knum_sh_cnt_postlock_10g";
		blksync_knum_sh_cnt_prelock	:	string	:=	"knum_sh_cnt_prelock_10g";
		blksync_pipeln	:	string	:=	"blksync_pipeln_dis";
		clr_errblk_cnt_en	:	string	:=	"disable";
		control_del	:	string	:=	"control_del_all";
		crcchk_bypass	:	string	:=	"crcchk_bypass_dis";
		crcchk_clken	:	string	:=	"crcchk_clk_dis";
		crcchk_inv	:	string	:=	"crcchk_inv_dis";
		crcchk_pipeln	:	string	:=	"crcchk_pipeln_dis";
		crcflag_pipeln	:	string	:=	"crcflag_pipeln_dis";
		ctrl_bit_reverse	:	string	:=	"ctrl_bit_reverse_dis";
		data_bit_reverse	:	string	:=	"data_bit_reverse_dis";
		dec64b66b_clken	:	string	:=	"dec64b66b_clk_dis";
		dec_64b66b_rxsm_bypass	:	string	:=	"dec_64b66b_rxsm_bypass_dis";
		descrm_bypass	:	string	:=	"descrm_bypass_en";
		descrm_clken	:	string	:=	"descrm_clk_dis";
		descrm_mode	:	string	:=	"async";
		descrm_pipeln	:	string	:=	"enable";
		dft_clk_out_sel	:	string	:=	"rx_master_clk";
		dis_signal_ok	:	string	:=	"dis_signal_ok_dis";
		dispchk_bypass	:	string	:=	"dispchk_bypass_dis";
		empty_flag_type	:	string	:=	"empty_rd_side";
		fast_path	:	string	:=	"fast_path_dis";
		fec_clken	:	string	:=	"fec_clk_dis";
		fec_enable	:	string	:=	"fec_dis";
		fifo_double_read	:	string	:=	"fifo_double_read_dis";
		fifo_stop_rd	:	string	:=	"n_rd_empty";
		fifo_stop_wr	:	string	:=	"n_wr_full";
		force_align	:	string	:=	"force_align_dis";
		frmsync_bypass	:	string	:=	"frmsync_bypass_dis";
		frmsync_clken	:	string	:=	"frmsync_clk_dis";
		frmsync_enum_scrm	:	string	:=	"enum_scrm_default";
		frmsync_enum_sync	:	string	:=	"enum_sync_default";
		frmsync_flag_type	:	string	:=	"all_framing_words";
		frmsync_knum_sync	:	string	:=	"knum_sync_default";
		frmsync_mfrm_length	:	bit_vector	:=	B"0000100000000000";
		frmsync_pipeln	:	string	:=	"frmsync_pipeln_dis";
		full_flag_type	:	string	:=	"full_wr_side";
		gb_rx_idwidth	:	string	:=	"width_32";
		gb_rx_odwidth	:	string	:=	"width_66";
		gbexp_clken	:	string	:=	"gbexp_clk_dis";
		low_latency_en	:	string	:=	"enable";
		lpbk_mode	:	string	:=	"lpbk_dis";
		master_clk_sel	:	string	:=	"master_rx_pma_clk";
		pempty_flag_type	:	string	:=	"pempty_rd_side";
		pfull_flag_type	:	string	:=	"pfull_wr_side";
		phcomp_rd_del	:	string	:=	"phcomp_rd_del2";
		pld_if_type	:	string	:=	"fifo";
		prot_mode	:	string	:=	"disable_mode";
		rand_clken	:	string	:=	"rand_clk_dis";
		rd_clk_sel	:	string	:=	"rd_rx_pma_clk";
		rdfifo_clken	:	string	:=	"rdfifo_clk_dis";
		reconfig_settings	:	string	:=	"{}";
		rx_fifo_write_ctrl	:	string	:=	"blklock_stops";
		rx_scrm_width	:	string	:=	"bit64";
		rx_sh_location	:	string	:=	"lsb";
		rx_signal_ok_sel	:	string	:=	"synchronized_ver";
		rx_sm_bypass	:	string	:=	"rx_sm_bypass_dis";
		rx_sm_hiber	:	string	:=	"rx_sm_hiber_en";
		rx_sm_pipeln	:	string	:=	"rx_sm_pipeln_dis";
		rx_testbus_sel	:	string	:=	"crc32_chk_testbus1";
		rx_true_b2b	:	string	:=	"b2b";
		rxfifo_empty	:	string	:=	"empty_default";
		rxfifo_full	:	string	:=	"full_default";
		rxfifo_mode	:	string	:=	"phase_comp";
		rxfifo_pempty	:	bit_vector	:=	B"00010";
		rxfifo_pfull	:	bit_vector	:=	B"10111";
		silicon_rev	:	string	:=	"20nm5es";
		stretch_num_stages	:	string	:=	"zero_stage";
		sup_mode	:	string	:=	"user_mode";
		test_mode	:	string	:=	"test_off";
		wrfifo_clken	:	string	:=	"wrfifo_clk_dis"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		krfec_refclk_dig	:	in	std_logic	:=	'0';
		r_rx_diag_word	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		r_rx_scrm_word	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		r_rx_skip_word	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		r_rx_sync_word	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		refclk_dig	:	in	std_logic	:=	'0';
		rx_align_clr	:	in	std_logic	:=	'0';
		rx_bitslip	:	in	std_logic	:=	'0';
		rx_clr_ber_count	:	in	std_logic	:=	'0';
		rx_clr_errblk_cnt	:	in	std_logic	:=	'0';
		rx_control_fb	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		rx_control_in_krfec	:	in	std_logic_vector(9 downto 0)	:=	"0000000000";
		rx_data_fb	:	in	std_logic_vector(127 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		rx_data_in_krfec	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		rx_data_valid_fb	:	in	std_logic	:=	'0';
		rx_data_valid_in_krfec	:	in	std_logic	:=	'0';
		rx_fifo_rd_data	:	in	std_logic_vector(73 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000";
		rx_fifo_rd_data_dw	:	in	std_logic_vector(73 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000";
		rx_pld_clk	:	in	std_logic	:=	'0';
		rx_pld_rst_n	:	in	std_logic	:=	'0';
		rx_pma_clk	:	in	std_logic	:=	'0';
		rx_pma_data	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		rx_prbs_err_clr	:	in	std_logic	:=	'0';
		rx_rd_en	:	in	std_logic	:=	'0';
		scan_mode_n	:	in	std_logic	:=	'0';
		signal_ok	:	in	std_logic	:=	'0';
		signal_ok_krfec	:	in	std_logic	:=	'0';
		tx_pma_clk	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_blk_lock_10g_reg	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_blk_lock_10g_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_clr_errblk_cnt_reg	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_clr_errblk_cnt_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_diag_data_status_10g_reg	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_diag_data_status_10g_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_frame_10g_reg	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_frame_10g_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_pld_rst_n_fifo	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_pld_rst_n_reg	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_pld_rst_n_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_align_clr_fifo	:	out	std_logic	:=	'0';
		pld_10g_rx_align_clr_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_align_clr_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_align_val_fifo	:	out	std_logic	:=	'0';
		pld_10g_rx_align_val_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_align_val_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_clr_ber_count_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_clr_ber_count_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_crc32_err_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_crc32_err_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_data_valid_10g_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_data_valid_fifo	:	out	std_logic	:=	'0';
		pld_10g_rx_data_valid_pcsdirect_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_data_valid_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_empty_fifo	:	out	std_logic	:=	'0';
		pld_10g_rx_fifo_del_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_fifo_del_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_fifo_insert_fifo	:	out	std_logic	:=	'0';
		pld_10g_rx_fifo_num_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_fifo_num_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_frame_lock_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_frame_lock_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_hi_ber_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_hi_ber_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_oflw_err_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_oflw_err_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_pempty_fifo	:	out	std_logic	:=	'0';
		pld_10g_rx_pfull_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_pfull_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_rd_en_fifo	:	out	std_logic	:=	'0';
		pld_pcs_rx_clk_out_10g_txclk_wire	:	out	std_logic	:=	'0';
		pld_pcs_rx_clk_out_10g_wire	:	out	std_logic	:=	'0';
		pld_rx_control_10g_reg	:	out	std_logic	:=	'0';
		pld_rx_control_10g_txclk_reg	:	out	std_logic	:=	'0';
		pld_rx_data_10g_reg	:	out	std_logic	:=	'0';
		pld_rx_data_10g_txclk_reg	:	out	std_logic	:=	'0';
		pld_rx_prbs_err_10g_txclk_reg	:	out	std_logic	:=	'0';
		pld_rx_prbs_err_clr_10g_txclk_reg	:	out	std_logic	:=	'0';
		rx_align_val	:	out	std_logic	:=	'0';
		rx_blk_lock	:	out	std_logic	:=	'0';
		rx_clk_out	:	out	std_logic	:=	'0';
		rx_clk_out_pld_if	:	out	std_logic	:=	'0';
		rx_control	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		rx_crc32_err	:	out	std_logic	:=	'0';
		rx_data	:	out	std_logic_vector(127 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		rx_data_valid	:	out	std_logic	:=	'0';
		rx_dft_clk_out	:	out	std_logic	:=	'0';
		rx_diag_status	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rx_empty	:	out	std_logic	:=	'0';
		rx_fec_clk	:	out	std_logic	:=	'0';
		rx_fifo_del	:	out	std_logic	:=	'0';
		rx_fifo_insert	:	out	std_logic	:=	'0';
		rx_fifo_num	:	out	std_logic_vector(4 downto 0)	:=	"00000";
		rx_fifo_rd_ptr	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rx_fifo_rd_ptr2	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rx_fifo_wr_clk	:	out	std_logic	:=	'0';
		rx_fifo_wr_data	:	out	std_logic_vector(73 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000";
		rx_fifo_wr_en	:	out	std_logic	:=	'0';
		rx_fifo_wr_ptr	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rx_fifo_wr_rst_n	:	out	std_logic	:=	'0';
		rx_frame_lock	:	out	std_logic	:=	'0';
		rx_hi_ber	:	out	std_logic	:=	'0';
		rx_master_clk	:	out	std_logic	:=	'0';
		rx_master_clk_rst_n	:	out	std_logic	:=	'0';
		rx_oflw_err	:	out	std_logic	:=	'0';
		rx_pempty	:	out	std_logic	:=	'0';
		rx_pfull	:	out	std_logic	:=	'0';
		rx_random_err	:	out	std_logic	:=	'0';
		rx_rx_frame	:	out	std_logic	:=	'0';
		rx_test_data	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000"
	);
end twentynm_hssi_10g_rx_pcs;

architecture behavior of twentynm_hssi_10g_rx_pcs	is

constant ber_xus_timer_window_int	:	integer	:=	bin2int(ber_xus_timer_window);
constant blksync_bitslip_wait_cnt_int	:	integer	:=	bin2int(blksync_bitslip_wait_cnt);
constant frmsync_mfrm_length_int	:	integer	:=	bin2int(frmsync_mfrm_length);
constant rxfifo_pempty_int	:	integer	:=	bin2int(rxfifo_pempty);
constant rxfifo_pfull_int	:	integer	:=	bin2int(rxfifo_pfull);



component	twentynm_hssi_10g_rx_pcs_encrypted
	generic (
		-- Architecture parameters
		advanced_user_mode	:	string	:=	"disable";
		align_del	:	string	:=	"align_del_en";
		ber_bit_err_total_cnt	:	string	:=	"bit_err_total_cnt_10g";
		ber_clken	:	string	:=	"ber_clk_dis";
		ber_xus_timer_window	:	integer	:=	19530;
		bitslip_mode	:	string	:=	"bitslip_dis";
		blksync_bitslip_type	:	string	:=	"bitslip_comb";
		blksync_bitslip_wait_cnt	:	integer	:=	1;
		blksync_bitslip_wait_type	:	string	:=	"bitslip_match";
		blksync_bypass	:	string	:=	"blksync_bypass_dis";
		blksync_clken	:	string	:=	"blksync_clk_dis";
		blksync_enum_invalid_sh_cnt	:	string	:=	"enum_invalid_sh_cnt_10g";
		blksync_knum_sh_cnt_postlock	:	string	:=	"knum_sh_cnt_postlock_10g";
		blksync_knum_sh_cnt_prelock	:	string	:=	"knum_sh_cnt_prelock_10g";
		blksync_pipeln	:	string	:=	"blksync_pipeln_dis";
		clr_errblk_cnt_en	:	string	:=	"disable";
		control_del	:	string	:=	"control_del_all";
		crcchk_bypass	:	string	:=	"crcchk_bypass_dis";
		crcchk_clken	:	string	:=	"crcchk_clk_dis";
		crcchk_inv	:	string	:=	"crcchk_inv_dis";
		crcchk_pipeln	:	string	:=	"crcchk_pipeln_dis";
		crcflag_pipeln	:	string	:=	"crcflag_pipeln_dis";
		ctrl_bit_reverse	:	string	:=	"ctrl_bit_reverse_dis";
		data_bit_reverse	:	string	:=	"data_bit_reverse_dis";
		dec64b66b_clken	:	string	:=	"dec64b66b_clk_dis";
		dec_64b66b_rxsm_bypass	:	string	:=	"dec_64b66b_rxsm_bypass_dis";
		descrm_bypass	:	string	:=	"descrm_bypass_en";
		descrm_clken	:	string	:=	"descrm_clk_dis";
		descrm_mode	:	string	:=	"async";
		descrm_pipeln	:	string	:=	"enable";
		dft_clk_out_sel	:	string	:=	"rx_master_clk";
		dis_signal_ok	:	string	:=	"dis_signal_ok_dis";
		dispchk_bypass	:	string	:=	"dispchk_bypass_dis";
		empty_flag_type	:	string	:=	"empty_rd_side";
		fast_path	:	string	:=	"fast_path_dis";
		fec_clken	:	string	:=	"fec_clk_dis";
		fec_enable	:	string	:=	"fec_dis";
		fifo_double_read	:	string	:=	"fifo_double_read_dis";
		fifo_stop_rd	:	string	:=	"n_rd_empty";
		fifo_stop_wr	:	string	:=	"n_wr_full";
		force_align	:	string	:=	"force_align_dis";
		frmsync_bypass	:	string	:=	"frmsync_bypass_dis";
		frmsync_clken	:	string	:=	"frmsync_clk_dis";
		frmsync_enum_scrm	:	string	:=	"enum_scrm_default";
		frmsync_enum_sync	:	string	:=	"enum_sync_default";
		frmsync_flag_type	:	string	:=	"all_framing_words";
		frmsync_knum_sync	:	string	:=	"knum_sync_default";
		frmsync_mfrm_length	:	integer	:=	2048;
		frmsync_pipeln	:	string	:=	"frmsync_pipeln_dis";
		full_flag_type	:	string	:=	"full_wr_side";
		gb_rx_idwidth	:	string	:=	"width_32";
		gb_rx_odwidth	:	string	:=	"width_66";
		gbexp_clken	:	string	:=	"gbexp_clk_dis";
		low_latency_en	:	string	:=	"enable";
		lpbk_mode	:	string	:=	"lpbk_dis";
		master_clk_sel	:	string	:=	"master_rx_pma_clk";
		pempty_flag_type	:	string	:=	"pempty_rd_side";
		pfull_flag_type	:	string	:=	"pfull_wr_side";
		phcomp_rd_del	:	string	:=	"phcomp_rd_del2";
		pld_if_type	:	string	:=	"fifo";
		prot_mode	:	string	:=	"disable_mode";
		rand_clken	:	string	:=	"rand_clk_dis";
		rd_clk_sel	:	string	:=	"rd_rx_pma_clk";
		rdfifo_clken	:	string	:=	"rdfifo_clk_dis";
		reconfig_settings	:	string	:=	"{}";
		rx_fifo_write_ctrl	:	string	:=	"blklock_stops";
		rx_scrm_width	:	string	:=	"bit64";
		rx_sh_location	:	string	:=	"lsb";
		rx_signal_ok_sel	:	string	:=	"synchronized_ver";
		rx_sm_bypass	:	string	:=	"rx_sm_bypass_dis";
		rx_sm_hiber	:	string	:=	"rx_sm_hiber_en";
		rx_sm_pipeln	:	string	:=	"rx_sm_pipeln_dis";
		rx_testbus_sel	:	string	:=	"crc32_chk_testbus1";
		rx_true_b2b	:	string	:=	"b2b";
		rxfifo_empty	:	string	:=	"empty_default";
		rxfifo_full	:	string	:=	"full_default";
		rxfifo_mode	:	string	:=	"phase_comp";
		rxfifo_pempty	:	integer	:=	2;
		rxfifo_pfull	:	integer	:=	23;
		silicon_rev	:	string	:=	"20nm5es";
		stretch_num_stages	:	string	:=	"zero_stage";
		sup_mode	:	string	:=	"user_mode";
		test_mode	:	string	:=	"test_off";
		wrfifo_clken	:	string	:=	"wrfifo_clk_dis"
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		krfec_refclk_dig	:	in	std_logic	:=	'0';
		r_rx_diag_word	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		r_rx_scrm_word	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		r_rx_skip_word	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		r_rx_sync_word	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		refclk_dig	:	in	std_logic	:=	'0';
		rx_align_clr	:	in	std_logic	:=	'0';
		rx_bitslip	:	in	std_logic	:=	'0';
		rx_clr_ber_count	:	in	std_logic	:=	'0';
		rx_clr_errblk_cnt	:	in	std_logic	:=	'0';
		rx_control_fb	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		rx_control_in_krfec	:	in	std_logic_vector(9 downto 0)	:=	"0000000000";
		rx_data_fb	:	in	std_logic_vector(127 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		rx_data_in_krfec	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		rx_data_valid_fb	:	in	std_logic	:=	'0';
		rx_data_valid_in_krfec	:	in	std_logic	:=	'0';
		rx_fifo_rd_data	:	in	std_logic_vector(73 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000";
		rx_fifo_rd_data_dw	:	in	std_logic_vector(73 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000";
		rx_pld_clk	:	in	std_logic	:=	'0';
		rx_pld_rst_n	:	in	std_logic	:=	'0';
		rx_pma_clk	:	in	std_logic	:=	'0';
		rx_pma_data	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		rx_prbs_err_clr	:	in	std_logic	:=	'0';
		rx_rd_en	:	in	std_logic	:=	'0';
		scan_mode_n	:	in	std_logic	:=	'0';
		signal_ok	:	in	std_logic	:=	'0';
		signal_ok_krfec	:	in	std_logic	:=	'0';
		tx_pma_clk	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_blk_lock_10g_reg	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_blk_lock_10g_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_clr_errblk_cnt_reg	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_clr_errblk_cnt_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_diag_data_status_10g_reg	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_diag_data_status_10g_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_frame_10g_reg	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_frame_10g_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_pld_rst_n_fifo	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_pld_rst_n_reg	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_pld_rst_n_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_align_clr_fifo	:	out	std_logic	:=	'0';
		pld_10g_rx_align_clr_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_align_clr_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_align_val_fifo	:	out	std_logic	:=	'0';
		pld_10g_rx_align_val_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_align_val_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_clr_ber_count_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_clr_ber_count_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_crc32_err_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_crc32_err_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_data_valid_10g_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_data_valid_fifo	:	out	std_logic	:=	'0';
		pld_10g_rx_data_valid_pcsdirect_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_data_valid_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_empty_fifo	:	out	std_logic	:=	'0';
		pld_10g_rx_fifo_del_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_fifo_del_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_fifo_insert_fifo	:	out	std_logic	:=	'0';
		pld_10g_rx_fifo_num_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_fifo_num_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_frame_lock_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_frame_lock_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_hi_ber_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_hi_ber_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_oflw_err_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_oflw_err_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_pempty_fifo	:	out	std_logic	:=	'0';
		pld_10g_rx_pfull_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_pfull_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_rx_rd_en_fifo	:	out	std_logic	:=	'0';
		pld_pcs_rx_clk_out_10g_txclk_wire	:	out	std_logic	:=	'0';
		pld_pcs_rx_clk_out_10g_wire	:	out	std_logic	:=	'0';
		pld_rx_control_10g_reg	:	out	std_logic	:=	'0';
		pld_rx_control_10g_txclk_reg	:	out	std_logic	:=	'0';
		pld_rx_data_10g_reg	:	out	std_logic	:=	'0';
		pld_rx_data_10g_txclk_reg	:	out	std_logic	:=	'0';
		pld_rx_prbs_err_10g_txclk_reg	:	out	std_logic	:=	'0';
		pld_rx_prbs_err_clr_10g_txclk_reg	:	out	std_logic	:=	'0';
		rx_align_val	:	out	std_logic	:=	'0';
		rx_blk_lock	:	out	std_logic	:=	'0';
		rx_clk_out	:	out	std_logic	:=	'0';
		rx_clk_out_pld_if	:	out	std_logic	:=	'0';
		rx_control	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		rx_crc32_err	:	out	std_logic	:=	'0';
		rx_data	:	out	std_logic_vector(127 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		rx_data_valid	:	out	std_logic	:=	'0';
		rx_dft_clk_out	:	out	std_logic	:=	'0';
		rx_diag_status	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rx_empty	:	out	std_logic	:=	'0';
		rx_fec_clk	:	out	std_logic	:=	'0';
		rx_fifo_del	:	out	std_logic	:=	'0';
		rx_fifo_insert	:	out	std_logic	:=	'0';
		rx_fifo_num	:	out	std_logic_vector(4 downto 0)	:=	"00000";
		rx_fifo_rd_ptr	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rx_fifo_rd_ptr2	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rx_fifo_wr_clk	:	out	std_logic	:=	'0';
		rx_fifo_wr_data	:	out	std_logic_vector(73 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000";
		rx_fifo_wr_en	:	out	std_logic	:=	'0';
		rx_fifo_wr_ptr	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rx_fifo_wr_rst_n	:	out	std_logic	:=	'0';
		rx_frame_lock	:	out	std_logic	:=	'0';
		rx_hi_ber	:	out	std_logic	:=	'0';
		rx_master_clk	:	out	std_logic	:=	'0';
		rx_master_clk_rst_n	:	out	std_logic	:=	'0';
		rx_oflw_err	:	out	std_logic	:=	'0';
		rx_pempty	:	out	std_logic	:=	'0';
		rx_pfull	:	out	std_logic	:=	'0';
		rx_random_err	:	out	std_logic	:=	'0';
		rx_rx_frame	:	out	std_logic	:=	'0';
		rx_test_data	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000"
	);
end component;

begin



inst : twentynm_hssi_10g_rx_pcs_encrypted
	generic map (
		-- Instance parameters
		advanced_user_mode	=>	advanced_user_mode,
		align_del	=>	align_del,
		ber_bit_err_total_cnt	=>	ber_bit_err_total_cnt,
		ber_clken	=>	ber_clken,
		ber_xus_timer_window	=>	ber_xus_timer_window_int,
		bitslip_mode	=>	bitslip_mode,
		blksync_bitslip_type	=>	blksync_bitslip_type,
		blksync_bitslip_wait_cnt	=>	blksync_bitslip_wait_cnt_int,
		blksync_bitslip_wait_type	=>	blksync_bitslip_wait_type,
		blksync_bypass	=>	blksync_bypass,
		blksync_clken	=>	blksync_clken,
		blksync_enum_invalid_sh_cnt	=>	blksync_enum_invalid_sh_cnt,
		blksync_knum_sh_cnt_postlock	=>	blksync_knum_sh_cnt_postlock,
		blksync_knum_sh_cnt_prelock	=>	blksync_knum_sh_cnt_prelock,
		blksync_pipeln	=>	blksync_pipeln,
		clr_errblk_cnt_en	=>	clr_errblk_cnt_en,
		control_del	=>	control_del,
		crcchk_bypass	=>	crcchk_bypass,
		crcchk_clken	=>	crcchk_clken,
		crcchk_inv	=>	crcchk_inv,
		crcchk_pipeln	=>	crcchk_pipeln,
		crcflag_pipeln	=>	crcflag_pipeln,
		ctrl_bit_reverse	=>	ctrl_bit_reverse,
		data_bit_reverse	=>	data_bit_reverse,
		dec64b66b_clken	=>	dec64b66b_clken,
		dec_64b66b_rxsm_bypass	=>	dec_64b66b_rxsm_bypass,
		descrm_bypass	=>	descrm_bypass,
		descrm_clken	=>	descrm_clken,
		descrm_mode	=>	descrm_mode,
		descrm_pipeln	=>	descrm_pipeln,
		dft_clk_out_sel	=>	dft_clk_out_sel,
		dis_signal_ok	=>	dis_signal_ok,
		dispchk_bypass	=>	dispchk_bypass,
		empty_flag_type	=>	empty_flag_type,
		fast_path	=>	fast_path,
		fec_clken	=>	fec_clken,
		fec_enable	=>	fec_enable,
		fifo_double_read	=>	fifo_double_read,
		fifo_stop_rd	=>	fifo_stop_rd,
		fifo_stop_wr	=>	fifo_stop_wr,
		force_align	=>	force_align,
		frmsync_bypass	=>	frmsync_bypass,
		frmsync_clken	=>	frmsync_clken,
		frmsync_enum_scrm	=>	frmsync_enum_scrm,
		frmsync_enum_sync	=>	frmsync_enum_sync,
		frmsync_flag_type	=>	frmsync_flag_type,
		frmsync_knum_sync	=>	frmsync_knum_sync,
		frmsync_mfrm_length	=>	frmsync_mfrm_length_int,
		frmsync_pipeln	=>	frmsync_pipeln,
		full_flag_type	=>	full_flag_type,
		gb_rx_idwidth	=>	gb_rx_idwidth,
		gb_rx_odwidth	=>	gb_rx_odwidth,
		gbexp_clken	=>	gbexp_clken,
		low_latency_en	=>	low_latency_en,
		lpbk_mode	=>	lpbk_mode,
		master_clk_sel	=>	master_clk_sel,
		pempty_flag_type	=>	pempty_flag_type,
		pfull_flag_type	=>	pfull_flag_type,
		phcomp_rd_del	=>	phcomp_rd_del,
		pld_if_type	=>	pld_if_type,
		prot_mode	=>	prot_mode,
		rand_clken	=>	rand_clken,
		rd_clk_sel	=>	rd_clk_sel,
		rdfifo_clken	=>	rdfifo_clken,
		reconfig_settings	=>	reconfig_settings,
		rx_fifo_write_ctrl	=>	rx_fifo_write_ctrl,
		rx_scrm_width	=>	rx_scrm_width,
		rx_sh_location	=>	rx_sh_location,
		rx_signal_ok_sel	=>	rx_signal_ok_sel,
		rx_sm_bypass	=>	rx_sm_bypass,
		rx_sm_hiber	=>	rx_sm_hiber,
		rx_sm_pipeln	=>	rx_sm_pipeln,
		rx_testbus_sel	=>	rx_testbus_sel,
		rx_true_b2b	=>	rx_true_b2b,
		rxfifo_empty	=>	rxfifo_empty,
		rxfifo_full	=>	rxfifo_full,
		rxfifo_mode	=>	rxfifo_mode,
		rxfifo_pempty	=>	rxfifo_pempty_int,
		rxfifo_pfull	=>	rxfifo_pfull_int,
		silicon_rev	=>	silicon_rev,
		stretch_num_stages	=>	stretch_num_stages,
		sup_mode	=>	sup_mode,
		test_mode	=>	test_mode,
		wrfifo_clken	=>	wrfifo_clken
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		krfec_refclk_dig	=>	krfec_refclk_dig,
		r_rx_diag_word	=>	r_rx_diag_word,
		r_rx_scrm_word	=>	r_rx_scrm_word,
		r_rx_skip_word	=>	r_rx_skip_word,
		r_rx_sync_word	=>	r_rx_sync_word,
		refclk_dig	=>	refclk_dig,
		rx_align_clr	=>	rx_align_clr,
		rx_bitslip	=>	rx_bitslip,
		rx_clr_ber_count	=>	rx_clr_ber_count,
		rx_clr_errblk_cnt	=>	rx_clr_errblk_cnt,
		rx_control_fb	=>	rx_control_fb,
		rx_control_in_krfec	=>	rx_control_in_krfec,
		rx_data_fb	=>	rx_data_fb,
		rx_data_in_krfec	=>	rx_data_in_krfec,
		rx_data_valid_fb	=>	rx_data_valid_fb,
		rx_data_valid_in_krfec	=>	rx_data_valid_in_krfec,
		rx_fifo_rd_data	=>	rx_fifo_rd_data,
		rx_fifo_rd_data_dw	=>	rx_fifo_rd_data_dw,
		rx_pld_clk	=>	rx_pld_clk,
		rx_pld_rst_n	=>	rx_pld_rst_n,
		rx_pma_clk	=>	rx_pma_clk,
		rx_pma_data	=>	rx_pma_data,
		rx_prbs_err_clr	=>	rx_prbs_err_clr,
		rx_rd_en	=>	rx_rd_en,
		scan_mode_n	=>	scan_mode_n,
		signal_ok	=>	signal_ok,
		signal_ok_krfec	=>	signal_ok_krfec,
		tx_pma_clk	=>	tx_pma_clk,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		pld_10g_krfec_rx_blk_lock_10g_reg	=>	pld_10g_krfec_rx_blk_lock_10g_reg,
		pld_10g_krfec_rx_blk_lock_10g_txclk_reg	=>	pld_10g_krfec_rx_blk_lock_10g_txclk_reg,
		pld_10g_krfec_rx_clr_errblk_cnt_reg	=>	pld_10g_krfec_rx_clr_errblk_cnt_reg,
		pld_10g_krfec_rx_clr_errblk_cnt_txclk_reg	=>	pld_10g_krfec_rx_clr_errblk_cnt_txclk_reg,
		pld_10g_krfec_rx_diag_data_status_10g_reg	=>	pld_10g_krfec_rx_diag_data_status_10g_reg,
		pld_10g_krfec_rx_diag_data_status_10g_txclk_reg	=>	pld_10g_krfec_rx_diag_data_status_10g_txclk_reg,
		pld_10g_krfec_rx_frame_10g_reg	=>	pld_10g_krfec_rx_frame_10g_reg,
		pld_10g_krfec_rx_frame_10g_txclk_reg	=>	pld_10g_krfec_rx_frame_10g_txclk_reg,
		pld_10g_krfec_rx_pld_rst_n_fifo	=>	pld_10g_krfec_rx_pld_rst_n_fifo,
		pld_10g_krfec_rx_pld_rst_n_reg	=>	pld_10g_krfec_rx_pld_rst_n_reg,
		pld_10g_krfec_rx_pld_rst_n_txclk_reg	=>	pld_10g_krfec_rx_pld_rst_n_txclk_reg,
		pld_10g_rx_align_clr_fifo	=>	pld_10g_rx_align_clr_fifo,
		pld_10g_rx_align_clr_reg	=>	pld_10g_rx_align_clr_reg,
		pld_10g_rx_align_clr_txclk_reg	=>	pld_10g_rx_align_clr_txclk_reg,
		pld_10g_rx_align_val_fifo	=>	pld_10g_rx_align_val_fifo,
		pld_10g_rx_align_val_reg	=>	pld_10g_rx_align_val_reg,
		pld_10g_rx_align_val_txclk_reg	=>	pld_10g_rx_align_val_txclk_reg,
		pld_10g_rx_clr_ber_count_reg	=>	pld_10g_rx_clr_ber_count_reg,
		pld_10g_rx_clr_ber_count_txclk_reg	=>	pld_10g_rx_clr_ber_count_txclk_reg,
		pld_10g_rx_crc32_err_reg	=>	pld_10g_rx_crc32_err_reg,
		pld_10g_rx_crc32_err_txclk_reg	=>	pld_10g_rx_crc32_err_txclk_reg,
		pld_10g_rx_data_valid_10g_reg	=>	pld_10g_rx_data_valid_10g_reg,
		pld_10g_rx_data_valid_fifo	=>	pld_10g_rx_data_valid_fifo,
		pld_10g_rx_data_valid_pcsdirect_reg	=>	pld_10g_rx_data_valid_pcsdirect_reg,
		pld_10g_rx_data_valid_txclk_reg	=>	pld_10g_rx_data_valid_txclk_reg,
		pld_10g_rx_empty_fifo	=>	pld_10g_rx_empty_fifo,
		pld_10g_rx_fifo_del_reg	=>	pld_10g_rx_fifo_del_reg,
		pld_10g_rx_fifo_del_txclk_reg	=>	pld_10g_rx_fifo_del_txclk_reg,
		pld_10g_rx_fifo_insert_fifo	=>	pld_10g_rx_fifo_insert_fifo,
		pld_10g_rx_fifo_num_reg	=>	pld_10g_rx_fifo_num_reg,
		pld_10g_rx_fifo_num_txclk_reg	=>	pld_10g_rx_fifo_num_txclk_reg,
		pld_10g_rx_frame_lock_reg	=>	pld_10g_rx_frame_lock_reg,
		pld_10g_rx_frame_lock_txclk_reg	=>	pld_10g_rx_frame_lock_txclk_reg,
		pld_10g_rx_hi_ber_reg	=>	pld_10g_rx_hi_ber_reg,
		pld_10g_rx_hi_ber_txclk_reg	=>	pld_10g_rx_hi_ber_txclk_reg,
		pld_10g_rx_oflw_err_reg	=>	pld_10g_rx_oflw_err_reg,
		pld_10g_rx_oflw_err_txclk_reg	=>	pld_10g_rx_oflw_err_txclk_reg,
		pld_10g_rx_pempty_fifo	=>	pld_10g_rx_pempty_fifo,
		pld_10g_rx_pfull_reg	=>	pld_10g_rx_pfull_reg,
		pld_10g_rx_pfull_txclk_reg	=>	pld_10g_rx_pfull_txclk_reg,
		pld_10g_rx_rd_en_fifo	=>	pld_10g_rx_rd_en_fifo,
		pld_pcs_rx_clk_out_10g_txclk_wire	=>	pld_pcs_rx_clk_out_10g_txclk_wire,
		pld_pcs_rx_clk_out_10g_wire	=>	pld_pcs_rx_clk_out_10g_wire,
		pld_rx_control_10g_reg	=>	pld_rx_control_10g_reg,
		pld_rx_control_10g_txclk_reg	=>	pld_rx_control_10g_txclk_reg,
		pld_rx_data_10g_reg	=>	pld_rx_data_10g_reg,
		pld_rx_data_10g_txclk_reg	=>	pld_rx_data_10g_txclk_reg,
		pld_rx_prbs_err_10g_txclk_reg	=>	pld_rx_prbs_err_10g_txclk_reg,
		pld_rx_prbs_err_clr_10g_txclk_reg	=>	pld_rx_prbs_err_clr_10g_txclk_reg,
		rx_align_val	=>	rx_align_val,
		rx_blk_lock	=>	rx_blk_lock,
		rx_clk_out	=>	rx_clk_out,
		rx_clk_out_pld_if	=>	rx_clk_out_pld_if,
		rx_control	=>	rx_control,
		rx_crc32_err	=>	rx_crc32_err,
		rx_data	=>	rx_data,
		rx_data_valid	=>	rx_data_valid,
		rx_dft_clk_out	=>	rx_dft_clk_out,
		rx_diag_status	=>	rx_diag_status,
		rx_empty	=>	rx_empty,
		rx_fec_clk	=>	rx_fec_clk,
		rx_fifo_del	=>	rx_fifo_del,
		rx_fifo_insert	=>	rx_fifo_insert,
		rx_fifo_num	=>	rx_fifo_num,
		rx_fifo_rd_ptr	=>	rx_fifo_rd_ptr,
		rx_fifo_rd_ptr2	=>	rx_fifo_rd_ptr2,
		rx_fifo_wr_clk	=>	rx_fifo_wr_clk,
		rx_fifo_wr_data	=>	rx_fifo_wr_data,
		rx_fifo_wr_en	=>	rx_fifo_wr_en,
		rx_fifo_wr_ptr	=>	rx_fifo_wr_ptr,
		rx_fifo_wr_rst_n	=>	rx_fifo_wr_rst_n,
		rx_frame_lock	=>	rx_frame_lock,
		rx_hi_ber	=>	rx_hi_ber,
		rx_master_clk	=>	rx_master_clk,
		rx_master_clk_rst_n	=>	rx_master_clk_rst_n,
		rx_oflw_err	=>	rx_oflw_err,
		rx_pempty	=>	rx_pempty,
		rx_pfull	=>	rx_pfull,
		rx_random_err	=>	rx_random_err,
		rx_rx_frame	=>	rx_rx_frame,
		rx_test_data	=>	rx_test_data
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_10g_tx_pcs	is
	generic (
		-- Entity parameters
		advanced_user_mode	:	string	:=	"disable";
		bitslip_en	:	string	:=	"bitslip_dis";
		bonding_dft_en	:	string	:=	"dft_dis";
		bonding_dft_val	:	string	:=	"dft_0";
		comp_cnt	:	bit_vector	:=	B"00000000";
		compin_sel	:	string	:=	"compin_master";
		crcgen_bypass	:	string	:=	"crcgen_bypass_dis";
		crcgen_clken	:	string	:=	"crcgen_clk_dis";
		crcgen_err	:	string	:=	"crcgen_err_dis";
		crcgen_inv	:	string	:=	"crcgen_inv_dis";
		ctrl_bit_reverse	:	string	:=	"ctrl_bit_reverse_dis";
		ctrl_plane_bonding	:	string	:=	"individual";
		data_bit_reverse	:	string	:=	"data_bit_reverse_dis";
		dft_clk_out_sel	:	string	:=	"tx_master_clk";
		dispgen_bypass	:	string	:=	"dispgen_bypass_dis";
		dispgen_clken	:	string	:=	"dispgen_clk_dis";
		dispgen_err	:	string	:=	"dispgen_err_dis";
		dispgen_pipeln	:	string	:=	"dispgen_pipeln_dis";
		distdwn_bypass_pipeln	:	string	:=	"distdwn_bypass_pipeln_dis";
		distdwn_master	:	string	:=	"distdwn_master_en";
		distup_bypass_pipeln	:	string	:=	"distup_bypass_pipeln_dis";
		distup_master	:	string	:=	"distup_master_en";
		dv_bond	:	string	:=	"dv_bond_dis";
		empty_flag_type	:	string	:=	"empty_rd_side";
		enc64b66b_txsm_clken	:	string	:=	"enc64b66b_txsm_clk_dis";
		enc_64b66b_txsm_bypass	:	string	:=	"enc_64b66b_txsm_bypass_dis";
		fastpath	:	string	:=	"fastpath_dis";
		fec_clken	:	string	:=	"fec_clk_dis";
		fec_enable	:	string	:=	"fec_dis";
		fifo_double_write	:	string	:=	"fifo_double_write_dis";
		fifo_reg_fast	:	string	:=	"fifo_reg_fast_dis";
		fifo_stop_rd	:	string	:=	"n_rd_empty";
		fifo_stop_wr	:	string	:=	"n_wr_full";
		frmgen_burst	:	string	:=	"frmgen_burst_dis";
		frmgen_bypass	:	string	:=	"frmgen_bypass_dis";
		frmgen_clken	:	string	:=	"frmgen_clk_dis";
		frmgen_mfrm_length	:	bit_vector	:=	B"0000100000000000";
		frmgen_pipeln	:	string	:=	"frmgen_pipeln_dis";
		frmgen_pyld_ins	:	string	:=	"frmgen_pyld_ins_dis";
		frmgen_wordslip	:	string	:=	"frmgen_wordslip_dis";
		full_flag_type	:	string	:=	"full_wr_side";
		gb_pipeln_bypass	:	string	:=	"enable";
		gb_tx_idwidth	:	string	:=	"width_50";
		gb_tx_odwidth	:	string	:=	"width_32";
		gbred_clken	:	string	:=	"gbred_clk_dis";
		indv	:	string	:=	"indv_en";
		low_latency_en	:	string	:=	"enable";
		master_clk_sel	:	string	:=	"master_tx_pma_clk";
		pempty_flag_type	:	string	:=	"pempty_rd_side";
		pfull_flag_type	:	string	:=	"pfull_wr_side";
		phcomp_rd_del	:	string	:=	"phcomp_rd_del2";
		pld_if_type	:	string	:=	"fifo";
		prot_mode	:	string	:=	"disable_mode";
		pseudo_random	:	string	:=	"all_0";
		pseudo_seed_a	:	string	:=	"1111111111111111111111111111111111111111111111111111111111";
		pseudo_seed_b	:	string	:=	"1111111111111111111111111111111111111111111111111111111111";
		random_disp	:	string	:=	"disable";
		rdfifo_clken	:	string	:=	"rdfifo_clk_dis";
		reconfig_settings	:	string	:=	"{}";
		scrm_bypass	:	string	:=	"scrm_bypass_dis";
		scrm_clken	:	string	:=	"scrm_clk_dis";
		scrm_mode	:	string	:=	"async";
		scrm_pipeln	:	string	:=	"enable";
		sh_err	:	string	:=	"sh_err_dis";
		silicon_rev	:	string	:=	"20nm5es";
		sop_mark	:	string	:=	"sop_mark_dis";
		stretch_num_stages	:	string	:=	"zero_stage";
		sup_mode	:	string	:=	"user_mode";
		test_mode	:	string	:=	"test_off";
		tx_scrm_err	:	string	:=	"scrm_err_dis";
		tx_scrm_width	:	string	:=	"bit64";
		tx_sh_location	:	string	:=	"lsb";
		tx_sm_bypass	:	string	:=	"tx_sm_bypass_dis";
		tx_sm_pipeln	:	string	:=	"tx_sm_pipeln_dis";
		tx_testbus_sel	:	string	:=	"crc32_gen_testbus1";
		txfifo_empty	:	string	:=	"empty_default";
		txfifo_full	:	string	:=	"full_default";
		txfifo_mode	:	string	:=	"phase_comp";
		txfifo_pempty	:	bit_vector	:=	B"0010";
		txfifo_pfull	:	bit_vector	:=	B"1011";
		wr_clk_sel	:	string	:=	"wr_tx_pma_clk";
		wrfifo_clken	:	string	:=	"wrfifo_clk_dis"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		distdwn_in_dv	:	in	std_logic	:=	'0';
		distdwn_in_rden	:	in	std_logic	:=	'0';
		distdwn_in_wren	:	in	std_logic	:=	'0';
		distup_in_dv	:	in	std_logic	:=	'0';
		distup_in_rden	:	in	std_logic	:=	'0';
		distup_in_wren	:	in	std_logic	:=	'0';
		krfec_refclk_dig	:	in	std_logic	:=	'0';
		r_tx_diag_word	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		r_tx_scrm_word	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		r_tx_skip_word	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		r_tx_sync_word	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		refclk_dig	:	in	std_logic	:=	'0';
		scan_mode_n	:	in	std_logic	:=	'0';
		tx_bitslip	:	in	std_logic_vector(6 downto 0)	:=	"0000000";
		tx_burst_en	:	in	std_logic	:=	'0';
		tx_control	:	in	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		tx_control_reg	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		tx_data	:	in	std_logic_vector(127 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		tx_data_in_krfec	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		tx_data_reg	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		tx_data_valid	:	in	std_logic	:=	'0';
		tx_data_valid_reg	:	in	std_logic	:=	'0';
		tx_diag_status	:	in	std_logic_vector(1 downto 0)	:=	"00";
		tx_fifo_rd_data	:	in	std_logic_vector(72 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000000000000";
		tx_pld_clk	:	in	std_logic	:=	'0';
		tx_pld_rst_n	:	in	std_logic	:=	'0';
		tx_pma_clk	:	in	std_logic	:=	'0';
		tx_wordslip	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		pld_10g_krfec_tx_frame_10g_reg	:	out	std_logic	:=	'0';
		pld_10g_krfec_tx_pld_rst_n_fifo	:	out	std_logic	:=	'0';
		pld_10g_krfec_tx_pld_rst_n_reg	:	out	std_logic	:=	'0';
		pld_10g_tx_bitslip_reg	:	out	std_logic	:=	'0';
		pld_10g_tx_burst_en_exe_reg	:	out	std_logic	:=	'0';
		pld_10g_tx_data_valid_10g_reg	:	out	std_logic	:=	'0';
		pld_10g_tx_data_valid_fifo	:	out	std_logic	:=	'0';
		pld_10g_tx_data_valid_reg	:	out	std_logic	:=	'0';
		pld_10g_tx_diag_status_reg	:	out	std_logic	:=	'0';
		pld_10g_tx_empty_reg	:	out	std_logic	:=	'0';
		pld_10g_tx_fifo_num_reg	:	out	std_logic	:=	'0';
		pld_10g_tx_full_fifo	:	out	std_logic	:=	'0';
		pld_10g_tx_full_reg	:	out	std_logic	:=	'0';
		pld_10g_tx_pempty_reg	:	out	std_logic	:=	'0';
		pld_10g_tx_pfull_fifo	:	out	std_logic	:=	'0';
		pld_10g_tx_wordslip_exe_reg	:	out	std_logic	:=	'0';
		pld_10g_tx_wordslip_reg	:	out	std_logic	:=	'0';
		pld_pcs_tx_clk_out_10g_wire	:	out	std_logic	:=	'0';
		pld_tx_burst_en_reg	:	out	std_logic	:=	'0';
		pld_tx_control_lo_10g_reg	:	out	std_logic	:=	'0';
		pld_tx_data_10g_fifo	:	out	std_logic	:=	'0';
		pld_tx_data_lo_10g_reg	:	out	std_logic	:=	'0';
		distdwn_out_dv	:	out	std_logic	:=	'0';
		distdwn_out_rden	:	out	std_logic	:=	'0';
		distdwn_out_wren	:	out	std_logic	:=	'0';
		distup_out_dv	:	out	std_logic	:=	'0';
		distup_out_rden	:	out	std_logic	:=	'0';
		distup_out_wren	:	out	std_logic	:=	'0';
		tx_burst_en_exe	:	out	std_logic	:=	'0';
		tx_clk_out	:	out	std_logic	:=	'0';
		tx_clk_out_pld_if	:	out	std_logic	:=	'0';
		tx_clk_out_pma_if	:	out	std_logic	:=	'0';
		tx_control_out_krfec	:	out	std_logic_vector(8 downto 0)	:=	"000000000";
		tx_data_out_krfec	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		tx_data_valid_out_krfec	:	out	std_logic	:=	'0';
		tx_dft_clk_out	:	out	std_logic	:=	'0';
		tx_empty	:	out	std_logic	:=	'0';
		tx_fec_clk	:	out	std_logic	:=	'0';
		tx_fifo_num	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		tx_fifo_rd_ptr	:	out	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		tx_fifo_wr_clk	:	out	std_logic	:=	'0';
		tx_fifo_wr_data	:	out	std_logic_vector(72 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000000000000";
		tx_fifo_wr_data_dw	:	out	std_logic_vector(72 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000000000000";
		tx_fifo_wr_en	:	out	std_logic	:=	'0';
		tx_fifo_wr_ptr	:	out	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		tx_fifo_wr_rst_n	:	out	std_logic	:=	'0';
		tx_frame	:	out	std_logic	:=	'0';
		tx_full	:	out	std_logic	:=	'0';
		tx_master_clk	:	out	std_logic	:=	'0';
		tx_master_clk_rst_n	:	out	std_logic	:=	'0';
		tx_pempty	:	out	std_logic	:=	'0';
		tx_pfull	:	out	std_logic	:=	'0';
		tx_pma_data	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		tx_pma_gating_val	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		tx_test_data	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		tx_wordslip_exe	:	out	std_logic	:=	'0'
	);
end twentynm_hssi_10g_tx_pcs;

architecture behavior of twentynm_hssi_10g_tx_pcs	is

constant comp_cnt_int	:	integer	:=	bin2int(comp_cnt);
constant frmgen_mfrm_length_int	:	integer	:=	bin2int(frmgen_mfrm_length);
constant txfifo_pempty_int	:	integer	:=	bin2int(txfifo_pempty);
constant txfifo_pfull_int	:	integer	:=	bin2int(txfifo_pfull);



component	twentynm_hssi_10g_tx_pcs_encrypted
	generic (
		-- Architecture parameters
		advanced_user_mode	:	string	:=	"disable";
		bitslip_en	:	string	:=	"bitslip_dis";
		bonding_dft_en	:	string	:=	"dft_dis";
		bonding_dft_val	:	string	:=	"dft_0";
		comp_cnt	:	integer	:=	0;
		compin_sel	:	string	:=	"compin_master";
		crcgen_bypass	:	string	:=	"crcgen_bypass_dis";
		crcgen_clken	:	string	:=	"crcgen_clk_dis";
		crcgen_err	:	string	:=	"crcgen_err_dis";
		crcgen_inv	:	string	:=	"crcgen_inv_dis";
		ctrl_bit_reverse	:	string	:=	"ctrl_bit_reverse_dis";
		ctrl_plane_bonding	:	string	:=	"individual";
		data_bit_reverse	:	string	:=	"data_bit_reverse_dis";
		dft_clk_out_sel	:	string	:=	"tx_master_clk";
		dispgen_bypass	:	string	:=	"dispgen_bypass_dis";
		dispgen_clken	:	string	:=	"dispgen_clk_dis";
		dispgen_err	:	string	:=	"dispgen_err_dis";
		dispgen_pipeln	:	string	:=	"dispgen_pipeln_dis";
		distdwn_bypass_pipeln	:	string	:=	"distdwn_bypass_pipeln_dis";
		distdwn_master	:	string	:=	"distdwn_master_en";
		distup_bypass_pipeln	:	string	:=	"distup_bypass_pipeln_dis";
		distup_master	:	string	:=	"distup_master_en";
		dv_bond	:	string	:=	"dv_bond_dis";
		empty_flag_type	:	string	:=	"empty_rd_side";
		enc64b66b_txsm_clken	:	string	:=	"enc64b66b_txsm_clk_dis";
		enc_64b66b_txsm_bypass	:	string	:=	"enc_64b66b_txsm_bypass_dis";
		fastpath	:	string	:=	"fastpath_dis";
		fec_clken	:	string	:=	"fec_clk_dis";
		fec_enable	:	string	:=	"fec_dis";
		fifo_double_write	:	string	:=	"fifo_double_write_dis";
		fifo_reg_fast	:	string	:=	"fifo_reg_fast_dis";
		fifo_stop_rd	:	string	:=	"n_rd_empty";
		fifo_stop_wr	:	string	:=	"n_wr_full";
		frmgen_burst	:	string	:=	"frmgen_burst_dis";
		frmgen_bypass	:	string	:=	"frmgen_bypass_dis";
		frmgen_clken	:	string	:=	"frmgen_clk_dis";
		frmgen_mfrm_length	:	integer	:=	2048;
		frmgen_pipeln	:	string	:=	"frmgen_pipeln_dis";
		frmgen_pyld_ins	:	string	:=	"frmgen_pyld_ins_dis";
		frmgen_wordslip	:	string	:=	"frmgen_wordslip_dis";
		full_flag_type	:	string	:=	"full_wr_side";
		gb_pipeln_bypass	:	string	:=	"enable";
		gb_tx_idwidth	:	string	:=	"width_50";
		gb_tx_odwidth	:	string	:=	"width_32";
		gbred_clken	:	string	:=	"gbred_clk_dis";
		indv	:	string	:=	"indv_en";
		low_latency_en	:	string	:=	"enable";
		master_clk_sel	:	string	:=	"master_tx_pma_clk";
		pempty_flag_type	:	string	:=	"pempty_rd_side";
		pfull_flag_type	:	string	:=	"pfull_wr_side";
		phcomp_rd_del	:	string	:=	"phcomp_rd_del2";
		pld_if_type	:	string	:=	"fifo";
		prot_mode	:	string	:=	"disable_mode";
		pseudo_random	:	string	:=	"all_0";
		pseudo_seed_a	:	string	:=	"1111111111111111111111111111111111111111111111111111111111";
		pseudo_seed_b	:	string	:=	"1111111111111111111111111111111111111111111111111111111111";
		random_disp	:	string	:=	"disable";
		rdfifo_clken	:	string	:=	"rdfifo_clk_dis";
		reconfig_settings	:	string	:=	"{}";
		scrm_bypass	:	string	:=	"scrm_bypass_dis";
		scrm_clken	:	string	:=	"scrm_clk_dis";
		scrm_mode	:	string	:=	"async";
		scrm_pipeln	:	string	:=	"enable";
		sh_err	:	string	:=	"sh_err_dis";
		silicon_rev	:	string	:=	"20nm5es";
		sop_mark	:	string	:=	"sop_mark_dis";
		stretch_num_stages	:	string	:=	"zero_stage";
		sup_mode	:	string	:=	"user_mode";
		test_mode	:	string	:=	"test_off";
		tx_scrm_err	:	string	:=	"scrm_err_dis";
		tx_scrm_width	:	string	:=	"bit64";
		tx_sh_location	:	string	:=	"lsb";
		tx_sm_bypass	:	string	:=	"tx_sm_bypass_dis";
		tx_sm_pipeln	:	string	:=	"tx_sm_pipeln_dis";
		tx_testbus_sel	:	string	:=	"crc32_gen_testbus1";
		txfifo_empty	:	string	:=	"empty_default";
		txfifo_full	:	string	:=	"full_default";
		txfifo_mode	:	string	:=	"phase_comp";
		txfifo_pempty	:	integer	:=	2;
		txfifo_pfull	:	integer	:=	11;
		wr_clk_sel	:	string	:=	"wr_tx_pma_clk";
		wrfifo_clken	:	string	:=	"wrfifo_clk_dis"
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		distdwn_in_dv	:	in	std_logic	:=	'0';
		distdwn_in_rden	:	in	std_logic	:=	'0';
		distdwn_in_wren	:	in	std_logic	:=	'0';
		distup_in_dv	:	in	std_logic	:=	'0';
		distup_in_rden	:	in	std_logic	:=	'0';
		distup_in_wren	:	in	std_logic	:=	'0';
		krfec_refclk_dig	:	in	std_logic	:=	'0';
		r_tx_diag_word	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		r_tx_scrm_word	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		r_tx_skip_word	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		r_tx_sync_word	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		refclk_dig	:	in	std_logic	:=	'0';
		scan_mode_n	:	in	std_logic	:=	'0';
		tx_bitslip	:	in	std_logic_vector(6 downto 0)	:=	"0000000";
		tx_burst_en	:	in	std_logic	:=	'0';
		tx_control	:	in	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		tx_control_reg	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		tx_data	:	in	std_logic_vector(127 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		tx_data_in_krfec	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		tx_data_reg	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		tx_data_valid	:	in	std_logic	:=	'0';
		tx_data_valid_reg	:	in	std_logic	:=	'0';
		tx_diag_status	:	in	std_logic_vector(1 downto 0)	:=	"00";
		tx_fifo_rd_data	:	in	std_logic_vector(72 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000000000000";
		tx_pld_clk	:	in	std_logic	:=	'0';
		tx_pld_rst_n	:	in	std_logic	:=	'0';
		tx_pma_clk	:	in	std_logic	:=	'0';
		tx_wordslip	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		pld_10g_krfec_tx_frame_10g_reg	:	out	std_logic	:=	'0';
		pld_10g_krfec_tx_pld_rst_n_fifo	:	out	std_logic	:=	'0';
		pld_10g_krfec_tx_pld_rst_n_reg	:	out	std_logic	:=	'0';
		pld_10g_tx_bitslip_reg	:	out	std_logic	:=	'0';
		pld_10g_tx_burst_en_exe_reg	:	out	std_logic	:=	'0';
		pld_10g_tx_data_valid_10g_reg	:	out	std_logic	:=	'0';
		pld_10g_tx_data_valid_fifo	:	out	std_logic	:=	'0';
		pld_10g_tx_data_valid_reg	:	out	std_logic	:=	'0';
		pld_10g_tx_diag_status_reg	:	out	std_logic	:=	'0';
		pld_10g_tx_empty_reg	:	out	std_logic	:=	'0';
		pld_10g_tx_fifo_num_reg	:	out	std_logic	:=	'0';
		pld_10g_tx_full_fifo	:	out	std_logic	:=	'0';
		pld_10g_tx_full_reg	:	out	std_logic	:=	'0';
		pld_10g_tx_pempty_reg	:	out	std_logic	:=	'0';
		pld_10g_tx_pfull_fifo	:	out	std_logic	:=	'0';
		pld_10g_tx_wordslip_exe_reg	:	out	std_logic	:=	'0';
		pld_10g_tx_wordslip_reg	:	out	std_logic	:=	'0';
		pld_pcs_tx_clk_out_10g_wire	:	out	std_logic	:=	'0';
		pld_tx_burst_en_reg	:	out	std_logic	:=	'0';
		pld_tx_control_lo_10g_reg	:	out	std_logic	:=	'0';
		pld_tx_data_10g_fifo	:	out	std_logic	:=	'0';
		pld_tx_data_lo_10g_reg	:	out	std_logic	:=	'0';
		distdwn_out_dv	:	out	std_logic	:=	'0';
		distdwn_out_rden	:	out	std_logic	:=	'0';
		distdwn_out_wren	:	out	std_logic	:=	'0';
		distup_out_dv	:	out	std_logic	:=	'0';
		distup_out_rden	:	out	std_logic	:=	'0';
		distup_out_wren	:	out	std_logic	:=	'0';
		tx_burst_en_exe	:	out	std_logic	:=	'0';
		tx_clk_out	:	out	std_logic	:=	'0';
		tx_clk_out_pld_if	:	out	std_logic	:=	'0';
		tx_clk_out_pma_if	:	out	std_logic	:=	'0';
		tx_control_out_krfec	:	out	std_logic_vector(8 downto 0)	:=	"000000000";
		tx_data_out_krfec	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		tx_data_valid_out_krfec	:	out	std_logic	:=	'0';
		tx_dft_clk_out	:	out	std_logic	:=	'0';
		tx_empty	:	out	std_logic	:=	'0';
		tx_fec_clk	:	out	std_logic	:=	'0';
		tx_fifo_num	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		tx_fifo_rd_ptr	:	out	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		tx_fifo_wr_clk	:	out	std_logic	:=	'0';
		tx_fifo_wr_data	:	out	std_logic_vector(72 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000000000000";
		tx_fifo_wr_data_dw	:	out	std_logic_vector(72 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000000000000";
		tx_fifo_wr_en	:	out	std_logic	:=	'0';
		tx_fifo_wr_ptr	:	out	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		tx_fifo_wr_rst_n	:	out	std_logic	:=	'0';
		tx_frame	:	out	std_logic	:=	'0';
		tx_full	:	out	std_logic	:=	'0';
		tx_master_clk	:	out	std_logic	:=	'0';
		tx_master_clk_rst_n	:	out	std_logic	:=	'0';
		tx_pempty	:	out	std_logic	:=	'0';
		tx_pfull	:	out	std_logic	:=	'0';
		tx_pma_data	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		tx_pma_gating_val	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		tx_test_data	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		tx_wordslip_exe	:	out	std_logic	:=	'0'
	);
end component;

begin



inst : twentynm_hssi_10g_tx_pcs_encrypted
	generic map (
		-- Instance parameters
		advanced_user_mode	=>	advanced_user_mode,
		bitslip_en	=>	bitslip_en,
		bonding_dft_en	=>	bonding_dft_en,
		bonding_dft_val	=>	bonding_dft_val,
		comp_cnt	=>	comp_cnt_int,
		compin_sel	=>	compin_sel,
		crcgen_bypass	=>	crcgen_bypass,
		crcgen_clken	=>	crcgen_clken,
		crcgen_err	=>	crcgen_err,
		crcgen_inv	=>	crcgen_inv,
		ctrl_bit_reverse	=>	ctrl_bit_reverse,
		ctrl_plane_bonding	=>	ctrl_plane_bonding,
		data_bit_reverse	=>	data_bit_reverse,
		dft_clk_out_sel	=>	dft_clk_out_sel,
		dispgen_bypass	=>	dispgen_bypass,
		dispgen_clken	=>	dispgen_clken,
		dispgen_err	=>	dispgen_err,
		dispgen_pipeln	=>	dispgen_pipeln,
		distdwn_bypass_pipeln	=>	distdwn_bypass_pipeln,
		distdwn_master	=>	distdwn_master,
		distup_bypass_pipeln	=>	distup_bypass_pipeln,
		distup_master	=>	distup_master,
		dv_bond	=>	dv_bond,
		empty_flag_type	=>	empty_flag_type,
		enc64b66b_txsm_clken	=>	enc64b66b_txsm_clken,
		enc_64b66b_txsm_bypass	=>	enc_64b66b_txsm_bypass,
		fastpath	=>	fastpath,
		fec_clken	=>	fec_clken,
		fec_enable	=>	fec_enable,
		fifo_double_write	=>	fifo_double_write,
		fifo_reg_fast	=>	fifo_reg_fast,
		fifo_stop_rd	=>	fifo_stop_rd,
		fifo_stop_wr	=>	fifo_stop_wr,
		frmgen_burst	=>	frmgen_burst,
		frmgen_bypass	=>	frmgen_bypass,
		frmgen_clken	=>	frmgen_clken,
		frmgen_mfrm_length	=>	frmgen_mfrm_length_int,
		frmgen_pipeln	=>	frmgen_pipeln,
		frmgen_pyld_ins	=>	frmgen_pyld_ins,
		frmgen_wordslip	=>	frmgen_wordslip,
		full_flag_type	=>	full_flag_type,
		gb_pipeln_bypass	=>	gb_pipeln_bypass,
		gb_tx_idwidth	=>	gb_tx_idwidth,
		gb_tx_odwidth	=>	gb_tx_odwidth,
		gbred_clken	=>	gbred_clken,
		indv	=>	indv,
		low_latency_en	=>	low_latency_en,
		master_clk_sel	=>	master_clk_sel,
		pempty_flag_type	=>	pempty_flag_type,
		pfull_flag_type	=>	pfull_flag_type,
		phcomp_rd_del	=>	phcomp_rd_del,
		pld_if_type	=>	pld_if_type,
		prot_mode	=>	prot_mode,
		pseudo_random	=>	pseudo_random,
		pseudo_seed_a	=>	pseudo_seed_a,
		pseudo_seed_b	=>	pseudo_seed_b,
		random_disp	=>	random_disp,
		rdfifo_clken	=>	rdfifo_clken,
		reconfig_settings	=>	reconfig_settings,
		scrm_bypass	=>	scrm_bypass,
		scrm_clken	=>	scrm_clken,
		scrm_mode	=>	scrm_mode,
		scrm_pipeln	=>	scrm_pipeln,
		sh_err	=>	sh_err,
		silicon_rev	=>	silicon_rev,
		sop_mark	=>	sop_mark,
		stretch_num_stages	=>	stretch_num_stages,
		sup_mode	=>	sup_mode,
		test_mode	=>	test_mode,
		tx_scrm_err	=>	tx_scrm_err,
		tx_scrm_width	=>	tx_scrm_width,
		tx_sh_location	=>	tx_sh_location,
		tx_sm_bypass	=>	tx_sm_bypass,
		tx_sm_pipeln	=>	tx_sm_pipeln,
		tx_testbus_sel	=>	tx_testbus_sel,
		txfifo_empty	=>	txfifo_empty,
		txfifo_full	=>	txfifo_full,
		txfifo_mode	=>	txfifo_mode,
		txfifo_pempty	=>	txfifo_pempty_int,
		txfifo_pfull	=>	txfifo_pfull_int,
		wr_clk_sel	=>	wr_clk_sel,
		wrfifo_clken	=>	wrfifo_clken
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		distdwn_in_dv	=>	distdwn_in_dv,
		distdwn_in_rden	=>	distdwn_in_rden,
		distdwn_in_wren	=>	distdwn_in_wren,
		distup_in_dv	=>	distup_in_dv,
		distup_in_rden	=>	distup_in_rden,
		distup_in_wren	=>	distup_in_wren,
		krfec_refclk_dig	=>	krfec_refclk_dig,
		r_tx_diag_word	=>	r_tx_diag_word,
		r_tx_scrm_word	=>	r_tx_scrm_word,
		r_tx_skip_word	=>	r_tx_skip_word,
		r_tx_sync_word	=>	r_tx_sync_word,
		refclk_dig	=>	refclk_dig,
		scan_mode_n	=>	scan_mode_n,
		tx_bitslip	=>	tx_bitslip,
		tx_burst_en	=>	tx_burst_en,
		tx_control	=>	tx_control,
		tx_control_reg	=>	tx_control_reg,
		tx_data	=>	tx_data,
		tx_data_in_krfec	=>	tx_data_in_krfec,
		tx_data_reg	=>	tx_data_reg,
		tx_data_valid	=>	tx_data_valid,
		tx_data_valid_reg	=>	tx_data_valid_reg,
		tx_diag_status	=>	tx_diag_status,
		tx_fifo_rd_data	=>	tx_fifo_rd_data,
		tx_pld_clk	=>	tx_pld_clk,
		tx_pld_rst_n	=>	tx_pld_rst_n,
		tx_pma_clk	=>	tx_pma_clk,
		tx_wordslip	=>	tx_wordslip,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		pld_10g_krfec_tx_frame_10g_reg	=>	pld_10g_krfec_tx_frame_10g_reg,
		pld_10g_krfec_tx_pld_rst_n_fifo	=>	pld_10g_krfec_tx_pld_rst_n_fifo,
		pld_10g_krfec_tx_pld_rst_n_reg	=>	pld_10g_krfec_tx_pld_rst_n_reg,
		pld_10g_tx_bitslip_reg	=>	pld_10g_tx_bitslip_reg,
		pld_10g_tx_burst_en_exe_reg	=>	pld_10g_tx_burst_en_exe_reg,
		pld_10g_tx_data_valid_10g_reg	=>	pld_10g_tx_data_valid_10g_reg,
		pld_10g_tx_data_valid_fifo	=>	pld_10g_tx_data_valid_fifo,
		pld_10g_tx_data_valid_reg	=>	pld_10g_tx_data_valid_reg,
		pld_10g_tx_diag_status_reg	=>	pld_10g_tx_diag_status_reg,
		pld_10g_tx_empty_reg	=>	pld_10g_tx_empty_reg,
		pld_10g_tx_fifo_num_reg	=>	pld_10g_tx_fifo_num_reg,
		pld_10g_tx_full_fifo	=>	pld_10g_tx_full_fifo,
		pld_10g_tx_full_reg	=>	pld_10g_tx_full_reg,
		pld_10g_tx_pempty_reg	=>	pld_10g_tx_pempty_reg,
		pld_10g_tx_pfull_fifo	=>	pld_10g_tx_pfull_fifo,
		pld_10g_tx_wordslip_exe_reg	=>	pld_10g_tx_wordslip_exe_reg,
		pld_10g_tx_wordslip_reg	=>	pld_10g_tx_wordslip_reg,
		pld_pcs_tx_clk_out_10g_wire	=>	pld_pcs_tx_clk_out_10g_wire,
		pld_tx_burst_en_reg	=>	pld_tx_burst_en_reg,
		pld_tx_control_lo_10g_reg	=>	pld_tx_control_lo_10g_reg,
		pld_tx_data_10g_fifo	=>	pld_tx_data_10g_fifo,
		pld_tx_data_lo_10g_reg	=>	pld_tx_data_lo_10g_reg,
		distdwn_out_dv	=>	distdwn_out_dv,
		distdwn_out_rden	=>	distdwn_out_rden,
		distdwn_out_wren	=>	distdwn_out_wren,
		distup_out_dv	=>	distup_out_dv,
		distup_out_rden	=>	distup_out_rden,
		distup_out_wren	=>	distup_out_wren,
		tx_burst_en_exe	=>	tx_burst_en_exe,
		tx_clk_out	=>	tx_clk_out,
		tx_clk_out_pld_if	=>	tx_clk_out_pld_if,
		tx_clk_out_pma_if	=>	tx_clk_out_pma_if,
		tx_control_out_krfec	=>	tx_control_out_krfec,
		tx_data_out_krfec	=>	tx_data_out_krfec,
		tx_data_valid_out_krfec	=>	tx_data_valid_out_krfec,
		tx_dft_clk_out	=>	tx_dft_clk_out,
		tx_empty	=>	tx_empty,
		tx_fec_clk	=>	tx_fec_clk,
		tx_fifo_num	=>	tx_fifo_num,
		tx_fifo_rd_ptr	=>	tx_fifo_rd_ptr,
		tx_fifo_wr_clk	=>	tx_fifo_wr_clk,
		tx_fifo_wr_data	=>	tx_fifo_wr_data,
		tx_fifo_wr_data_dw	=>	tx_fifo_wr_data_dw,
		tx_fifo_wr_en	=>	tx_fifo_wr_en,
		tx_fifo_wr_ptr	=>	tx_fifo_wr_ptr,
		tx_fifo_wr_rst_n	=>	tx_fifo_wr_rst_n,
		tx_frame	=>	tx_frame,
		tx_full	=>	tx_full,
		tx_master_clk	=>	tx_master_clk,
		tx_master_clk_rst_n	=>	tx_master_clk_rst_n,
		tx_pempty	=>	tx_pempty,
		tx_pfull	=>	tx_pfull,
		tx_pma_data	=>	tx_pma_data,
		tx_pma_gating_val	=>	tx_pma_gating_val,
		tx_test_data	=>	tx_test_data,
		tx_wordslip_exe	=>	tx_wordslip_exe
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_8g_rx_pcs	is
	generic (
		-- Entity parameters
		auto_error_replacement	:	string	:=	"dis_err_replace";
		auto_speed_nego	:	string	:=	"dis_asn";
		bit_reversal	:	string	:=	"dis_bit_reversal";
		bonding_dft_en	:	string	:=	"dft_dis";
		bonding_dft_val	:	string	:=	"dft_0";
		bypass_pipeline_reg	:	string	:=	"dis_bypass_pipeline";
		byte_deserializer	:	string	:=	"dis_bds";
		cdr_ctrl_rxvalid_mask	:	string	:=	"dis_rxvalid_mask";
		clkcmp_pattern_n	:	bit_vector	:=	B"00000000000000000000";
		clkcmp_pattern_p	:	bit_vector	:=	B"00000000000000000000";
		clock_gate_bds_dec_asn	:	string	:=	"dis_bds_dec_asn_clk_gating";
		clock_gate_cdr_eidle	:	string	:=	"dis_cdr_eidle_clk_gating";
		clock_gate_dw_pc_wrclk	:	string	:=	"dis_dw_pc_wrclk_gating";
		clock_gate_dw_rm_rd	:	string	:=	"dis_dw_rm_rdclk_gating";
		clock_gate_dw_rm_wr	:	string	:=	"dis_dw_rm_wrclk_gating";
		clock_gate_dw_wa	:	string	:=	"dis_dw_wa_clk_gating";
		clock_gate_pc_rdclk	:	string	:=	"dis_pc_rdclk_gating";
		clock_gate_sw_pc_wrclk	:	string	:=	"dis_sw_pc_wrclk_gating";
		clock_gate_sw_rm_rd	:	string	:=	"dis_sw_rm_rdclk_gating";
		clock_gate_sw_rm_wr	:	string	:=	"dis_sw_rm_wrclk_gating";
		clock_gate_sw_wa	:	string	:=	"dis_sw_wa_clk_gating";
		clock_observation_in_pld_core	:	string	:=	"internal_sw_wa_clk";
		ctrl_plane_bonding_compensation	:	string	:=	"dis_compensation";
		ctrl_plane_bonding_consumption	:	string	:=	"individual";
		ctrl_plane_bonding_distribution	:	string	:=	"not_master_chnl_distr";
		eidle_entry_eios	:	string	:=	"dis_eidle_eios";
		eidle_entry_iei	:	string	:=	"dis_eidle_iei";
		eidle_entry_sd	:	string	:=	"dis_eidle_sd";
		eightb_tenb_decoder	:	string	:=	"dis_8b10b";
		err_flags_sel	:	string	:=	"err_flags_wa";
		fixed_pat_det	:	string	:=	"dis_fixed_patdet";
		fixed_pat_num	:	bit_vector	:=	B"1111";
		force_signal_detect	:	string	:=	"en_force_signal_detect";
		gen3_clk_en	:	string	:=	"disable_clk";
		gen3_rx_clk_sel	:	string	:=	"rcvd_clk";
		gen3_tx_clk_sel	:	string	:=	"tx_pma_clk";
		hip_mode	:	string	:=	"dis_hip";
		ibm_invalid_code	:	string	:=	"dis_ibm_invalid_code";
		invalid_code_flag_only	:	string	:=	"dis_invalid_code_only";
		pad_or_edb_error_replace	:	string	:=	"replace_edb";
		pcs_bypass	:	string	:=	"dis_pcs_bypass";
		phase_comp_rdptr	:	string	:=	"enable_rdptr";
		phase_compensation_fifo	:	string	:=	"low_latency";
		pipe_if_enable	:	string	:=	"dis_pipe_rx";
		pma_dw	:	string	:=	"eight_bit";
		polinv_8b10b_dec	:	string	:=	"dis_polinv_8b10b_dec";
		prot_mode	:	string	:=	"gige";
		rate_match	:	string	:=	"dis_rm";
		rate_match_del_thres	:	string	:=	"dis_rm_del_thres";
		rate_match_empty_thres	:	string	:=	"dis_rm_empty_thres";
		rate_match_full_thres	:	string	:=	"dis_rm_full_thres";
		rate_match_ins_thres	:	string	:=	"dis_rm_ins_thres";
		rate_match_start_thres	:	string	:=	"dis_rm_start_thres";
		reconfig_settings	:	string	:=	"{}";
		rx_clk2	:	string	:=	"rcvd_clk_clk2";
		rx_clk_free_running	:	string	:=	"en_rx_clk_free_run";
		rx_pcs_urst	:	string	:=	"en_rx_pcs_urst";
		rx_rcvd_clk	:	string	:=	"rcvd_clk_rcvd_clk";
		rx_rd_clk	:	string	:=	"pld_rx_clk";
		rx_refclk	:	string	:=	"dis_refclk_sel";
		rx_wr_clk	:	string	:=	"rx_clk2_div_1_2_4";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode";
		symbol_swap	:	string	:=	"dis_symbol_swap";
		sync_sm_idle_eios	:	string	:=	"dis_syncsm_idle";
		test_bus_sel	:	string	:=	"tx_testbus";
		tx_rx_parallel_loopback	:	string	:=	"dis_plpbk";
		wa_boundary_lock_ctrl	:	string	:=	"bit_slip";
		wa_clk_slip_spacing	:	bit_vector	:=	B"0000010000";
		wa_det_latency_sync_status_beh	:	string	:=	"assert_sync_status_non_imm";
		wa_disp_err_flag	:	string	:=	"dis_disp_err_flag";
		wa_kchar	:	string	:=	"dis_kchar";
		wa_pd	:	string	:=	"wa_pd_10";
		wa_pd_data	:	string	:=	"0000000000000000000000000000000000000000";
		wa_pd_polarity	:	string	:=	"dis_pd_both_pol";
		wa_pld_controlled	:	string	:=	"dis_pld_ctrl";
		wa_renumber_data	:	bit_vector	:=	B"000000";
		wa_rgnumber_data	:	bit_vector	:=	B"00000000";
		wa_rknumber_data	:	bit_vector	:=	B"00000000";
		wa_rosnumber_data	:	bit_vector	:=	B"00";
		wa_rvnumber_data	:	bit_vector	:=	B"0000000000000";
		wa_sync_sm_ctrl	:	string	:=	"gige_sync_sm";
		wait_cnt	:	bit_vector	:=	B"000000000000"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		a1a2_size	:	in	std_logic	:=	'0';
		bit_reversal_enable	:	in	std_logic	:=	'0';
		bitslip	:	in	std_logic	:=	'0';
		byte_rev_en	:	in	std_logic	:=	'0';
		disable_pc_fifo_byte_serdes	:	in	std_logic	:=	'0';
		dyn_clk_switch_n	:	in	std_logic	:=	'0';
		eidleinfersel	:	in	std_logic_vector(2 downto 0)	:=	"000";
		eios_detected_cdr_ctrl	:	in	std_logic	:=	'0';
		enable_comma_detect	:	in	std_logic	:=	'0';
		gen3_clk_sel	:	in	std_logic	:=	'0';
		hrd_rst	:	in	std_logic	:=	'0';
		inferred_rxvalid_cdr_ctrl	:	in	std_logic	:=	'0';
		pcie_switch	:	in	std_logic	:=	'0';
		pcs_rst	:	in	std_logic	:=	'0';
		phystatus_int	:	in	std_logic	:=	'0';
		phystatus_pcs_gen3	:	in	std_logic	:=	'0';
		pipe_loopbk	:	in	std_logic	:=	'0';
		pld_rx_clk	:	in	std_logic	:=	'0';
		polarity_inversion	:	in	std_logic	:=	'0';
		datain	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		rcvd_clk_pma	:	in	std_logic	:=	'0';
		rd_data1_rx_rmfifo	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rd_data2_rx_rmfifo	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rd_data_rx_phfifo	:	in	std_logic_vector(79 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
		rd_enable_in_chnl_down	:	in	std_logic	:=	'0';
		rd_enable_in_chnl_up	:	in	std_logic	:=	'0';
		rm_fifo_read_enable	:	in	std_logic	:=	'0';
		pc_fifo_rd_enable	:	in	std_logic	:=	'0';
		refclk_dig	:	in	std_logic	:=	'0';
		refclk_dig2	:	in	std_logic	:=	'0';
		reset_pc_ptrs_asn	:	in	std_logic	:=	'0';
		reset_pc_ptrs_in_chnl_down	:	in	std_logic	:=	'0';
		reset_pc_ptrs_in_chnl_up	:	in	std_logic	:=	'0';
		reset_ppm_cntrs_pcs_pma	:	in	std_logic	:=	'0';
		rx_blk_start_pcs_gen3	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rx_data_pcs_gen3	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		rx_data_valid_pcs_gen3	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rx_div_sync_in_chnl_down	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rx_div_sync_in_chnl_up	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rx_sync_hdr_pcs_gen3	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rx_we_in_chnl_down	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rx_we_in_chnl_up	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxstatus_int	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus_pcs_gen3	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rx_pcs_rst	:	in	std_logic	:=	'0';
		rxvalid_int	:	in	std_logic	:=	'0';
		rxvalid_pcs_gen3	:	in	std_logic	:=	'0';
		scan_mode_n	:	in	std_logic	:=	'0';
		sig_det_from_pma	:	in	std_logic	:=	'0';
		soft_reset_wclk1_n	:	in	std_logic	:=	'0';
		speed_change	:	in	std_logic	:=	'0';
		sw_fifo_wr_clk	:	in	std_logic	:=	'0';
		syncsm_en	:	in	std_logic	:=	'0';
		tx_clk_out	:	in	std_logic	:=	'0';
		tx_ctrlplane_testbus	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		tx_div_sync	:	in	std_logic_vector(1 downto 0)	:=	"00";
		tx_pma_clk	:	in	std_logic	:=	'0';
		tx_testbus	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		wr_enable_in_chnl_down	:	in	std_logic	:=	'0';
		wr_enable_in_chnl_up	:	in	std_logic	:=	'0';
		pc_fifo_wrdisable	:	in	std_logic	:=	'0';
		rm_fifo_write_enable	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		byte_deserializer_pcs_clk_div_by_2_reg	:	out	std_logic	:=	'0';
		byte_deserializer_pcs_clk_div_by_2_txclk_reg	:	out	std_logic	:=	'0';
		byte_deserializer_pcs_clk_div_by_2_txclk_wire	:	out	std_logic	:=	'0';
		byte_deserializer_pcs_clk_div_by_2_wire	:	out	std_logic	:=	'0';
		byte_deserializer_pcs_clk_div_by_4_txclk_reg	:	out	std_logic	:=	'0';
		byte_deserializer_pld_clk_div_by_2_reg	:	out	std_logic	:=	'0';
		byte_deserializer_pld_clk_div_by_2_txclk_reg	:	out	std_logic	:=	'0';
		byte_deserializer_pld_clk_div_by_4_txclk_reg	:	out	std_logic	:=	'0';
		pld_8g_a1a2_k1k2_flag_reg	:	out	std_logic	:=	'0';
		pld_8g_a1a2_k1k2_flag_txclk_reg	:	out	std_logic	:=	'0';
		pld_8g_a1a2_size_reg	:	out	std_logic	:=	'0';
		pld_8g_a1a2_size_txclk_reg	:	out	std_logic	:=	'0';
		pld_8g_bitloc_rev_en_reg	:	out	std_logic	:=	'0';
		pld_8g_bitloc_rev_en_txclk_reg	:	out	std_logic	:=	'0';
		pld_8g_byte_rev_en_reg	:	out	std_logic	:=	'0';
		pld_8g_byte_rev_en_txclk_reg	:	out	std_logic	:=	'0';
		pld_8g_elecidle_reg	:	out	std_logic	:=	'0';
		pld_8g_empty_rmf_lowlatency_reg	:	out	std_logic	:=	'0';
		pld_8g_empty_rmf_lowlatency_txclk_reg	:	out	std_logic	:=	'0';
		pld_8g_empty_rmf_reg	:	out	std_logic	:=	'0';
		pld_8g_empty_rmf_txclk_reg	:	out	std_logic	:=	'0';
		pld_8g_empty_rx_fifo	:	out	std_logic	:=	'0';
		pld_8g_empty_rx_reg	:	out	std_logic	:=	'0';
		pld_8g_empty_rx_txclk_reg	:	out	std_logic	:=	'0';
		pld_8g_encdt_reg	:	out	std_logic	:=	'0';
		pld_8g_encdt_txclk_reg	:	out	std_logic	:=	'0';
		pld_8g_full_rmf_reg	:	out	std_logic	:=	'0';
		pld_8g_full_rmf_txclk_reg	:	out	std_logic	:=	'0';
		pld_8g_full_rx_fifo	:	out	std_logic	:=	'0';
		pld_8g_full_rx_reg	:	out	std_logic	:=	'0';
		pld_8g_full_rx_txclk_reg	:	out	std_logic	:=	'0';
		pld_8g_g3_rx_pld_rst_n_reg	:	out	std_logic	:=	'0';
		pld_8g_g3_rx_pld_rst_n_txclk_reg	:	out	std_logic	:=	'0';
		pld_8g_rxelecidle_txclk_reg	:	out	std_logic	:=	'0';
		pld_8g_rxpolarity_reg	:	out	std_logic	:=	'0';
		pld_8g_rxpolarity_txclk_reg	:	out	std_logic	:=	'0';
		pld_8g_wa_boundary_reg	:	out	std_logic	:=	'0';
		pld_8g_wrdisable_rx_reg	:	out	std_logic	:=	'0';
		pld_8g_wrdisable_rx_txclk_reg	:	out	std_logic	:=	'0';
		pld_pcs_rx_clk_out_8g_div_by_2_txclk_wire	:	out	std_logic	:=	'0';
		pld_pcs_rx_clk_out_8g_div_by_2_wire	:	out	std_logic	:=	'0';
		pld_pcs_rx_clk_out_8g_txclk_wire	:	out	std_logic	:=	'0';
		pld_pcs_rx_clk_out_8g_wire	:	out	std_logic	:=	'0';
		pld_rx_control_8g_reg	:	out	std_logic	:=	'0';
		pld_rx_control_8g_txclk_reg	:	out	std_logic	:=	'0';
		pld_rx_data_8g_reg	:	out	std_logic	:=	'0';
		pld_rx_data_8g_txclk_reg	:	out	std_logic	:=	'0';
		pld_syncsm_en_reg	:	out	std_logic	:=	'0';
		pld_syncsm_en_txclk_reg	:	out	std_logic	:=	'0';
		sta_rx_clk2_by2_1	:	out	std_logic	:=	'0';
		sta_rx_clk2_by2_1_out	:	out	std_logic	:=	'0';
		sta_rx_clk2_by2_2	:	out	std_logic	:=	'0';
		sta_rx_clk2_by2_2_out	:	out	std_logic	:=	'0';
		sta_rx_clk2_by4_1	:	out	std_logic	:=	'0';
		sta_rx_clk2_by4_1_out	:	out	std_logic	:=	'0';
		a1a2k1k2flag	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		rm_fifo_partial_full	:	out	std_logic	:=	'0';
		rm_fifo_partial_empty	:	out	std_logic	:=	'0';
		chnl_test_bus_out	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		dis_pc_byte	:	out	std_logic	:=	'0';
		eios_det_cdr_ctrl	:	out	std_logic_vector(2 downto 0)	:=	"000";
		rm_fifo_empty	:	out	std_logic	:=	'0';
		pc_fifo_empty	:	out	std_logic	:=	'0';
		rm_fifo_full	:	out	std_logic	:=	'0';
		pcfifofull	:	out	std_logic	:=	'0';
		g3_rx_pma_rstn	:	out	std_logic	:=	'0';
		g3_rx_rcvd_rstn	:	out	std_logic	:=	'0';
		gen2ngen1	:	out	std_logic	:=	'0';
		phystatus	:	out	std_logic	:=	'0';
		pipe_data	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		rd_enable_out_chnl_down	:	out	std_logic	:=	'0';
		rd_enable_out_chnl_up	:	out	std_logic	:=	'0';
		rd_ptr1_rx_rmfifo	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		rd_ptr2_rx_rmfifo	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		rd_ptr_rx_phfifo	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		reset_pc_ptrs	:	out	std_logic	:=	'0';
		reset_pc_ptrs_in_chnl_down_pipe	:	out	std_logic	:=	'0';
		reset_pc_ptrs_in_chnl_up_pipe	:	out	std_logic	:=	'0';
		reset_pc_ptrs_out_chnl_down	:	out	std_logic	:=	'0';
		reset_pc_ptrs_out_chnl_up	:	out	std_logic	:=	'0';
		parallel_rev_loopback	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		rx_blk_start	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		clock_to_pld	:	out	std_logic	:=	'0';
		rx_clk_out_pld_if	:	out	std_logic	:=	'0';
		rx_clk_to_observation_ff_in_pld_if	:	out	std_logic	:=	'0';
		rx_clkslip	:	out	std_logic	:=	'0';
		rx_data_valid	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		rx_div_sync_out_chnl_down	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rx_div_sync_out_chnl_up	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rx_pipe_clk	:	out	std_logic	:=	'0';
		rx_pipe_soft_reset	:	out	std_logic	:=	'0';
		rx_pma_clk_gen3	:	out	std_logic	:=	'0';
		rx_rcvd_clk_gen3	:	out	std_logic	:=	'0';
		rx_rstn_sync2wrfifo_8g	:	out	std_logic	:=	'0';
		rx_sync_hdr	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rx_we_out_chnl_down	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rx_we_out_chnl_up	:	out	std_logic_vector(1 downto 0)	:=	"00";
		dataout	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		eidle_detected	:	out	std_logic	:=	'0';
		rxstatus	:	out	std_logic_vector(2 downto 0)	:=	"000";
		rxvalid	:	out	std_logic	:=	'0';
		signal_detect_out	:	out	std_logic	:=	'0';
		word_align_boundary	:	out	std_logic_vector(4 downto 0)	:=	"00000";
		wr_clk_rx_phfifo_dw_clk	:	out	std_logic	:=	'0';
		wr_clk_rx_phfifo_sw_clk	:	out	std_logic	:=	'0';
		wr_clk_rx_rmfifo_dw_clk	:	out	std_logic	:=	'0';
		wr_clk_rx_rmfifo_sw_clk	:	out	std_logic	:=	'0';
		wr_data_rx_phfifo	:	out	std_logic_vector(79 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
		wr_data_rx_rmfifo	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		wr_en_rx_phfifo	:	out	std_logic	:=	'0';
		wr_en_rx_rmfifo	:	out	std_logic	:=	'0';
		wr_enable_out_chnl_down	:	out	std_logic	:=	'0';
		wr_enable_out_chnl_up	:	out	std_logic	:=	'0';
		wr_ptr_rx_phfifo	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		wr_ptr_rx_rmfifo	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		wr_rst_n_rx_phfifo	:	out	std_logic	:=	'0';
		wr_rst_rx_rmfifo	:	out	std_logic	:=	'0'
	);
end twentynm_hssi_8g_rx_pcs;

architecture behavior of twentynm_hssi_8g_rx_pcs	is

constant clkcmp_pattern_n_int	:	integer	:=	bin2int(clkcmp_pattern_n);
constant clkcmp_pattern_p_int	:	integer	:=	bin2int(clkcmp_pattern_p);
constant fixed_pat_num_int	:	integer	:=	bin2int(fixed_pat_num);
constant wa_clk_slip_spacing_int	:	integer	:=	bin2int(wa_clk_slip_spacing);
constant wa_renumber_data_int	:	integer	:=	bin2int(wa_renumber_data);
constant wa_rgnumber_data_int	:	integer	:=	bin2int(wa_rgnumber_data);
constant wa_rknumber_data_int	:	integer	:=	bin2int(wa_rknumber_data);
constant wa_rosnumber_data_int	:	integer	:=	bin2int(wa_rosnumber_data);
constant wa_rvnumber_data_int	:	integer	:=	bin2int(wa_rvnumber_data);
constant wait_cnt_int	:	integer	:=	bin2int(wait_cnt);



component	twentynm_hssi_8g_rx_pcs_encrypted
	generic (
		-- Architecture parameters
		auto_error_replacement	:	string	:=	"dis_err_replace";
		auto_speed_nego	:	string	:=	"dis_asn";
		bit_reversal	:	string	:=	"dis_bit_reversal";
		bonding_dft_en	:	string	:=	"dft_dis";
		bonding_dft_val	:	string	:=	"dft_0";
		bypass_pipeline_reg	:	string	:=	"dis_bypass_pipeline";
		byte_deserializer	:	string	:=	"dis_bds";
		cdr_ctrl_rxvalid_mask	:	string	:=	"dis_rxvalid_mask";
		clkcmp_pattern_n	:	integer	:=	0;
		clkcmp_pattern_p	:	integer	:=	0;
		clock_gate_bds_dec_asn	:	string	:=	"dis_bds_dec_asn_clk_gating";
		clock_gate_cdr_eidle	:	string	:=	"dis_cdr_eidle_clk_gating";
		clock_gate_dw_pc_wrclk	:	string	:=	"dis_dw_pc_wrclk_gating";
		clock_gate_dw_rm_rd	:	string	:=	"dis_dw_rm_rdclk_gating";
		clock_gate_dw_rm_wr	:	string	:=	"dis_dw_rm_wrclk_gating";
		clock_gate_dw_wa	:	string	:=	"dis_dw_wa_clk_gating";
		clock_gate_pc_rdclk	:	string	:=	"dis_pc_rdclk_gating";
		clock_gate_sw_pc_wrclk	:	string	:=	"dis_sw_pc_wrclk_gating";
		clock_gate_sw_rm_rd	:	string	:=	"dis_sw_rm_rdclk_gating";
		clock_gate_sw_rm_wr	:	string	:=	"dis_sw_rm_wrclk_gating";
		clock_gate_sw_wa	:	string	:=	"dis_sw_wa_clk_gating";
		clock_observation_in_pld_core	:	string	:=	"internal_sw_wa_clk";
		ctrl_plane_bonding_compensation	:	string	:=	"dis_compensation";
		ctrl_plane_bonding_consumption	:	string	:=	"individual";
		ctrl_plane_bonding_distribution	:	string	:=	"not_master_chnl_distr";
		eidle_entry_eios	:	string	:=	"dis_eidle_eios";
		eidle_entry_iei	:	string	:=	"dis_eidle_iei";
		eidle_entry_sd	:	string	:=	"dis_eidle_sd";
		eightb_tenb_decoder	:	string	:=	"dis_8b10b";
		err_flags_sel	:	string	:=	"err_flags_wa";
		fixed_pat_det	:	string	:=	"dis_fixed_patdet";
		fixed_pat_num	:	integer	:=	15;
		force_signal_detect	:	string	:=	"en_force_signal_detect";
		gen3_clk_en	:	string	:=	"disable_clk";
		gen3_rx_clk_sel	:	string	:=	"rcvd_clk";
		gen3_tx_clk_sel	:	string	:=	"tx_pma_clk";
		hip_mode	:	string	:=	"dis_hip";
		ibm_invalid_code	:	string	:=	"dis_ibm_invalid_code";
		invalid_code_flag_only	:	string	:=	"dis_invalid_code_only";
		pad_or_edb_error_replace	:	string	:=	"replace_edb";
		pcs_bypass	:	string	:=	"dis_pcs_bypass";
		phase_comp_rdptr	:	string	:=	"enable_rdptr";
		phase_compensation_fifo	:	string	:=	"low_latency";
		pipe_if_enable	:	string	:=	"dis_pipe_rx";
		pma_dw	:	string	:=	"eight_bit";
		polinv_8b10b_dec	:	string	:=	"dis_polinv_8b10b_dec";
		prot_mode	:	string	:=	"gige";
		rate_match	:	string	:=	"dis_rm";
		rate_match_del_thres	:	string	:=	"dis_rm_del_thres";
		rate_match_empty_thres	:	string	:=	"dis_rm_empty_thres";
		rate_match_full_thres	:	string	:=	"dis_rm_full_thres";
		rate_match_ins_thres	:	string	:=	"dis_rm_ins_thres";
		rate_match_start_thres	:	string	:=	"dis_rm_start_thres";
		reconfig_settings	:	string	:=	"{}";
		rx_clk2	:	string	:=	"rcvd_clk_clk2";
		rx_clk_free_running	:	string	:=	"en_rx_clk_free_run";
		rx_pcs_urst	:	string	:=	"en_rx_pcs_urst";
		rx_rcvd_clk	:	string	:=	"rcvd_clk_rcvd_clk";
		rx_rd_clk	:	string	:=	"pld_rx_clk";
		rx_refclk	:	string	:=	"dis_refclk_sel";
		rx_wr_clk	:	string	:=	"rx_clk2_div_1_2_4";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode";
		symbol_swap	:	string	:=	"dis_symbol_swap";
		sync_sm_idle_eios	:	string	:=	"dis_syncsm_idle";
		test_bus_sel	:	string	:=	"tx_testbus";
		tx_rx_parallel_loopback	:	string	:=	"dis_plpbk";
		wa_boundary_lock_ctrl	:	string	:=	"bit_slip";
		wa_clk_slip_spacing	:	integer	:=	16;
		wa_det_latency_sync_status_beh	:	string	:=	"assert_sync_status_non_imm";
		wa_disp_err_flag	:	string	:=	"dis_disp_err_flag";
		wa_kchar	:	string	:=	"dis_kchar";
		wa_pd	:	string	:=	"wa_pd_10";
		wa_pd_data	:	string	:=	"0000000000000000000000000000000000000000";
		wa_pd_polarity	:	string	:=	"dis_pd_both_pol";
		wa_pld_controlled	:	string	:=	"dis_pld_ctrl";
		wa_renumber_data	:	integer	:=	0;
		wa_rgnumber_data	:	integer	:=	0;
		wa_rknumber_data	:	integer	:=	0;
		wa_rosnumber_data	:	integer	:=	0;
		wa_rvnumber_data	:	integer	:=	0;
		wa_sync_sm_ctrl	:	string	:=	"gige_sync_sm";
		wait_cnt	:	integer	:=	0
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		a1a2_size	:	in	std_logic	:=	'0';
		bit_reversal_enable	:	in	std_logic	:=	'0';
		bitslip	:	in	std_logic	:=	'0';
		byte_rev_en	:	in	std_logic	:=	'0';
		disable_pc_fifo_byte_serdes	:	in	std_logic	:=	'0';
		dyn_clk_switch_n	:	in	std_logic	:=	'0';
		eidleinfersel	:	in	std_logic_vector(2 downto 0)	:=	"000";
		eios_detected_cdr_ctrl	:	in	std_logic	:=	'0';
		enable_comma_detect	:	in	std_logic	:=	'0';
		gen3_clk_sel	:	in	std_logic	:=	'0';
		hrd_rst	:	in	std_logic	:=	'0';
		inferred_rxvalid_cdr_ctrl	:	in	std_logic	:=	'0';
		pcie_switch	:	in	std_logic	:=	'0';
		pcs_rst	:	in	std_logic	:=	'0';
		phystatus_int	:	in	std_logic	:=	'0';
		phystatus_pcs_gen3	:	in	std_logic	:=	'0';
		pipe_loopbk	:	in	std_logic	:=	'0';
		pld_rx_clk	:	in	std_logic	:=	'0';
		polarity_inversion	:	in	std_logic	:=	'0';
		datain	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		rcvd_clk_pma	:	in	std_logic	:=	'0';
		rd_data1_rx_rmfifo	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rd_data2_rx_rmfifo	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rd_data_rx_phfifo	:	in	std_logic_vector(79 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
		rd_enable_in_chnl_down	:	in	std_logic	:=	'0';
		rd_enable_in_chnl_up	:	in	std_logic	:=	'0';
		rm_fifo_read_enable	:	in	std_logic	:=	'0';
		pc_fifo_rd_enable	:	in	std_logic	:=	'0';
		refclk_dig	:	in	std_logic	:=	'0';
		refclk_dig2	:	in	std_logic	:=	'0';
		reset_pc_ptrs_asn	:	in	std_logic	:=	'0';
		reset_pc_ptrs_in_chnl_down	:	in	std_logic	:=	'0';
		reset_pc_ptrs_in_chnl_up	:	in	std_logic	:=	'0';
		reset_ppm_cntrs_pcs_pma	:	in	std_logic	:=	'0';
		rx_blk_start_pcs_gen3	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rx_data_pcs_gen3	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		rx_data_valid_pcs_gen3	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rx_div_sync_in_chnl_down	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rx_div_sync_in_chnl_up	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rx_sync_hdr_pcs_gen3	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rx_we_in_chnl_down	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rx_we_in_chnl_up	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxstatus_int	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus_pcs_gen3	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rx_pcs_rst	:	in	std_logic	:=	'0';
		rxvalid_int	:	in	std_logic	:=	'0';
		rxvalid_pcs_gen3	:	in	std_logic	:=	'0';
		scan_mode_n	:	in	std_logic	:=	'0';
		sig_det_from_pma	:	in	std_logic	:=	'0';
		soft_reset_wclk1_n	:	in	std_logic	:=	'0';
		speed_change	:	in	std_logic	:=	'0';
		sw_fifo_wr_clk	:	in	std_logic	:=	'0';
		syncsm_en	:	in	std_logic	:=	'0';
		tx_clk_out	:	in	std_logic	:=	'0';
		tx_ctrlplane_testbus	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		tx_div_sync	:	in	std_logic_vector(1 downto 0)	:=	"00";
		tx_pma_clk	:	in	std_logic	:=	'0';
		tx_testbus	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		wr_enable_in_chnl_down	:	in	std_logic	:=	'0';
		wr_enable_in_chnl_up	:	in	std_logic	:=	'0';
		pc_fifo_wrdisable	:	in	std_logic	:=	'0';
		rm_fifo_write_enable	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		byte_deserializer_pcs_clk_div_by_2_reg	:	out	std_logic	:=	'0';
		byte_deserializer_pcs_clk_div_by_2_txclk_reg	:	out	std_logic	:=	'0';
		byte_deserializer_pcs_clk_div_by_2_txclk_wire	:	out	std_logic	:=	'0';
		byte_deserializer_pcs_clk_div_by_2_wire	:	out	std_logic	:=	'0';
		byte_deserializer_pcs_clk_div_by_4_txclk_reg	:	out	std_logic	:=	'0';
		byte_deserializer_pld_clk_div_by_2_reg	:	out	std_logic	:=	'0';
		byte_deserializer_pld_clk_div_by_2_txclk_reg	:	out	std_logic	:=	'0';
		byte_deserializer_pld_clk_div_by_4_txclk_reg	:	out	std_logic	:=	'0';
		pld_8g_a1a2_k1k2_flag_reg	:	out	std_logic	:=	'0';
		pld_8g_a1a2_k1k2_flag_txclk_reg	:	out	std_logic	:=	'0';
		pld_8g_a1a2_size_reg	:	out	std_logic	:=	'0';
		pld_8g_a1a2_size_txclk_reg	:	out	std_logic	:=	'0';
		pld_8g_bitloc_rev_en_reg	:	out	std_logic	:=	'0';
		pld_8g_bitloc_rev_en_txclk_reg	:	out	std_logic	:=	'0';
		pld_8g_byte_rev_en_reg	:	out	std_logic	:=	'0';
		pld_8g_byte_rev_en_txclk_reg	:	out	std_logic	:=	'0';
		pld_8g_elecidle_reg	:	out	std_logic	:=	'0';
		pld_8g_empty_rmf_lowlatency_reg	:	out	std_logic	:=	'0';
		pld_8g_empty_rmf_lowlatency_txclk_reg	:	out	std_logic	:=	'0';
		pld_8g_empty_rmf_reg	:	out	std_logic	:=	'0';
		pld_8g_empty_rmf_txclk_reg	:	out	std_logic	:=	'0';
		pld_8g_empty_rx_fifo	:	out	std_logic	:=	'0';
		pld_8g_empty_rx_reg	:	out	std_logic	:=	'0';
		pld_8g_empty_rx_txclk_reg	:	out	std_logic	:=	'0';
		pld_8g_encdt_reg	:	out	std_logic	:=	'0';
		pld_8g_encdt_txclk_reg	:	out	std_logic	:=	'0';
		pld_8g_full_rmf_reg	:	out	std_logic	:=	'0';
		pld_8g_full_rmf_txclk_reg	:	out	std_logic	:=	'0';
		pld_8g_full_rx_fifo	:	out	std_logic	:=	'0';
		pld_8g_full_rx_reg	:	out	std_logic	:=	'0';
		pld_8g_full_rx_txclk_reg	:	out	std_logic	:=	'0';
		pld_8g_g3_rx_pld_rst_n_reg	:	out	std_logic	:=	'0';
		pld_8g_g3_rx_pld_rst_n_txclk_reg	:	out	std_logic	:=	'0';
		pld_8g_rxelecidle_txclk_reg	:	out	std_logic	:=	'0';
		pld_8g_rxpolarity_reg	:	out	std_logic	:=	'0';
		pld_8g_rxpolarity_txclk_reg	:	out	std_logic	:=	'0';
		pld_8g_wa_boundary_reg	:	out	std_logic	:=	'0';
		pld_8g_wrdisable_rx_reg	:	out	std_logic	:=	'0';
		pld_8g_wrdisable_rx_txclk_reg	:	out	std_logic	:=	'0';
		pld_pcs_rx_clk_out_8g_div_by_2_txclk_wire	:	out	std_logic	:=	'0';
		pld_pcs_rx_clk_out_8g_div_by_2_wire	:	out	std_logic	:=	'0';
		pld_pcs_rx_clk_out_8g_txclk_wire	:	out	std_logic	:=	'0';
		pld_pcs_rx_clk_out_8g_wire	:	out	std_logic	:=	'0';
		pld_rx_control_8g_reg	:	out	std_logic	:=	'0';
		pld_rx_control_8g_txclk_reg	:	out	std_logic	:=	'0';
		pld_rx_data_8g_reg	:	out	std_logic	:=	'0';
		pld_rx_data_8g_txclk_reg	:	out	std_logic	:=	'0';
		pld_syncsm_en_reg	:	out	std_logic	:=	'0';
		pld_syncsm_en_txclk_reg	:	out	std_logic	:=	'0';
		sta_rx_clk2_by2_1	:	out	std_logic	:=	'0';
		sta_rx_clk2_by2_1_out	:	out	std_logic	:=	'0';
		sta_rx_clk2_by2_2	:	out	std_logic	:=	'0';
		sta_rx_clk2_by2_2_out	:	out	std_logic	:=	'0';
		sta_rx_clk2_by4_1	:	out	std_logic	:=	'0';
		sta_rx_clk2_by4_1_out	:	out	std_logic	:=	'0';
		a1a2k1k2flag	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		rm_fifo_partial_full	:	out	std_logic	:=	'0';
		rm_fifo_partial_empty	:	out	std_logic	:=	'0';
		chnl_test_bus_out	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		dis_pc_byte	:	out	std_logic	:=	'0';
		eios_det_cdr_ctrl	:	out	std_logic_vector(2 downto 0)	:=	"000";
		rm_fifo_empty	:	out	std_logic	:=	'0';
		pc_fifo_empty	:	out	std_logic	:=	'0';
		rm_fifo_full	:	out	std_logic	:=	'0';
		pcfifofull	:	out	std_logic	:=	'0';
		g3_rx_pma_rstn	:	out	std_logic	:=	'0';
		g3_rx_rcvd_rstn	:	out	std_logic	:=	'0';
		gen2ngen1	:	out	std_logic	:=	'0';
		phystatus	:	out	std_logic	:=	'0';
		pipe_data	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		rd_enable_out_chnl_down	:	out	std_logic	:=	'0';
		rd_enable_out_chnl_up	:	out	std_logic	:=	'0';
		rd_ptr1_rx_rmfifo	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		rd_ptr2_rx_rmfifo	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		rd_ptr_rx_phfifo	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		reset_pc_ptrs	:	out	std_logic	:=	'0';
		reset_pc_ptrs_in_chnl_down_pipe	:	out	std_logic	:=	'0';
		reset_pc_ptrs_in_chnl_up_pipe	:	out	std_logic	:=	'0';
		reset_pc_ptrs_out_chnl_down	:	out	std_logic	:=	'0';
		reset_pc_ptrs_out_chnl_up	:	out	std_logic	:=	'0';
		parallel_rev_loopback	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		rx_blk_start	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		clock_to_pld	:	out	std_logic	:=	'0';
		rx_clk_out_pld_if	:	out	std_logic	:=	'0';
		rx_clk_to_observation_ff_in_pld_if	:	out	std_logic	:=	'0';
		rx_clkslip	:	out	std_logic	:=	'0';
		rx_data_valid	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		rx_div_sync_out_chnl_down	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rx_div_sync_out_chnl_up	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rx_pipe_clk	:	out	std_logic	:=	'0';
		rx_pipe_soft_reset	:	out	std_logic	:=	'0';
		rx_pma_clk_gen3	:	out	std_logic	:=	'0';
		rx_rcvd_clk_gen3	:	out	std_logic	:=	'0';
		rx_rstn_sync2wrfifo_8g	:	out	std_logic	:=	'0';
		rx_sync_hdr	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rx_we_out_chnl_down	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rx_we_out_chnl_up	:	out	std_logic_vector(1 downto 0)	:=	"00";
		dataout	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		eidle_detected	:	out	std_logic	:=	'0';
		rxstatus	:	out	std_logic_vector(2 downto 0)	:=	"000";
		rxvalid	:	out	std_logic	:=	'0';
		signal_detect_out	:	out	std_logic	:=	'0';
		word_align_boundary	:	out	std_logic_vector(4 downto 0)	:=	"00000";
		wr_clk_rx_phfifo_dw_clk	:	out	std_logic	:=	'0';
		wr_clk_rx_phfifo_sw_clk	:	out	std_logic	:=	'0';
		wr_clk_rx_rmfifo_dw_clk	:	out	std_logic	:=	'0';
		wr_clk_rx_rmfifo_sw_clk	:	out	std_logic	:=	'0';
		wr_data_rx_phfifo	:	out	std_logic_vector(79 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
		wr_data_rx_rmfifo	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		wr_en_rx_phfifo	:	out	std_logic	:=	'0';
		wr_en_rx_rmfifo	:	out	std_logic	:=	'0';
		wr_enable_out_chnl_down	:	out	std_logic	:=	'0';
		wr_enable_out_chnl_up	:	out	std_logic	:=	'0';
		wr_ptr_rx_phfifo	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		wr_ptr_rx_rmfifo	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		wr_rst_n_rx_phfifo	:	out	std_logic	:=	'0';
		wr_rst_rx_rmfifo	:	out	std_logic	:=	'0'
	);
end component;

begin



inst : twentynm_hssi_8g_rx_pcs_encrypted
	generic map (
		-- Instance parameters
		auto_error_replacement	=>	auto_error_replacement,
		auto_speed_nego	=>	auto_speed_nego,
		bit_reversal	=>	bit_reversal,
		bonding_dft_en	=>	bonding_dft_en,
		bonding_dft_val	=>	bonding_dft_val,
		bypass_pipeline_reg	=>	bypass_pipeline_reg,
		byte_deserializer	=>	byte_deserializer,
		cdr_ctrl_rxvalid_mask	=>	cdr_ctrl_rxvalid_mask,
		clkcmp_pattern_n	=>	clkcmp_pattern_n_int,
		clkcmp_pattern_p	=>	clkcmp_pattern_p_int,
		clock_gate_bds_dec_asn	=>	clock_gate_bds_dec_asn,
		clock_gate_cdr_eidle	=>	clock_gate_cdr_eidle,
		clock_gate_dw_pc_wrclk	=>	clock_gate_dw_pc_wrclk,
		clock_gate_dw_rm_rd	=>	clock_gate_dw_rm_rd,
		clock_gate_dw_rm_wr	=>	clock_gate_dw_rm_wr,
		clock_gate_dw_wa	=>	clock_gate_dw_wa,
		clock_gate_pc_rdclk	=>	clock_gate_pc_rdclk,
		clock_gate_sw_pc_wrclk	=>	clock_gate_sw_pc_wrclk,
		clock_gate_sw_rm_rd	=>	clock_gate_sw_rm_rd,
		clock_gate_sw_rm_wr	=>	clock_gate_sw_rm_wr,
		clock_gate_sw_wa	=>	clock_gate_sw_wa,
		clock_observation_in_pld_core	=>	clock_observation_in_pld_core,
		ctrl_plane_bonding_compensation	=>	ctrl_plane_bonding_compensation,
		ctrl_plane_bonding_consumption	=>	ctrl_plane_bonding_consumption,
		ctrl_plane_bonding_distribution	=>	ctrl_plane_bonding_distribution,
		eidle_entry_eios	=>	eidle_entry_eios,
		eidle_entry_iei	=>	eidle_entry_iei,
		eidle_entry_sd	=>	eidle_entry_sd,
		eightb_tenb_decoder	=>	eightb_tenb_decoder,
		err_flags_sel	=>	err_flags_sel,
		fixed_pat_det	=>	fixed_pat_det,
		fixed_pat_num	=>	fixed_pat_num_int,
		force_signal_detect	=>	force_signal_detect,
		gen3_clk_en	=>	gen3_clk_en,
		gen3_rx_clk_sel	=>	gen3_rx_clk_sel,
		gen3_tx_clk_sel	=>	gen3_tx_clk_sel,
		hip_mode	=>	hip_mode,
		ibm_invalid_code	=>	ibm_invalid_code,
		invalid_code_flag_only	=>	invalid_code_flag_only,
		pad_or_edb_error_replace	=>	pad_or_edb_error_replace,
		pcs_bypass	=>	pcs_bypass,
		phase_comp_rdptr	=>	phase_comp_rdptr,
		phase_compensation_fifo	=>	phase_compensation_fifo,
		pipe_if_enable	=>	pipe_if_enable,
		pma_dw	=>	pma_dw,
		polinv_8b10b_dec	=>	polinv_8b10b_dec,
		prot_mode	=>	prot_mode,
		rate_match	=>	rate_match,
		rate_match_del_thres	=>	rate_match_del_thres,
		rate_match_empty_thres	=>	rate_match_empty_thres,
		rate_match_full_thres	=>	rate_match_full_thres,
		rate_match_ins_thres	=>	rate_match_ins_thres,
		rate_match_start_thres	=>	rate_match_start_thres,
		reconfig_settings	=>	reconfig_settings,
		rx_clk2	=>	rx_clk2,
		rx_clk_free_running	=>	rx_clk_free_running,
		rx_pcs_urst	=>	rx_pcs_urst,
		rx_rcvd_clk	=>	rx_rcvd_clk,
		rx_rd_clk	=>	rx_rd_clk,
		rx_refclk	=>	rx_refclk,
		rx_wr_clk	=>	rx_wr_clk,
		silicon_rev	=>	silicon_rev,
		sup_mode	=>	sup_mode,
		symbol_swap	=>	symbol_swap,
		sync_sm_idle_eios	=>	sync_sm_idle_eios,
		test_bus_sel	=>	test_bus_sel,
		tx_rx_parallel_loopback	=>	tx_rx_parallel_loopback,
		wa_boundary_lock_ctrl	=>	wa_boundary_lock_ctrl,
		wa_clk_slip_spacing	=>	wa_clk_slip_spacing_int,
		wa_det_latency_sync_status_beh	=>	wa_det_latency_sync_status_beh,
		wa_disp_err_flag	=>	wa_disp_err_flag,
		wa_kchar	=>	wa_kchar,
		wa_pd	=>	wa_pd,
		wa_pd_data	=>	wa_pd_data,
		wa_pd_polarity	=>	wa_pd_polarity,
		wa_pld_controlled	=>	wa_pld_controlled,
		wa_renumber_data	=>	wa_renumber_data_int,
		wa_rgnumber_data	=>	wa_rgnumber_data_int,
		wa_rknumber_data	=>	wa_rknumber_data_int,
		wa_rosnumber_data	=>	wa_rosnumber_data_int,
		wa_rvnumber_data	=>	wa_rvnumber_data_int,
		wa_sync_sm_ctrl	=>	wa_sync_sm_ctrl,
		wait_cnt	=>	wait_cnt_int
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		a1a2_size	=>	a1a2_size,
		bit_reversal_enable	=>	bit_reversal_enable,
		bitslip	=>	bitslip,
		byte_rev_en	=>	byte_rev_en,
		disable_pc_fifo_byte_serdes	=>	disable_pc_fifo_byte_serdes,
		dyn_clk_switch_n	=>	dyn_clk_switch_n,
		eidleinfersel	=>	eidleinfersel,
		eios_detected_cdr_ctrl	=>	eios_detected_cdr_ctrl,
		enable_comma_detect	=>	enable_comma_detect,
		gen3_clk_sel	=>	gen3_clk_sel,
		hrd_rst	=>	hrd_rst,
		inferred_rxvalid_cdr_ctrl	=>	inferred_rxvalid_cdr_ctrl,
		pcie_switch	=>	pcie_switch,
		pcs_rst	=>	pcs_rst,
		phystatus_int	=>	phystatus_int,
		phystatus_pcs_gen3	=>	phystatus_pcs_gen3,
		pipe_loopbk	=>	pipe_loopbk,
		pld_rx_clk	=>	pld_rx_clk,
		polarity_inversion	=>	polarity_inversion,
		datain	=>	datain,
		rcvd_clk_pma	=>	rcvd_clk_pma,
		rd_data1_rx_rmfifo	=>	rd_data1_rx_rmfifo,
		rd_data2_rx_rmfifo	=>	rd_data2_rx_rmfifo,
		rd_data_rx_phfifo	=>	rd_data_rx_phfifo,
		rd_enable_in_chnl_down	=>	rd_enable_in_chnl_down,
		rd_enable_in_chnl_up	=>	rd_enable_in_chnl_up,
		rm_fifo_read_enable	=>	rm_fifo_read_enable,
		pc_fifo_rd_enable	=>	pc_fifo_rd_enable,
		refclk_dig	=>	refclk_dig,
		refclk_dig2	=>	refclk_dig2,
		reset_pc_ptrs_asn	=>	reset_pc_ptrs_asn,
		reset_pc_ptrs_in_chnl_down	=>	reset_pc_ptrs_in_chnl_down,
		reset_pc_ptrs_in_chnl_up	=>	reset_pc_ptrs_in_chnl_up,
		reset_ppm_cntrs_pcs_pma	=>	reset_ppm_cntrs_pcs_pma,
		rx_blk_start_pcs_gen3	=>	rx_blk_start_pcs_gen3,
		rx_data_pcs_gen3	=>	rx_data_pcs_gen3,
		rx_data_valid_pcs_gen3	=>	rx_data_valid_pcs_gen3,
		rx_div_sync_in_chnl_down	=>	rx_div_sync_in_chnl_down,
		rx_div_sync_in_chnl_up	=>	rx_div_sync_in_chnl_up,
		rx_sync_hdr_pcs_gen3	=>	rx_sync_hdr_pcs_gen3,
		rx_we_in_chnl_down	=>	rx_we_in_chnl_down,
		rx_we_in_chnl_up	=>	rx_we_in_chnl_up,
		rxstatus_int	=>	rxstatus_int,
		rxstatus_pcs_gen3	=>	rxstatus_pcs_gen3,
		rx_pcs_rst	=>	rx_pcs_rst,
		rxvalid_int	=>	rxvalid_int,
		rxvalid_pcs_gen3	=>	rxvalid_pcs_gen3,
		scan_mode_n	=>	scan_mode_n,
		sig_det_from_pma	=>	sig_det_from_pma,
		soft_reset_wclk1_n	=>	soft_reset_wclk1_n,
		speed_change	=>	speed_change,
		sw_fifo_wr_clk	=>	sw_fifo_wr_clk,
		syncsm_en	=>	syncsm_en,
		tx_clk_out	=>	tx_clk_out,
		tx_ctrlplane_testbus	=>	tx_ctrlplane_testbus,
		tx_div_sync	=>	tx_div_sync,
		tx_pma_clk	=>	tx_pma_clk,
		tx_testbus	=>	tx_testbus,
		wr_enable_in_chnl_down	=>	wr_enable_in_chnl_down,
		wr_enable_in_chnl_up	=>	wr_enable_in_chnl_up,
		pc_fifo_wrdisable	=>	pc_fifo_wrdisable,
		rm_fifo_write_enable	=>	rm_fifo_write_enable,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		byte_deserializer_pcs_clk_div_by_2_reg	=>	byte_deserializer_pcs_clk_div_by_2_reg,
		byte_deserializer_pcs_clk_div_by_2_txclk_reg	=>	byte_deserializer_pcs_clk_div_by_2_txclk_reg,
		byte_deserializer_pcs_clk_div_by_2_txclk_wire	=>	byte_deserializer_pcs_clk_div_by_2_txclk_wire,
		byte_deserializer_pcs_clk_div_by_2_wire	=>	byte_deserializer_pcs_clk_div_by_2_wire,
		byte_deserializer_pcs_clk_div_by_4_txclk_reg	=>	byte_deserializer_pcs_clk_div_by_4_txclk_reg,
		byte_deserializer_pld_clk_div_by_2_reg	=>	byte_deserializer_pld_clk_div_by_2_reg,
		byte_deserializer_pld_clk_div_by_2_txclk_reg	=>	byte_deserializer_pld_clk_div_by_2_txclk_reg,
		byte_deserializer_pld_clk_div_by_4_txclk_reg	=>	byte_deserializer_pld_clk_div_by_4_txclk_reg,
		pld_8g_a1a2_k1k2_flag_reg	=>	pld_8g_a1a2_k1k2_flag_reg,
		pld_8g_a1a2_k1k2_flag_txclk_reg	=>	pld_8g_a1a2_k1k2_flag_txclk_reg,
		pld_8g_a1a2_size_reg	=>	pld_8g_a1a2_size_reg,
		pld_8g_a1a2_size_txclk_reg	=>	pld_8g_a1a2_size_txclk_reg,
		pld_8g_bitloc_rev_en_reg	=>	pld_8g_bitloc_rev_en_reg,
		pld_8g_bitloc_rev_en_txclk_reg	=>	pld_8g_bitloc_rev_en_txclk_reg,
		pld_8g_byte_rev_en_reg	=>	pld_8g_byte_rev_en_reg,
		pld_8g_byte_rev_en_txclk_reg	=>	pld_8g_byte_rev_en_txclk_reg,
		pld_8g_elecidle_reg	=>	pld_8g_elecidle_reg,
		pld_8g_empty_rmf_lowlatency_reg	=>	pld_8g_empty_rmf_lowlatency_reg,
		pld_8g_empty_rmf_lowlatency_txclk_reg	=>	pld_8g_empty_rmf_lowlatency_txclk_reg,
		pld_8g_empty_rmf_reg	=>	pld_8g_empty_rmf_reg,
		pld_8g_empty_rmf_txclk_reg	=>	pld_8g_empty_rmf_txclk_reg,
		pld_8g_empty_rx_fifo	=>	pld_8g_empty_rx_fifo,
		pld_8g_empty_rx_reg	=>	pld_8g_empty_rx_reg,
		pld_8g_empty_rx_txclk_reg	=>	pld_8g_empty_rx_txclk_reg,
		pld_8g_encdt_reg	=>	pld_8g_encdt_reg,
		pld_8g_encdt_txclk_reg	=>	pld_8g_encdt_txclk_reg,
		pld_8g_full_rmf_reg	=>	pld_8g_full_rmf_reg,
		pld_8g_full_rmf_txclk_reg	=>	pld_8g_full_rmf_txclk_reg,
		pld_8g_full_rx_fifo	=>	pld_8g_full_rx_fifo,
		pld_8g_full_rx_reg	=>	pld_8g_full_rx_reg,
		pld_8g_full_rx_txclk_reg	=>	pld_8g_full_rx_txclk_reg,
		pld_8g_g3_rx_pld_rst_n_reg	=>	pld_8g_g3_rx_pld_rst_n_reg,
		pld_8g_g3_rx_pld_rst_n_txclk_reg	=>	pld_8g_g3_rx_pld_rst_n_txclk_reg,
		pld_8g_rxelecidle_txclk_reg	=>	pld_8g_rxelecidle_txclk_reg,
		pld_8g_rxpolarity_reg	=>	pld_8g_rxpolarity_reg,
		pld_8g_rxpolarity_txclk_reg	=>	pld_8g_rxpolarity_txclk_reg,
		pld_8g_wa_boundary_reg	=>	pld_8g_wa_boundary_reg,
		pld_8g_wrdisable_rx_reg	=>	pld_8g_wrdisable_rx_reg,
		pld_8g_wrdisable_rx_txclk_reg	=>	pld_8g_wrdisable_rx_txclk_reg,
		pld_pcs_rx_clk_out_8g_div_by_2_txclk_wire	=>	pld_pcs_rx_clk_out_8g_div_by_2_txclk_wire,
		pld_pcs_rx_clk_out_8g_div_by_2_wire	=>	pld_pcs_rx_clk_out_8g_div_by_2_wire,
		pld_pcs_rx_clk_out_8g_txclk_wire	=>	pld_pcs_rx_clk_out_8g_txclk_wire,
		pld_pcs_rx_clk_out_8g_wire	=>	pld_pcs_rx_clk_out_8g_wire,
		pld_rx_control_8g_reg	=>	pld_rx_control_8g_reg,
		pld_rx_control_8g_txclk_reg	=>	pld_rx_control_8g_txclk_reg,
		pld_rx_data_8g_reg	=>	pld_rx_data_8g_reg,
		pld_rx_data_8g_txclk_reg	=>	pld_rx_data_8g_txclk_reg,
		pld_syncsm_en_reg	=>	pld_syncsm_en_reg,
		pld_syncsm_en_txclk_reg	=>	pld_syncsm_en_txclk_reg,
		sta_rx_clk2_by2_1	=>	sta_rx_clk2_by2_1,
		sta_rx_clk2_by2_1_out	=>	sta_rx_clk2_by2_1_out,
		sta_rx_clk2_by2_2	=>	sta_rx_clk2_by2_2,
		sta_rx_clk2_by2_2_out	=>	sta_rx_clk2_by2_2_out,
		sta_rx_clk2_by4_1	=>	sta_rx_clk2_by4_1,
		sta_rx_clk2_by4_1_out	=>	sta_rx_clk2_by4_1_out,
		a1a2k1k2flag	=>	a1a2k1k2flag,
		rm_fifo_partial_full	=>	rm_fifo_partial_full,
		rm_fifo_partial_empty	=>	rm_fifo_partial_empty,
		chnl_test_bus_out	=>	chnl_test_bus_out,
		dis_pc_byte	=>	dis_pc_byte,
		eios_det_cdr_ctrl	=>	eios_det_cdr_ctrl,
		rm_fifo_empty	=>	rm_fifo_empty,
		pc_fifo_empty	=>	pc_fifo_empty,
		rm_fifo_full	=>	rm_fifo_full,
		pcfifofull	=>	pcfifofull,
		g3_rx_pma_rstn	=>	g3_rx_pma_rstn,
		g3_rx_rcvd_rstn	=>	g3_rx_rcvd_rstn,
		gen2ngen1	=>	gen2ngen1,
		phystatus	=>	phystatus,
		pipe_data	=>	pipe_data,
		rd_enable_out_chnl_down	=>	rd_enable_out_chnl_down,
		rd_enable_out_chnl_up	=>	rd_enable_out_chnl_up,
		rd_ptr1_rx_rmfifo	=>	rd_ptr1_rx_rmfifo,
		rd_ptr2_rx_rmfifo	=>	rd_ptr2_rx_rmfifo,
		rd_ptr_rx_phfifo	=>	rd_ptr_rx_phfifo,
		reset_pc_ptrs	=>	reset_pc_ptrs,
		reset_pc_ptrs_in_chnl_down_pipe	=>	reset_pc_ptrs_in_chnl_down_pipe,
		reset_pc_ptrs_in_chnl_up_pipe	=>	reset_pc_ptrs_in_chnl_up_pipe,
		reset_pc_ptrs_out_chnl_down	=>	reset_pc_ptrs_out_chnl_down,
		reset_pc_ptrs_out_chnl_up	=>	reset_pc_ptrs_out_chnl_up,
		parallel_rev_loopback	=>	parallel_rev_loopback,
		rx_blk_start	=>	rx_blk_start,
		clock_to_pld	=>	clock_to_pld,
		rx_clk_out_pld_if	=>	rx_clk_out_pld_if,
		rx_clk_to_observation_ff_in_pld_if	=>	rx_clk_to_observation_ff_in_pld_if,
		rx_clkslip	=>	rx_clkslip,
		rx_data_valid	=>	rx_data_valid,
		rx_div_sync_out_chnl_down	=>	rx_div_sync_out_chnl_down,
		rx_div_sync_out_chnl_up	=>	rx_div_sync_out_chnl_up,
		rx_pipe_clk	=>	rx_pipe_clk,
		rx_pipe_soft_reset	=>	rx_pipe_soft_reset,
		rx_pma_clk_gen3	=>	rx_pma_clk_gen3,
		rx_rcvd_clk_gen3	=>	rx_rcvd_clk_gen3,
		rx_rstn_sync2wrfifo_8g	=>	rx_rstn_sync2wrfifo_8g,
		rx_sync_hdr	=>	rx_sync_hdr,
		rx_we_out_chnl_down	=>	rx_we_out_chnl_down,
		rx_we_out_chnl_up	=>	rx_we_out_chnl_up,
		dataout	=>	dataout,
		eidle_detected	=>	eidle_detected,
		rxstatus	=>	rxstatus,
		rxvalid	=>	rxvalid,
		signal_detect_out	=>	signal_detect_out,
		word_align_boundary	=>	word_align_boundary,
		wr_clk_rx_phfifo_dw_clk	=>	wr_clk_rx_phfifo_dw_clk,
		wr_clk_rx_phfifo_sw_clk	=>	wr_clk_rx_phfifo_sw_clk,
		wr_clk_rx_rmfifo_dw_clk	=>	wr_clk_rx_rmfifo_dw_clk,
		wr_clk_rx_rmfifo_sw_clk	=>	wr_clk_rx_rmfifo_sw_clk,
		wr_data_rx_phfifo	=>	wr_data_rx_phfifo,
		wr_data_rx_rmfifo	=>	wr_data_rx_rmfifo,
		wr_en_rx_phfifo	=>	wr_en_rx_phfifo,
		wr_en_rx_rmfifo	=>	wr_en_rx_rmfifo,
		wr_enable_out_chnl_down	=>	wr_enable_out_chnl_down,
		wr_enable_out_chnl_up	=>	wr_enable_out_chnl_up,
		wr_ptr_rx_phfifo	=>	wr_ptr_rx_phfifo,
		wr_ptr_rx_rmfifo	=>	wr_ptr_rx_rmfifo,
		wr_rst_n_rx_phfifo	=>	wr_rst_n_rx_phfifo,
		wr_rst_rx_rmfifo	=>	wr_rst_rx_rmfifo
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_8g_tx_pcs	is
	generic (
		-- Entity parameters
		auto_speed_nego_gen2	:	string	:=	"dis_asn_g2";
		bit_reversal	:	string	:=	"dis_bit_reversal";
		bonding_dft_en	:	string	:=	"dft_dis";
		bonding_dft_val	:	string	:=	"dft_0";
		bypass_pipeline_reg	:	string	:=	"dis_bypass_pipeline";
		byte_serializer	:	string	:=	"dis_bs";
		clock_gate_bs_enc	:	string	:=	"dis_bs_enc_clk_gating";
		clock_gate_dw_fifowr	:	string	:=	"dis_dw_fifowr_clk_gating";
		clock_gate_fiford	:	string	:=	"dis_fiford_clk_gating";
		clock_gate_sw_fifowr	:	string	:=	"dis_sw_fifowr_clk_gating";
		clock_observation_in_pld_core	:	string	:=	"internal_refclk_b";
		ctrl_plane_bonding_compensation	:	string	:=	"dis_compensation";
		ctrl_plane_bonding_consumption	:	string	:=	"individual";
		ctrl_plane_bonding_distribution	:	string	:=	"not_master_chnl_distr";
		data_selection_8b10b_encoder_input	:	string	:=	"normal_data_path";
		dynamic_clk_switch	:	string	:=	"dis_dyn_clk_switch";
		eightb_tenb_disp_ctrl	:	string	:=	"dis_disp_ctrl";
		eightb_tenb_encoder	:	string	:=	"dis_8b10b";
		force_echar	:	string	:=	"dis_force_echar";
		force_kchar	:	string	:=	"dis_force_kchar";
		gen3_tx_clk_sel	:	string	:=	"tx_pma_clk";
		gen3_tx_pipe_clk_sel	:	string	:=	"func_clk";
		hip_mode	:	string	:=	"dis_hip";
		pcs_bypass	:	string	:=	"dis_pcs_bypass";
		phase_comp_rdptr	:	string	:=	"enable_rdptr";
		phase_compensation_fifo	:	string	:=	"low_latency";
		phfifo_write_clk_sel	:	string	:=	"pld_tx_clk";
		pma_dw	:	string	:=	"eight_bit";
		prot_mode	:	string	:=	"basic";
		reconfig_settings	:	string	:=	"{}";
		refclk_b_clk_sel	:	string	:=	"tx_pma_clock";
		revloop_back_rm	:	string	:=	"dis_rev_loopback_rx_rm";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode";
		symbol_swap	:	string	:=	"dis_symbol_swap";
		tx_bitslip	:	string	:=	"dis_tx_bitslip";
		tx_compliance_controlled_disparity	:	string	:=	"dis_txcompliance";
		tx_fast_pld_reg	:	string	:=	"dis_tx_fast_pld_reg";
		txclk_freerun	:	string	:=	"dis_freerun_tx";
		txpcs_urst	:	string	:=	"en_txpcs_urst"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		clk_sel_gen3	:	in	std_logic	:=	'0';
		dis_pc_byte	:	in	std_logic	:=	'0';
		eidleinfersel	:	in	std_logic_vector(2 downto 0)	:=	"000";
		fifo_select_in_chnl_down	:	in	std_logic_vector(1 downto 0)	:=	"00";
		fifo_select_in_chnl_up	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rate_switch	:	in	std_logic	:=	'0';
		hrdrst	:	in	std_logic	:=	'0';
		pcs_rst	:	in	std_logic	:=	'0';
		pipe_tx_deemph	:	in	std_logic	:=	'0';
		pipe_tx_margin	:	in	std_logic_vector(2 downto 0)	:=	"000";
		coreclk	:	in	std_logic	:=	'0';
		powerdn	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rd_data_tx_phfifo	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		rd_enable_in_chnl_down	:	in	std_logic	:=	'0';
		rd_enable_in_chnl_up	:	in	std_logic	:=	'0';
		ph_fifo_rd_disable	:	in	std_logic	:=	'0';
		refclk_dig	:	in	std_logic	:=	'0';
		reset_pc_ptrs	:	in	std_logic	:=	'0';
		reset_pc_ptrs_in_chnl_down	:	in	std_logic	:=	'0';
		reset_pc_ptrs_in_chnl_up	:	in	std_logic	:=	'0';
		rev_parallel_lpbk_data	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		en_rev_parallel_lpbk	:	in	std_logic	:=	'0';
		pipe_en_rev_parallel_lpbk_in	:	in	std_logic	:=	'0';
		rxpolarity	:	in	std_logic	:=	'0';
		scan_mode_n	:	in	std_logic	:=	'0';
		tx_blk_start	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		bitslip_boundary_select	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		tx_data_valid	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		tx_div_sync_in_chnl_down	:	in	std_logic_vector(1 downto 0)	:=	"00";
		tx_div_sync_in_chnl_up	:	in	std_logic_vector(1 downto 0)	:=	"00";
		tx_sync_hdr	:	in	std_logic_vector(1 downto 0)	:=	"00";
		datain	:	in	std_logic_vector(43 downto 0)	:=	"00000000000000000000000000000000000000000000";
		txd_fast_reg	:	in	std_logic_vector(43 downto 0)	:=	"00000000000000000000000000000000000000000000";
		detectrxloopin	:	in	std_logic	:=	'0';
		txpma_local_clk	:	in	std_logic	:=	'0';
		txswing	:	in	std_logic	:=	'0';
		tx_pcs_reset	:	in	std_logic	:=	'0';
		wr_enable_in_chnl_down	:	in	std_logic	:=	'0';
		wr_enable_in_chnl_up	:	in	std_logic	:=	'0';
		wrenable_tx	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		byte_serializer_pcs_clk_div_by_2_reg	:	out	std_logic	:=	'0';
		byte_serializer_pcs_clk_div_by_2_wire	:	out	std_logic	:=	'0';
		byte_serializer_pcs_clk_div_by_4_reg	:	out	std_logic	:=	'0';
		byte_serializer_pld_clk_div_by_2_reg	:	out	std_logic	:=	'0';
		byte_serializer_pld_clk_div_by_4_reg	:	out	std_logic	:=	'0';
		pld_8g_empty_tx_fifo	:	out	std_logic	:=	'0';
		pld_8g_empty_tx_reg	:	out	std_logic	:=	'0';
		pld_8g_full_tx_fifo	:	out	std_logic	:=	'0';
		pld_8g_full_tx_reg	:	out	std_logic	:=	'0';
		pld_8g_g3_tx_pld_rst_n_reg	:	out	std_logic	:=	'0';
		pld_8g_rddisable_tx_reg	:	out	std_logic	:=	'0';
		pld_8g_tx_boundary_sel_reg	:	out	std_logic	:=	'0';
		pld_pcs_tx_clk_out_8g_div_by_2_wire	:	out	std_logic	:=	'0';
		pld_pcs_tx_clk_out_8g_wire	:	out	std_logic	:=	'0';
		pld_tx_data_8g_fifo	:	out	std_logic	:=	'0';
		pld_tx_data_lo_8g_reg	:	out	std_logic	:=	'0';
		sta_tx_clk2_by2_1	:	out	std_logic	:=	'0';
		sta_tx_clk2_by2_1_out	:	out	std_logic	:=	'0';
		sta_tx_clk2_by4_1	:	out	std_logic	:=	'0';
		sta_tx_clk2_by4_1_out	:	out	std_logic	:=	'0';
		dyn_clk_switch_n	:	out	std_logic	:=	'0';
		ph_fifo_underflow	:	out	std_logic	:=	'0';
		fifo_select_out_chnl_down	:	out	std_logic_vector(1 downto 0)	:=	"00";
		fifo_select_out_chnl_up	:	out	std_logic_vector(1 downto 0)	:=	"00";
		ph_fifo_overflow	:	out	std_logic	:=	'0';
		g3_pipe_tx_pma_rstn	:	out	std_logic	:=	'0';
		g3_tx_pma_rstn	:	out	std_logic	:=	'0';
		non_gray_eidleinfersel	:	out	std_logic_vector(2 downto 0)	:=	"000";
		phfifo_txdeemph	:	out	std_logic	:=	'0';
		phfifo_txmargin	:	out	std_logic_vector(2 downto 0)	:=	"000";
		phfifo_txswing	:	out	std_logic	:=	'0';
		pipe_tx_clk_out_gen3	:	out	std_logic	:=	'0';
		pmaif_asn_rstn	:	out	std_logic	:=	'0';
		pipe_power_down_out	:	out	std_logic_vector(1 downto 0)	:=	"00";
		dataout	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		rd_enable_out_chnl_down	:	out	std_logic	:=	'0';
		rd_enable_out_chnl_up	:	out	std_logic	:=	'0';
		rd_ptr_tx_phfifo	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		refclk_b	:	out	std_logic	:=	'0';
		refclk_b_reset	:	out	std_logic	:=	'0';
		pipe_en_rev_parallel_lpbk_out	:	out	std_logic	:=	'0';
		rxpolarity_int	:	out	std_logic	:=	'0';
		soft_reset_wclk1_n	:	out	std_logic	:=	'0';
		sw_fifo_wr_clk	:	out	std_logic	:=	'0';
		tx_blk_start_out	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		clk_out	:	out	std_logic	:=	'0';
		tx_clk_out_8g_pmaif	:	out	std_logic	:=	'0';
		clk_out_gen3	:	out	std_logic	:=	'0';
		tx_clk_out_pld_if	:	out	std_logic	:=	'0';
		tx_clk_out_pmaif	:	out	std_logic	:=	'0';
		tx_clk_to_observation_ff_in_pld_if	:	out	std_logic	:=	'0';
		tx_ctrlplane_testbus	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		tx_data_out	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		tx_data_valid_out	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		tx_datak_out	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		tx_div_sync	:	out	std_logic_vector(1 downto 0)	:=	"00";
		tx_div_sync_out_chnl_down	:	out	std_logic_vector(1 downto 0)	:=	"00";
		tx_div_sync_out_chnl_up	:	out	std_logic_vector(1 downto 0)	:=	"00";
		tx_pipe_clk	:	out	std_logic	:=	'0';
		tx_pipe_electidle	:	out	std_logic	:=	'0';
		tx_pipe_soft_reset	:	out	std_logic	:=	'0';
		tx_sync_hdr_out	:	out	std_logic_vector(1 downto 0)	:=	"00";
		tx_testbus	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		txcompliance_out	:	out	std_logic	:=	'0';
		tx_detect_rxloopback_int	:	out	std_logic	:=	'0';
		txelecidle_out	:	out	std_logic	:=	'0';
		wr_clk_tx_phfifo_dw_clk	:	out	std_logic	:=	'0';
		wr_clk_tx_phfifo_sw_clk	:	out	std_logic	:=	'0';
		wr_data_tx_phfifo	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		wr_en_tx_phfifo	:	out	std_logic	:=	'0';
		wr_enable_out_chnl_down	:	out	std_logic	:=	'0';
		wr_enable_out_chnl_up	:	out	std_logic	:=	'0';
		wr_ptr_tx_phfifo	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		wr_rst_n_tx_phfifo	:	out	std_logic	:=	'0'
	);
end twentynm_hssi_8g_tx_pcs;

architecture behavior of twentynm_hssi_8g_tx_pcs	is




component	twentynm_hssi_8g_tx_pcs_encrypted
	generic (
		-- Architecture parameters
		auto_speed_nego_gen2	:	string	:=	"dis_asn_g2";
		bit_reversal	:	string	:=	"dis_bit_reversal";
		bonding_dft_en	:	string	:=	"dft_dis";
		bonding_dft_val	:	string	:=	"dft_0";
		bypass_pipeline_reg	:	string	:=	"dis_bypass_pipeline";
		byte_serializer	:	string	:=	"dis_bs";
		clock_gate_bs_enc	:	string	:=	"dis_bs_enc_clk_gating";
		clock_gate_dw_fifowr	:	string	:=	"dis_dw_fifowr_clk_gating";
		clock_gate_fiford	:	string	:=	"dis_fiford_clk_gating";
		clock_gate_sw_fifowr	:	string	:=	"dis_sw_fifowr_clk_gating";
		clock_observation_in_pld_core	:	string	:=	"internal_refclk_b";
		ctrl_plane_bonding_compensation	:	string	:=	"dis_compensation";
		ctrl_plane_bonding_consumption	:	string	:=	"individual";
		ctrl_plane_bonding_distribution	:	string	:=	"not_master_chnl_distr";
		data_selection_8b10b_encoder_input	:	string	:=	"normal_data_path";
		dynamic_clk_switch	:	string	:=	"dis_dyn_clk_switch";
		eightb_tenb_disp_ctrl	:	string	:=	"dis_disp_ctrl";
		eightb_tenb_encoder	:	string	:=	"dis_8b10b";
		force_echar	:	string	:=	"dis_force_echar";
		force_kchar	:	string	:=	"dis_force_kchar";
		gen3_tx_clk_sel	:	string	:=	"tx_pma_clk";
		gen3_tx_pipe_clk_sel	:	string	:=	"func_clk";
		hip_mode	:	string	:=	"dis_hip";
		pcs_bypass	:	string	:=	"dis_pcs_bypass";
		phase_comp_rdptr	:	string	:=	"enable_rdptr";
		phase_compensation_fifo	:	string	:=	"low_latency";
		phfifo_write_clk_sel	:	string	:=	"pld_tx_clk";
		pma_dw	:	string	:=	"eight_bit";
		prot_mode	:	string	:=	"basic";
		reconfig_settings	:	string	:=	"{}";
		refclk_b_clk_sel	:	string	:=	"tx_pma_clock";
		revloop_back_rm	:	string	:=	"dis_rev_loopback_rx_rm";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode";
		symbol_swap	:	string	:=	"dis_symbol_swap";
		tx_bitslip	:	string	:=	"dis_tx_bitslip";
		tx_compliance_controlled_disparity	:	string	:=	"dis_txcompliance";
		tx_fast_pld_reg	:	string	:=	"dis_tx_fast_pld_reg";
		txclk_freerun	:	string	:=	"dis_freerun_tx";
		txpcs_urst	:	string	:=	"en_txpcs_urst"
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		clk_sel_gen3	:	in	std_logic	:=	'0';
		dis_pc_byte	:	in	std_logic	:=	'0';
		eidleinfersel	:	in	std_logic_vector(2 downto 0)	:=	"000";
		fifo_select_in_chnl_down	:	in	std_logic_vector(1 downto 0)	:=	"00";
		fifo_select_in_chnl_up	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rate_switch	:	in	std_logic	:=	'0';
		hrdrst	:	in	std_logic	:=	'0';
		pcs_rst	:	in	std_logic	:=	'0';
		pipe_tx_deemph	:	in	std_logic	:=	'0';
		pipe_tx_margin	:	in	std_logic_vector(2 downto 0)	:=	"000";
		coreclk	:	in	std_logic	:=	'0';
		powerdn	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rd_data_tx_phfifo	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		rd_enable_in_chnl_down	:	in	std_logic	:=	'0';
		rd_enable_in_chnl_up	:	in	std_logic	:=	'0';
		ph_fifo_rd_disable	:	in	std_logic	:=	'0';
		refclk_dig	:	in	std_logic	:=	'0';
		reset_pc_ptrs	:	in	std_logic	:=	'0';
		reset_pc_ptrs_in_chnl_down	:	in	std_logic	:=	'0';
		reset_pc_ptrs_in_chnl_up	:	in	std_logic	:=	'0';
		rev_parallel_lpbk_data	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		en_rev_parallel_lpbk	:	in	std_logic	:=	'0';
		pipe_en_rev_parallel_lpbk_in	:	in	std_logic	:=	'0';
		rxpolarity	:	in	std_logic	:=	'0';
		scan_mode_n	:	in	std_logic	:=	'0';
		tx_blk_start	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		bitslip_boundary_select	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		tx_data_valid	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		tx_div_sync_in_chnl_down	:	in	std_logic_vector(1 downto 0)	:=	"00";
		tx_div_sync_in_chnl_up	:	in	std_logic_vector(1 downto 0)	:=	"00";
		tx_sync_hdr	:	in	std_logic_vector(1 downto 0)	:=	"00";
		datain	:	in	std_logic_vector(43 downto 0)	:=	"00000000000000000000000000000000000000000000";
		txd_fast_reg	:	in	std_logic_vector(43 downto 0)	:=	"00000000000000000000000000000000000000000000";
		detectrxloopin	:	in	std_logic	:=	'0';
		txpma_local_clk	:	in	std_logic	:=	'0';
		txswing	:	in	std_logic	:=	'0';
		tx_pcs_reset	:	in	std_logic	:=	'0';
		wr_enable_in_chnl_down	:	in	std_logic	:=	'0';
		wr_enable_in_chnl_up	:	in	std_logic	:=	'0';
		wrenable_tx	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		byte_serializer_pcs_clk_div_by_2_reg	:	out	std_logic	:=	'0';
		byte_serializer_pcs_clk_div_by_2_wire	:	out	std_logic	:=	'0';
		byte_serializer_pcs_clk_div_by_4_reg	:	out	std_logic	:=	'0';
		byte_serializer_pld_clk_div_by_2_reg	:	out	std_logic	:=	'0';
		byte_serializer_pld_clk_div_by_4_reg	:	out	std_logic	:=	'0';
		pld_8g_empty_tx_fifo	:	out	std_logic	:=	'0';
		pld_8g_empty_tx_reg	:	out	std_logic	:=	'0';
		pld_8g_full_tx_fifo	:	out	std_logic	:=	'0';
		pld_8g_full_tx_reg	:	out	std_logic	:=	'0';
		pld_8g_g3_tx_pld_rst_n_reg	:	out	std_logic	:=	'0';
		pld_8g_rddisable_tx_reg	:	out	std_logic	:=	'0';
		pld_8g_tx_boundary_sel_reg	:	out	std_logic	:=	'0';
		pld_pcs_tx_clk_out_8g_div_by_2_wire	:	out	std_logic	:=	'0';
		pld_pcs_tx_clk_out_8g_wire	:	out	std_logic	:=	'0';
		pld_tx_data_8g_fifo	:	out	std_logic	:=	'0';
		pld_tx_data_lo_8g_reg	:	out	std_logic	:=	'0';
		sta_tx_clk2_by2_1	:	out	std_logic	:=	'0';
		sta_tx_clk2_by2_1_out	:	out	std_logic	:=	'0';
		sta_tx_clk2_by4_1	:	out	std_logic	:=	'0';
		sta_tx_clk2_by4_1_out	:	out	std_logic	:=	'0';
		dyn_clk_switch_n	:	out	std_logic	:=	'0';
		ph_fifo_underflow	:	out	std_logic	:=	'0';
		fifo_select_out_chnl_down	:	out	std_logic_vector(1 downto 0)	:=	"00";
		fifo_select_out_chnl_up	:	out	std_logic_vector(1 downto 0)	:=	"00";
		ph_fifo_overflow	:	out	std_logic	:=	'0';
		g3_pipe_tx_pma_rstn	:	out	std_logic	:=	'0';
		g3_tx_pma_rstn	:	out	std_logic	:=	'0';
		non_gray_eidleinfersel	:	out	std_logic_vector(2 downto 0)	:=	"000";
		phfifo_txdeemph	:	out	std_logic	:=	'0';
		phfifo_txmargin	:	out	std_logic_vector(2 downto 0)	:=	"000";
		phfifo_txswing	:	out	std_logic	:=	'0';
		pipe_tx_clk_out_gen3	:	out	std_logic	:=	'0';
		pmaif_asn_rstn	:	out	std_logic	:=	'0';
		pipe_power_down_out	:	out	std_logic_vector(1 downto 0)	:=	"00";
		dataout	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		rd_enable_out_chnl_down	:	out	std_logic	:=	'0';
		rd_enable_out_chnl_up	:	out	std_logic	:=	'0';
		rd_ptr_tx_phfifo	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		refclk_b	:	out	std_logic	:=	'0';
		refclk_b_reset	:	out	std_logic	:=	'0';
		pipe_en_rev_parallel_lpbk_out	:	out	std_logic	:=	'0';
		rxpolarity_int	:	out	std_logic	:=	'0';
		soft_reset_wclk1_n	:	out	std_logic	:=	'0';
		sw_fifo_wr_clk	:	out	std_logic	:=	'0';
		tx_blk_start_out	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		clk_out	:	out	std_logic	:=	'0';
		tx_clk_out_8g_pmaif	:	out	std_logic	:=	'0';
		clk_out_gen3	:	out	std_logic	:=	'0';
		tx_clk_out_pld_if	:	out	std_logic	:=	'0';
		tx_clk_out_pmaif	:	out	std_logic	:=	'0';
		tx_clk_to_observation_ff_in_pld_if	:	out	std_logic	:=	'0';
		tx_ctrlplane_testbus	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		tx_data_out	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		tx_data_valid_out	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		tx_datak_out	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		tx_div_sync	:	out	std_logic_vector(1 downto 0)	:=	"00";
		tx_div_sync_out_chnl_down	:	out	std_logic_vector(1 downto 0)	:=	"00";
		tx_div_sync_out_chnl_up	:	out	std_logic_vector(1 downto 0)	:=	"00";
		tx_pipe_clk	:	out	std_logic	:=	'0';
		tx_pipe_electidle	:	out	std_logic	:=	'0';
		tx_pipe_soft_reset	:	out	std_logic	:=	'0';
		tx_sync_hdr_out	:	out	std_logic_vector(1 downto 0)	:=	"00";
		tx_testbus	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		txcompliance_out	:	out	std_logic	:=	'0';
		tx_detect_rxloopback_int	:	out	std_logic	:=	'0';
		txelecidle_out	:	out	std_logic	:=	'0';
		wr_clk_tx_phfifo_dw_clk	:	out	std_logic	:=	'0';
		wr_clk_tx_phfifo_sw_clk	:	out	std_logic	:=	'0';
		wr_data_tx_phfifo	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		wr_en_tx_phfifo	:	out	std_logic	:=	'0';
		wr_enable_out_chnl_down	:	out	std_logic	:=	'0';
		wr_enable_out_chnl_up	:	out	std_logic	:=	'0';
		wr_ptr_tx_phfifo	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		wr_rst_n_tx_phfifo	:	out	std_logic	:=	'0'
	);
end component;

begin



inst : twentynm_hssi_8g_tx_pcs_encrypted
	generic map (
		-- Instance parameters
		auto_speed_nego_gen2	=>	auto_speed_nego_gen2,
		bit_reversal	=>	bit_reversal,
		bonding_dft_en	=>	bonding_dft_en,
		bonding_dft_val	=>	bonding_dft_val,
		bypass_pipeline_reg	=>	bypass_pipeline_reg,
		byte_serializer	=>	byte_serializer,
		clock_gate_bs_enc	=>	clock_gate_bs_enc,
		clock_gate_dw_fifowr	=>	clock_gate_dw_fifowr,
		clock_gate_fiford	=>	clock_gate_fiford,
		clock_gate_sw_fifowr	=>	clock_gate_sw_fifowr,
		clock_observation_in_pld_core	=>	clock_observation_in_pld_core,
		ctrl_plane_bonding_compensation	=>	ctrl_plane_bonding_compensation,
		ctrl_plane_bonding_consumption	=>	ctrl_plane_bonding_consumption,
		ctrl_plane_bonding_distribution	=>	ctrl_plane_bonding_distribution,
		data_selection_8b10b_encoder_input	=>	data_selection_8b10b_encoder_input,
		dynamic_clk_switch	=>	dynamic_clk_switch,
		eightb_tenb_disp_ctrl	=>	eightb_tenb_disp_ctrl,
		eightb_tenb_encoder	=>	eightb_tenb_encoder,
		force_echar	=>	force_echar,
		force_kchar	=>	force_kchar,
		gen3_tx_clk_sel	=>	gen3_tx_clk_sel,
		gen3_tx_pipe_clk_sel	=>	gen3_tx_pipe_clk_sel,
		hip_mode	=>	hip_mode,
		pcs_bypass	=>	pcs_bypass,
		phase_comp_rdptr	=>	phase_comp_rdptr,
		phase_compensation_fifo	=>	phase_compensation_fifo,
		phfifo_write_clk_sel	=>	phfifo_write_clk_sel,
		pma_dw	=>	pma_dw,
		prot_mode	=>	prot_mode,
		reconfig_settings	=>	reconfig_settings,
		refclk_b_clk_sel	=>	refclk_b_clk_sel,
		revloop_back_rm	=>	revloop_back_rm,
		silicon_rev	=>	silicon_rev,
		sup_mode	=>	sup_mode,
		symbol_swap	=>	symbol_swap,
		tx_bitslip	=>	tx_bitslip,
		tx_compliance_controlled_disparity	=>	tx_compliance_controlled_disparity,
		tx_fast_pld_reg	=>	tx_fast_pld_reg,
		txclk_freerun	=>	txclk_freerun,
		txpcs_urst	=>	txpcs_urst
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		clk_sel_gen3	=>	clk_sel_gen3,
		dis_pc_byte	=>	dis_pc_byte,
		eidleinfersel	=>	eidleinfersel,
		fifo_select_in_chnl_down	=>	fifo_select_in_chnl_down,
		fifo_select_in_chnl_up	=>	fifo_select_in_chnl_up,
		rate_switch	=>	rate_switch,
		hrdrst	=>	hrdrst,
		pcs_rst	=>	pcs_rst,
		pipe_tx_deemph	=>	pipe_tx_deemph,
		pipe_tx_margin	=>	pipe_tx_margin,
		coreclk	=>	coreclk,
		powerdn	=>	powerdn,
		rd_data_tx_phfifo	=>	rd_data_tx_phfifo,
		rd_enable_in_chnl_down	=>	rd_enable_in_chnl_down,
		rd_enable_in_chnl_up	=>	rd_enable_in_chnl_up,
		ph_fifo_rd_disable	=>	ph_fifo_rd_disable,
		refclk_dig	=>	refclk_dig,
		reset_pc_ptrs	=>	reset_pc_ptrs,
		reset_pc_ptrs_in_chnl_down	=>	reset_pc_ptrs_in_chnl_down,
		reset_pc_ptrs_in_chnl_up	=>	reset_pc_ptrs_in_chnl_up,
		rev_parallel_lpbk_data	=>	rev_parallel_lpbk_data,
		en_rev_parallel_lpbk	=>	en_rev_parallel_lpbk,
		pipe_en_rev_parallel_lpbk_in	=>	pipe_en_rev_parallel_lpbk_in,
		rxpolarity	=>	rxpolarity,
		scan_mode_n	=>	scan_mode_n,
		tx_blk_start	=>	tx_blk_start,
		bitslip_boundary_select	=>	bitslip_boundary_select,
		tx_data_valid	=>	tx_data_valid,
		tx_div_sync_in_chnl_down	=>	tx_div_sync_in_chnl_down,
		tx_div_sync_in_chnl_up	=>	tx_div_sync_in_chnl_up,
		tx_sync_hdr	=>	tx_sync_hdr,
		datain	=>	datain,
		txd_fast_reg	=>	txd_fast_reg,
		detectrxloopin	=>	detectrxloopin,
		txpma_local_clk	=>	txpma_local_clk,
		txswing	=>	txswing,
		tx_pcs_reset	=>	tx_pcs_reset,
		wr_enable_in_chnl_down	=>	wr_enable_in_chnl_down,
		wr_enable_in_chnl_up	=>	wr_enable_in_chnl_up,
		wrenable_tx	=>	wrenable_tx,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		byte_serializer_pcs_clk_div_by_2_reg	=>	byte_serializer_pcs_clk_div_by_2_reg,
		byte_serializer_pcs_clk_div_by_2_wire	=>	byte_serializer_pcs_clk_div_by_2_wire,
		byte_serializer_pcs_clk_div_by_4_reg	=>	byte_serializer_pcs_clk_div_by_4_reg,
		byte_serializer_pld_clk_div_by_2_reg	=>	byte_serializer_pld_clk_div_by_2_reg,
		byte_serializer_pld_clk_div_by_4_reg	=>	byte_serializer_pld_clk_div_by_4_reg,
		pld_8g_empty_tx_fifo	=>	pld_8g_empty_tx_fifo,
		pld_8g_empty_tx_reg	=>	pld_8g_empty_tx_reg,
		pld_8g_full_tx_fifo	=>	pld_8g_full_tx_fifo,
		pld_8g_full_tx_reg	=>	pld_8g_full_tx_reg,
		pld_8g_g3_tx_pld_rst_n_reg	=>	pld_8g_g3_tx_pld_rst_n_reg,
		pld_8g_rddisable_tx_reg	=>	pld_8g_rddisable_tx_reg,
		pld_8g_tx_boundary_sel_reg	=>	pld_8g_tx_boundary_sel_reg,
		pld_pcs_tx_clk_out_8g_div_by_2_wire	=>	pld_pcs_tx_clk_out_8g_div_by_2_wire,
		pld_pcs_tx_clk_out_8g_wire	=>	pld_pcs_tx_clk_out_8g_wire,
		pld_tx_data_8g_fifo	=>	pld_tx_data_8g_fifo,
		pld_tx_data_lo_8g_reg	=>	pld_tx_data_lo_8g_reg,
		sta_tx_clk2_by2_1	=>	sta_tx_clk2_by2_1,
		sta_tx_clk2_by2_1_out	=>	sta_tx_clk2_by2_1_out,
		sta_tx_clk2_by4_1	=>	sta_tx_clk2_by4_1,
		sta_tx_clk2_by4_1_out	=>	sta_tx_clk2_by4_1_out,
		dyn_clk_switch_n	=>	dyn_clk_switch_n,
		ph_fifo_underflow	=>	ph_fifo_underflow,
		fifo_select_out_chnl_down	=>	fifo_select_out_chnl_down,
		fifo_select_out_chnl_up	=>	fifo_select_out_chnl_up,
		ph_fifo_overflow	=>	ph_fifo_overflow,
		g3_pipe_tx_pma_rstn	=>	g3_pipe_tx_pma_rstn,
		g3_tx_pma_rstn	=>	g3_tx_pma_rstn,
		non_gray_eidleinfersel	=>	non_gray_eidleinfersel,
		phfifo_txdeemph	=>	phfifo_txdeemph,
		phfifo_txmargin	=>	phfifo_txmargin,
		phfifo_txswing	=>	phfifo_txswing,
		pipe_tx_clk_out_gen3	=>	pipe_tx_clk_out_gen3,
		pmaif_asn_rstn	=>	pmaif_asn_rstn,
		pipe_power_down_out	=>	pipe_power_down_out,
		dataout	=>	dataout,
		rd_enable_out_chnl_down	=>	rd_enable_out_chnl_down,
		rd_enable_out_chnl_up	=>	rd_enable_out_chnl_up,
		rd_ptr_tx_phfifo	=>	rd_ptr_tx_phfifo,
		refclk_b	=>	refclk_b,
		refclk_b_reset	=>	refclk_b_reset,
		pipe_en_rev_parallel_lpbk_out	=>	pipe_en_rev_parallel_lpbk_out,
		rxpolarity_int	=>	rxpolarity_int,
		soft_reset_wclk1_n	=>	soft_reset_wclk1_n,
		sw_fifo_wr_clk	=>	sw_fifo_wr_clk,
		tx_blk_start_out	=>	tx_blk_start_out,
		clk_out	=>	clk_out,
		tx_clk_out_8g_pmaif	=>	tx_clk_out_8g_pmaif,
		clk_out_gen3	=>	clk_out_gen3,
		tx_clk_out_pld_if	=>	tx_clk_out_pld_if,
		tx_clk_out_pmaif	=>	tx_clk_out_pmaif,
		tx_clk_to_observation_ff_in_pld_if	=>	tx_clk_to_observation_ff_in_pld_if,
		tx_ctrlplane_testbus	=>	tx_ctrlplane_testbus,
		tx_data_out	=>	tx_data_out,
		tx_data_valid_out	=>	tx_data_valid_out,
		tx_datak_out	=>	tx_datak_out,
		tx_div_sync	=>	tx_div_sync,
		tx_div_sync_out_chnl_down	=>	tx_div_sync_out_chnl_down,
		tx_div_sync_out_chnl_up	=>	tx_div_sync_out_chnl_up,
		tx_pipe_clk	=>	tx_pipe_clk,
		tx_pipe_electidle	=>	tx_pipe_electidle,
		tx_pipe_soft_reset	=>	tx_pipe_soft_reset,
		tx_sync_hdr_out	=>	tx_sync_hdr_out,
		tx_testbus	=>	tx_testbus,
		txcompliance_out	=>	txcompliance_out,
		tx_detect_rxloopback_int	=>	tx_detect_rxloopback_int,
		txelecidle_out	=>	txelecidle_out,
		wr_clk_tx_phfifo_dw_clk	=>	wr_clk_tx_phfifo_dw_clk,
		wr_clk_tx_phfifo_sw_clk	=>	wr_clk_tx_phfifo_sw_clk,
		wr_data_tx_phfifo	=>	wr_data_tx_phfifo,
		wr_en_tx_phfifo	=>	wr_en_tx_phfifo,
		wr_enable_out_chnl_down	=>	wr_enable_out_chnl_down,
		wr_enable_out_chnl_up	=>	wr_enable_out_chnl_up,
		wr_ptr_tx_phfifo	=>	wr_ptr_tx_phfifo,
		wr_rst_n_tx_phfifo	=>	wr_rst_n_tx_phfifo
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_common_pcs_pma_interface	is
	generic (
		-- Entity parameters
		asn_clk_enable	:	string	:=	"false";
		asn_enable	:	string	:=	"dis_asn";
		block_sel	:	string	:=	"eight_g_pcs";
		bypass_early_eios	:	string	:=	"false";
		bypass_pcie_switch	:	string	:=	"false";
		bypass_pma_ltr	:	string	:=	"false";
		bypass_pma_sw_done	:	string	:=	"false";
		bypass_ppm_lock	:	string	:=	"false";
		bypass_send_syncp_fbkp	:	string	:=	"false";
		bypass_txdetectrx	:	string	:=	"false";
		cdr_control	:	string	:=	"en_cdr_ctrl";
		cid_enable	:	string	:=	"en_cid_mode";
		cp_cons_sel	:	string	:=	"cp_cons_default";
		cp_dwn_mstr	:	string	:=	"true";
		cp_up_mstr	:	string	:=	"true";
		ctrl_plane_bonding	:	string	:=	"individual";
		data_mask_count	:	bit_vector	:=	B"0000100111000100";
		data_mask_count_multi	:	bit_vector	:=	B"001";
		dft_observation_clock_selection	:	string	:=	"dft_clk_obsrv_tx0";
		early_eios_counter	:	bit_vector	:=	B"00110010";
		force_freqdet	:	string	:=	"force_freqdet_dis";
		free_run_clk_enable	:	string	:=	"true";
		ignore_sigdet_g23	:	string	:=	"false";
		pc_en_counter	:	bit_vector	:=	B"0110111";
		pc_rst_counter	:	bit_vector	:=	B"10111";
		pcie_hip_mode	:	string	:=	"hip_disable";
		ph_fifo_reg_mode	:	string	:=	"phfifo_reg_mode_dis";
		phfifo_flush_wait	:	bit_vector	:=	B"100100";
		pipe_if_g3pcs	:	string	:=	"pipe_if_8gpcs";
		pma_done_counter	:	bit_vector	:=	B"101010101110011000";
		pma_if_dft_en	:	string	:=	"dft_dis";
		pma_if_dft_val	:	string	:=	"dft_0";
		ppm_cnt_rst	:	string	:=	"ppm_cnt_rst_dis";
		ppm_deassert_early	:	string	:=	"deassert_early_dis";
		ppm_det_buckets	:	string	:=	"ppm_100_bucket";
		ppm_gen1_2_cnt	:	string	:=	"cnt_32k";
		ppm_post_eidle_delay	:	string	:=	"cnt_200_cycles";
		ppmsel	:	string	:=	"ppmsel_300";
		prot_mode	:	string	:=	"disable_prot_mode";
		reconfig_settings	:	string	:=	"{}";
		rxvalid_mask	:	string	:=	"rxvalid_mask_en";
		sigdet_wait_counter	:	bit_vector	:=	B"100111000100";
		sigdet_wait_counter_multi	:	bit_vector	:=	B"001";
		silicon_rev	:	string	:=	"20nm5es";
		sim_mode	:	string	:=	"disable";
		spd_chg_rst_wait_cnt_en	:	string	:=	"true";
		sup_mode	:	string	:=	"user_mode";
		testout_sel	:	string	:=	"ppm_det_test";
		wait_clk_on_off_timer	:	bit_vector	:=	B"0100";
		wait_pipe_synchronizing	:	bit_vector	:=	B"10111";
		wait_send_syncp_fbkp	:	bit_vector	:=	B"00011111010"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		int_pmaif_8g_current_coeff	:	in	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		int_pmaif_8g_eios_det	:	in	std_logic_vector(2 downto 0)	:=	"000";
		int_pmaif_8g_pipe_tx_pma_rstn	:	in	std_logic	:=	'0';
		int_pmaif_8g_rev_lpbk	:	in	std_logic	:=	'0';
		int_pmaif_8g_tx_clk_out_gen3	:	in	std_logic	:=	'0';
		int_pmaif_8g_txdetectrx	:	in	std_logic	:=	'0';
		int_pmaif_g3_eios_det	:	in	std_logic_vector(2 downto 0)	:=	"000";
		int_pmaif_g3_pma_current_coeff	:	in	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		int_pmaif_g3_pma_current_rxpreset	:	in	std_logic_vector(2 downto 0)	:=	"000";
		int_pmaif_g3_pma_txdetectrx	:	in	std_logic	:=	'0';
		int_pmaif_g3_rev_lpbk	:	in	std_logic	:=	'0';
		int_pmaif_pldif_8g_tx_pld_rstn	:	in	std_logic	:=	'0';
		int_pmaif_pldif_adapt_start	:	in	std_logic	:=	'0';
		int_pmaif_pldif_atpg_los_en_n	:	in	std_logic	:=	'0';
		int_pmaif_pldif_csr_test_dis	:	in	std_logic	:=	'0';
		int_pmaif_pldif_early_eios	:	in	std_logic	:=	'0';
		int_pmaif_pldif_interface_select	:	in	std_logic_vector(1 downto 0)	:=	"00";
		int_pmaif_pldif_ltd_b	:	in	std_logic	:=	'0';
		int_pmaif_pldif_ltr	:	in	std_logic	:=	'0';
		int_pmaif_pldif_nfrzdrv	:	in	std_logic	:=	'0';
		int_pmaif_pldif_nrpi_freeze	:	in	std_logic	:=	'0';
		int_pmaif_pldif_pcie_switch	:	in	std_logic_vector(1 downto 0)	:=	"00";
		int_pmaif_pldif_pma_reserved_out	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		int_pmaif_pldif_pma_scan_mode_n	:	in	std_logic	:=	'0';
		int_pmaif_pldif_pma_scan_shift_n	:	in	std_logic	:=	'0';
		int_pmaif_pldif_ppm_lock	:	in	std_logic	:=	'0';
		int_pmaif_pldif_rate	:	in	std_logic_vector(1 downto 0)	:=	"00";
		int_pmaif_pldif_refclk_dig	:	in	std_logic	:=	'0';
		int_pmaif_pldif_rs_lpbk_b	:	in	std_logic	:=	'0';
		int_pmaif_pldif_rx_qpi_pullup	:	in	std_logic	:=	'0';
		int_pmaif_pldif_rxpma_rstb	:	in	std_logic	:=	'0';
		int_pmaif_pldif_tx_bitslip	:	in	std_logic	:=	'0';
		int_pmaif_pldif_tx_bonding_rstb	:	in	std_logic	:=	'0';
		int_pmaif_pldif_tx_pma_syncp_hip	:	in	std_logic	:=	'0';
		int_pmaif_pldif_tx_qpi_pulldn	:	in	std_logic	:=	'0';
		int_pmaif_pldif_tx_qpi_pullup	:	in	std_logic	:=	'0';
		int_pmaif_pldif_txdetectrx	:	in	std_logic	:=	'0';
		int_pmaif_scan_mode_n	:	in	std_logic	:=	'0';
		int_rx_dft_obsrv_clk	:	in	std_logic	:=	'0';
		int_tx_dft_obsrv_clk	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		iocsr_clk	:	in	std_logic	:=	'0';
		iocsr_config	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		iocsr_rdy	:	in	std_logic	:=	'0';
		iocsr_rdy_dly	:	in	std_logic	:=	'0';
		pma_adapt_done	:	in	std_logic	:=	'0';
		pma_clklow	:	in	std_logic	:=	'0';
		pma_fref	:	in	std_logic	:=	'0';
		pma_hclk	:	in	std_logic	:=	'0';
		pma_pcie_sw_done	:	in	std_logic_vector(1 downto 0)	:=	"00";
		pma_pfdmode_lock	:	in	std_logic	:=	'0';
		pma_reserved_in	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		pma_signal_det	:	in	std_logic	:=	'0';
		pma_testbus	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		pmaif_bundling_in_down	:	in	std_logic_vector(11 downto 0)	:=	"000000000000";
		pmaif_bundling_in_up	:	in	std_logic_vector(11 downto 0)	:=	"000000000000";
		rx_pmaif_test_out	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		rx_prbs_ver_test	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		tx_prbs_gen_test	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		uhsif_test_out_1	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		uhsif_test_out_2	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		uhsif_test_out_3	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		sta_pma_hclk_by2	:	out	std_logic	:=	'0';
		int_pmaif_8g_asn_bundling_in	:	out	std_logic_vector(8 downto 0)	:=	"000000000";
		int_pmaif_8g_eios_detected	:	out	std_logic	:=	'0';
		int_pmaif_8g_inferred_rxvalid	:	out	std_logic	:=	'0';
		int_pmaif_8g_power_state_transition_done	:	out	std_logic	:=	'0';
		int_pmaif_avmm_iocsr_clk	:	out	std_logic	:=	'0';
		int_pmaif_avmm_iocsr_config	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		int_pmaif_avmm_iocsr_rdy	:	out	std_logic	:=	'0';
		int_pmaif_avmm_iocsr_rdy_dly	:	out	std_logic	:=	'0';
		int_pmaif_g3_data_sel	:	out	std_logic	:=	'0';
		int_pmaif_g3_inferred_rxvalid	:	out	std_logic	:=	'0';
		int_pmaif_g3_pcs_asn_bundling_in	:	out	std_logic_vector(8 downto 0)	:=	"000000000";
		int_pmaif_pldif_adapt_done	:	out	std_logic	:=	'0';
		int_pmaif_pldif_dft_obsrv_clk	:	out	std_logic	:=	'0';
		int_pmaif_pldif_mask_tx_pll	:	out	std_logic	:=	'0';
		int_pmaif_pldif_pcie_sw_done	:	out	std_logic_vector(1 downto 0)	:=	"00";
		int_pmaif_pldif_pfdmode_lock	:	out	std_logic	:=	'0';
		int_pmaif_pldif_pma_clklow	:	out	std_logic	:=	'0';
		int_pmaif_pldif_pma_fref	:	out	std_logic	:=	'0';
		int_pmaif_pldif_pma_hclk	:	out	std_logic	:=	'0';
		int_pmaif_pldif_pma_reserved_in	:	out	std_logic_vector(4 downto 0)	:=	"00000";
		int_pmaif_pldif_test_out	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		int_pmaif_pldif_testbus	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		pma_adapt_start	:	out	std_logic	:=	'0';
		pma_atpg_los_en_n	:	out	std_logic	:=	'0';
		pma_csr_test_dis	:	out	std_logic	:=	'0';
		pma_current_coeff	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		pma_current_rxpreset	:	out	std_logic_vector(2 downto 0)	:=	"000";
		pma_early_eios	:	out	std_logic	:=	'0';
		pma_interface_select	:	out	std_logic_vector(1 downto 0)	:=	"00";
		pma_ltd_b	:	out	std_logic	:=	'0';
		pma_ltr	:	out	std_logic	:=	'0';
		pma_nfrzdrv	:	out	std_logic	:=	'0';
		pma_nrpi_freeze	:	out	std_logic	:=	'0';
		pma_pcie_switch	:	out	std_logic_vector(1 downto 0)	:=	"00";
		pma_ppm_lock	:	out	std_logic	:=	'0';
		pma_reserved_out	:	out	std_logic_vector(4 downto 0)	:=	"00000";
		pma_rs_lpbk_b	:	out	std_logic	:=	'0';
		pma_rx_qpi_pullup	:	out	std_logic	:=	'0';
		pma_scan_mode_n	:	out	std_logic	:=	'0';
		pma_scan_shift_n	:	out	std_logic	:=	'0';
		pma_tx_bitslip	:	out	std_logic	:=	'0';
		pma_tx_bonding_rstb	:	out	std_logic	:=	'0';
		pma_tx_pma_syncp	:	out	std_logic	:=	'0';
		pma_tx_qpi_pulldn	:	out	std_logic	:=	'0';
		pma_tx_qpi_pullup	:	out	std_logic	:=	'0';
		pma_tx_txdetectrx	:	out	std_logic	:=	'0';
		pmaif_bundling_out_down	:	out	std_logic_vector(11 downto 0)	:=	"000000000000";
		pmaif_bundling_out_up	:	out	std_logic_vector(11 downto 0)	:=	"000000000000"
	);
end twentynm_hssi_common_pcs_pma_interface;

architecture behavior of twentynm_hssi_common_pcs_pma_interface	is

constant data_mask_count_int	:	integer	:=	bin2int(data_mask_count);
constant data_mask_count_multi_int	:	integer	:=	bin2int(data_mask_count_multi);
constant early_eios_counter_int	:	integer	:=	bin2int(early_eios_counter);
constant pc_en_counter_int	:	integer	:=	bin2int(pc_en_counter);
constant pc_rst_counter_int	:	integer	:=	bin2int(pc_rst_counter);
constant phfifo_flush_wait_int	:	integer	:=	bin2int(phfifo_flush_wait);
constant pma_done_counter_int	:	integer	:=	bin2int(pma_done_counter);
constant sigdet_wait_counter_int	:	integer	:=	bin2int(sigdet_wait_counter);
constant sigdet_wait_counter_multi_int	:	integer	:=	bin2int(sigdet_wait_counter_multi);
constant wait_clk_on_off_timer_int	:	integer	:=	bin2int(wait_clk_on_off_timer);
constant wait_pipe_synchronizing_int	:	integer	:=	bin2int(wait_pipe_synchronizing);
constant wait_send_syncp_fbkp_int	:	integer	:=	bin2int(wait_send_syncp_fbkp);



component	twentynm_hssi_common_pcs_pma_interface_encrypted
	generic (
		-- Architecture parameters
		asn_clk_enable	:	string	:=	"false";
		asn_enable	:	string	:=	"dis_asn";
		block_sel	:	string	:=	"eight_g_pcs";
		bypass_early_eios	:	string	:=	"false";
		bypass_pcie_switch	:	string	:=	"false";
		bypass_pma_ltr	:	string	:=	"false";
		bypass_pma_sw_done	:	string	:=	"false";
		bypass_ppm_lock	:	string	:=	"false";
		bypass_send_syncp_fbkp	:	string	:=	"false";
		bypass_txdetectrx	:	string	:=	"false";
		cdr_control	:	string	:=	"en_cdr_ctrl";
		cid_enable	:	string	:=	"en_cid_mode";
		cp_cons_sel	:	string	:=	"cp_cons_default";
		cp_dwn_mstr	:	string	:=	"true";
		cp_up_mstr	:	string	:=	"true";
		ctrl_plane_bonding	:	string	:=	"individual";
		data_mask_count	:	integer	:=	2500;
		data_mask_count_multi	:	integer	:=	1;
		dft_observation_clock_selection	:	string	:=	"dft_clk_obsrv_tx0";
		early_eios_counter	:	integer	:=	50;
		force_freqdet	:	string	:=	"force_freqdet_dis";
		free_run_clk_enable	:	string	:=	"true";
		ignore_sigdet_g23	:	string	:=	"false";
		pc_en_counter	:	integer	:=	55;
		pc_rst_counter	:	integer	:=	23;
		pcie_hip_mode	:	string	:=	"hip_disable";
		ph_fifo_reg_mode	:	string	:=	"phfifo_reg_mode_dis";
		phfifo_flush_wait	:	integer	:=	36;
		pipe_if_g3pcs	:	string	:=	"pipe_if_8gpcs";
		pma_done_counter	:	integer	:=	175000;
		pma_if_dft_en	:	string	:=	"dft_dis";
		pma_if_dft_val	:	string	:=	"dft_0";
		ppm_cnt_rst	:	string	:=	"ppm_cnt_rst_dis";
		ppm_deassert_early	:	string	:=	"deassert_early_dis";
		ppm_det_buckets	:	string	:=	"ppm_100_bucket";
		ppm_gen1_2_cnt	:	string	:=	"cnt_32k";
		ppm_post_eidle_delay	:	string	:=	"cnt_200_cycles";
		ppmsel	:	string	:=	"ppmsel_300";
		prot_mode	:	string	:=	"disable_prot_mode";
		reconfig_settings	:	string	:=	"{}";
		rxvalid_mask	:	string	:=	"rxvalid_mask_en";
		sigdet_wait_counter	:	integer	:=	2500;
		sigdet_wait_counter_multi	:	integer	:=	1;
		silicon_rev	:	string	:=	"20nm5es";
		sim_mode	:	string	:=	"disable";
		spd_chg_rst_wait_cnt_en	:	string	:=	"true";
		sup_mode	:	string	:=	"user_mode";
		testout_sel	:	string	:=	"ppm_det_test";
		wait_clk_on_off_timer	:	integer	:=	4;
		wait_pipe_synchronizing	:	integer	:=	23;
		wait_send_syncp_fbkp	:	integer	:=	250
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		int_pmaif_8g_current_coeff	:	in	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		int_pmaif_8g_eios_det	:	in	std_logic_vector(2 downto 0)	:=	"000";
		int_pmaif_8g_pipe_tx_pma_rstn	:	in	std_logic	:=	'0';
		int_pmaif_8g_rev_lpbk	:	in	std_logic	:=	'0';
		int_pmaif_8g_tx_clk_out_gen3	:	in	std_logic	:=	'0';
		int_pmaif_8g_txdetectrx	:	in	std_logic	:=	'0';
		int_pmaif_g3_eios_det	:	in	std_logic_vector(2 downto 0)	:=	"000";
		int_pmaif_g3_pma_current_coeff	:	in	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		int_pmaif_g3_pma_current_rxpreset	:	in	std_logic_vector(2 downto 0)	:=	"000";
		int_pmaif_g3_pma_txdetectrx	:	in	std_logic	:=	'0';
		int_pmaif_g3_rev_lpbk	:	in	std_logic	:=	'0';
		int_pmaif_pldif_8g_tx_pld_rstn	:	in	std_logic	:=	'0';
		int_pmaif_pldif_adapt_start	:	in	std_logic	:=	'0';
		int_pmaif_pldif_atpg_los_en_n	:	in	std_logic	:=	'0';
		int_pmaif_pldif_csr_test_dis	:	in	std_logic	:=	'0';
		int_pmaif_pldif_early_eios	:	in	std_logic	:=	'0';
		int_pmaif_pldif_interface_select	:	in	std_logic_vector(1 downto 0)	:=	"00";
		int_pmaif_pldif_ltd_b	:	in	std_logic	:=	'0';
		int_pmaif_pldif_ltr	:	in	std_logic	:=	'0';
		int_pmaif_pldif_nfrzdrv	:	in	std_logic	:=	'0';
		int_pmaif_pldif_nrpi_freeze	:	in	std_logic	:=	'0';
		int_pmaif_pldif_pcie_switch	:	in	std_logic_vector(1 downto 0)	:=	"00";
		int_pmaif_pldif_pma_reserved_out	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		int_pmaif_pldif_pma_scan_mode_n	:	in	std_logic	:=	'0';
		int_pmaif_pldif_pma_scan_shift_n	:	in	std_logic	:=	'0';
		int_pmaif_pldif_ppm_lock	:	in	std_logic	:=	'0';
		int_pmaif_pldif_rate	:	in	std_logic_vector(1 downto 0)	:=	"00";
		int_pmaif_pldif_refclk_dig	:	in	std_logic	:=	'0';
		int_pmaif_pldif_rs_lpbk_b	:	in	std_logic	:=	'0';
		int_pmaif_pldif_rx_qpi_pullup	:	in	std_logic	:=	'0';
		int_pmaif_pldif_rxpma_rstb	:	in	std_logic	:=	'0';
		int_pmaif_pldif_tx_bitslip	:	in	std_logic	:=	'0';
		int_pmaif_pldif_tx_bonding_rstb	:	in	std_logic	:=	'0';
		int_pmaif_pldif_tx_pma_syncp_hip	:	in	std_logic	:=	'0';
		int_pmaif_pldif_tx_qpi_pulldn	:	in	std_logic	:=	'0';
		int_pmaif_pldif_tx_qpi_pullup	:	in	std_logic	:=	'0';
		int_pmaif_pldif_txdetectrx	:	in	std_logic	:=	'0';
		int_pmaif_scan_mode_n	:	in	std_logic	:=	'0';
		int_rx_dft_obsrv_clk	:	in	std_logic	:=	'0';
		int_tx_dft_obsrv_clk	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		iocsr_clk	:	in	std_logic	:=	'0';
		iocsr_config	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		iocsr_rdy	:	in	std_logic	:=	'0';
		iocsr_rdy_dly	:	in	std_logic	:=	'0';
		pma_adapt_done	:	in	std_logic	:=	'0';
		pma_clklow	:	in	std_logic	:=	'0';
		pma_fref	:	in	std_logic	:=	'0';
		pma_hclk	:	in	std_logic	:=	'0';
		pma_pcie_sw_done	:	in	std_logic_vector(1 downto 0)	:=	"00";
		pma_pfdmode_lock	:	in	std_logic	:=	'0';
		pma_reserved_in	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		pma_signal_det	:	in	std_logic	:=	'0';
		pma_testbus	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		pmaif_bundling_in_down	:	in	std_logic_vector(11 downto 0)	:=	"000000000000";
		pmaif_bundling_in_up	:	in	std_logic_vector(11 downto 0)	:=	"000000000000";
		rx_pmaif_test_out	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		rx_prbs_ver_test	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		tx_prbs_gen_test	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		uhsif_test_out_1	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		uhsif_test_out_2	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		uhsif_test_out_3	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		sta_pma_hclk_by2	:	out	std_logic	:=	'0';
		int_pmaif_8g_asn_bundling_in	:	out	std_logic_vector(8 downto 0)	:=	"000000000";
		int_pmaif_8g_eios_detected	:	out	std_logic	:=	'0';
		int_pmaif_8g_inferred_rxvalid	:	out	std_logic	:=	'0';
		int_pmaif_8g_power_state_transition_done	:	out	std_logic	:=	'0';
		int_pmaif_avmm_iocsr_clk	:	out	std_logic	:=	'0';
		int_pmaif_avmm_iocsr_config	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		int_pmaif_avmm_iocsr_rdy	:	out	std_logic	:=	'0';
		int_pmaif_avmm_iocsr_rdy_dly	:	out	std_logic	:=	'0';
		int_pmaif_g3_data_sel	:	out	std_logic	:=	'0';
		int_pmaif_g3_inferred_rxvalid	:	out	std_logic	:=	'0';
		int_pmaif_g3_pcs_asn_bundling_in	:	out	std_logic_vector(8 downto 0)	:=	"000000000";
		int_pmaif_pldif_adapt_done	:	out	std_logic	:=	'0';
		int_pmaif_pldif_dft_obsrv_clk	:	out	std_logic	:=	'0';
		int_pmaif_pldif_mask_tx_pll	:	out	std_logic	:=	'0';
		int_pmaif_pldif_pcie_sw_done	:	out	std_logic_vector(1 downto 0)	:=	"00";
		int_pmaif_pldif_pfdmode_lock	:	out	std_logic	:=	'0';
		int_pmaif_pldif_pma_clklow	:	out	std_logic	:=	'0';
		int_pmaif_pldif_pma_fref	:	out	std_logic	:=	'0';
		int_pmaif_pldif_pma_hclk	:	out	std_logic	:=	'0';
		int_pmaif_pldif_pma_reserved_in	:	out	std_logic_vector(4 downto 0)	:=	"00000";
		int_pmaif_pldif_test_out	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		int_pmaif_pldif_testbus	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		pma_adapt_start	:	out	std_logic	:=	'0';
		pma_atpg_los_en_n	:	out	std_logic	:=	'0';
		pma_csr_test_dis	:	out	std_logic	:=	'0';
		pma_current_coeff	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		pma_current_rxpreset	:	out	std_logic_vector(2 downto 0)	:=	"000";
		pma_early_eios	:	out	std_logic	:=	'0';
		pma_interface_select	:	out	std_logic_vector(1 downto 0)	:=	"00";
		pma_ltd_b	:	out	std_logic	:=	'0';
		pma_ltr	:	out	std_logic	:=	'0';
		pma_nfrzdrv	:	out	std_logic	:=	'0';
		pma_nrpi_freeze	:	out	std_logic	:=	'0';
		pma_pcie_switch	:	out	std_logic_vector(1 downto 0)	:=	"00";
		pma_ppm_lock	:	out	std_logic	:=	'0';
		pma_reserved_out	:	out	std_logic_vector(4 downto 0)	:=	"00000";
		pma_rs_lpbk_b	:	out	std_logic	:=	'0';
		pma_rx_qpi_pullup	:	out	std_logic	:=	'0';
		pma_scan_mode_n	:	out	std_logic	:=	'0';
		pma_scan_shift_n	:	out	std_logic	:=	'0';
		pma_tx_bitslip	:	out	std_logic	:=	'0';
		pma_tx_bonding_rstb	:	out	std_logic	:=	'0';
		pma_tx_pma_syncp	:	out	std_logic	:=	'0';
		pma_tx_qpi_pulldn	:	out	std_logic	:=	'0';
		pma_tx_qpi_pullup	:	out	std_logic	:=	'0';
		pma_tx_txdetectrx	:	out	std_logic	:=	'0';
		pmaif_bundling_out_down	:	out	std_logic_vector(11 downto 0)	:=	"000000000000";
		pmaif_bundling_out_up	:	out	std_logic_vector(11 downto 0)	:=	"000000000000"
	);
end component;

begin



inst : twentynm_hssi_common_pcs_pma_interface_encrypted
	generic map (
		-- Instance parameters
		asn_clk_enable	=>	asn_clk_enable,
		asn_enable	=>	asn_enable,
		block_sel	=>	block_sel,
		bypass_early_eios	=>	bypass_early_eios,
		bypass_pcie_switch	=>	bypass_pcie_switch,
		bypass_pma_ltr	=>	bypass_pma_ltr,
		bypass_pma_sw_done	=>	bypass_pma_sw_done,
		bypass_ppm_lock	=>	bypass_ppm_lock,
		bypass_send_syncp_fbkp	=>	bypass_send_syncp_fbkp,
		bypass_txdetectrx	=>	bypass_txdetectrx,
		cdr_control	=>	cdr_control,
		cid_enable	=>	cid_enable,
		cp_cons_sel	=>	cp_cons_sel,
		cp_dwn_mstr	=>	cp_dwn_mstr,
		cp_up_mstr	=>	cp_up_mstr,
		ctrl_plane_bonding	=>	ctrl_plane_bonding,
		data_mask_count	=>	data_mask_count_int,
		data_mask_count_multi	=>	data_mask_count_multi_int,
		dft_observation_clock_selection	=>	dft_observation_clock_selection,
		early_eios_counter	=>	early_eios_counter_int,
		force_freqdet	=>	force_freqdet,
		free_run_clk_enable	=>	free_run_clk_enable,
		ignore_sigdet_g23	=>	ignore_sigdet_g23,
		pc_en_counter	=>	pc_en_counter_int,
		pc_rst_counter	=>	pc_rst_counter_int,
		pcie_hip_mode	=>	pcie_hip_mode,
		ph_fifo_reg_mode	=>	ph_fifo_reg_mode,
		phfifo_flush_wait	=>	phfifo_flush_wait_int,
		pipe_if_g3pcs	=>	pipe_if_g3pcs,
		pma_done_counter	=>	pma_done_counter_int,
		pma_if_dft_en	=>	pma_if_dft_en,
		pma_if_dft_val	=>	pma_if_dft_val,
		ppm_cnt_rst	=>	ppm_cnt_rst,
		ppm_deassert_early	=>	ppm_deassert_early,
		ppm_det_buckets	=>	ppm_det_buckets,
		ppm_gen1_2_cnt	=>	ppm_gen1_2_cnt,
		ppm_post_eidle_delay	=>	ppm_post_eidle_delay,
		ppmsel	=>	ppmsel,
		prot_mode	=>	prot_mode,
		reconfig_settings	=>	reconfig_settings,
		rxvalid_mask	=>	rxvalid_mask,
		sigdet_wait_counter	=>	sigdet_wait_counter_int,
		sigdet_wait_counter_multi	=>	sigdet_wait_counter_multi_int,
		silicon_rev	=>	silicon_rev,
		sim_mode	=>	sim_mode,
		spd_chg_rst_wait_cnt_en	=>	spd_chg_rst_wait_cnt_en,
		sup_mode	=>	sup_mode,
		testout_sel	=>	testout_sel,
		wait_clk_on_off_timer	=>	wait_clk_on_off_timer_int,
		wait_pipe_synchronizing	=>	wait_pipe_synchronizing_int,
		wait_send_syncp_fbkp	=>	wait_send_syncp_fbkp_int
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		int_pmaif_8g_current_coeff	=>	int_pmaif_8g_current_coeff,
		int_pmaif_8g_eios_det	=>	int_pmaif_8g_eios_det,
		int_pmaif_8g_pipe_tx_pma_rstn	=>	int_pmaif_8g_pipe_tx_pma_rstn,
		int_pmaif_8g_rev_lpbk	=>	int_pmaif_8g_rev_lpbk,
		int_pmaif_8g_tx_clk_out_gen3	=>	int_pmaif_8g_tx_clk_out_gen3,
		int_pmaif_8g_txdetectrx	=>	int_pmaif_8g_txdetectrx,
		int_pmaif_g3_eios_det	=>	int_pmaif_g3_eios_det,
		int_pmaif_g3_pma_current_coeff	=>	int_pmaif_g3_pma_current_coeff,
		int_pmaif_g3_pma_current_rxpreset	=>	int_pmaif_g3_pma_current_rxpreset,
		int_pmaif_g3_pma_txdetectrx	=>	int_pmaif_g3_pma_txdetectrx,
		int_pmaif_g3_rev_lpbk	=>	int_pmaif_g3_rev_lpbk,
		int_pmaif_pldif_8g_tx_pld_rstn	=>	int_pmaif_pldif_8g_tx_pld_rstn,
		int_pmaif_pldif_adapt_start	=>	int_pmaif_pldif_adapt_start,
		int_pmaif_pldif_atpg_los_en_n	=>	int_pmaif_pldif_atpg_los_en_n,
		int_pmaif_pldif_csr_test_dis	=>	int_pmaif_pldif_csr_test_dis,
		int_pmaif_pldif_early_eios	=>	int_pmaif_pldif_early_eios,
		int_pmaif_pldif_interface_select	=>	int_pmaif_pldif_interface_select,
		int_pmaif_pldif_ltd_b	=>	int_pmaif_pldif_ltd_b,
		int_pmaif_pldif_ltr	=>	int_pmaif_pldif_ltr,
		int_pmaif_pldif_nfrzdrv	=>	int_pmaif_pldif_nfrzdrv,
		int_pmaif_pldif_nrpi_freeze	=>	int_pmaif_pldif_nrpi_freeze,
		int_pmaif_pldif_pcie_switch	=>	int_pmaif_pldif_pcie_switch,
		int_pmaif_pldif_pma_reserved_out	=>	int_pmaif_pldif_pma_reserved_out,
		int_pmaif_pldif_pma_scan_mode_n	=>	int_pmaif_pldif_pma_scan_mode_n,
		int_pmaif_pldif_pma_scan_shift_n	=>	int_pmaif_pldif_pma_scan_shift_n,
		int_pmaif_pldif_ppm_lock	=>	int_pmaif_pldif_ppm_lock,
		int_pmaif_pldif_rate	=>	int_pmaif_pldif_rate,
		int_pmaif_pldif_refclk_dig	=>	int_pmaif_pldif_refclk_dig,
		int_pmaif_pldif_rs_lpbk_b	=>	int_pmaif_pldif_rs_lpbk_b,
		int_pmaif_pldif_rx_qpi_pullup	=>	int_pmaif_pldif_rx_qpi_pullup,
		int_pmaif_pldif_rxpma_rstb	=>	int_pmaif_pldif_rxpma_rstb,
		int_pmaif_pldif_tx_bitslip	=>	int_pmaif_pldif_tx_bitslip,
		int_pmaif_pldif_tx_bonding_rstb	=>	int_pmaif_pldif_tx_bonding_rstb,
		int_pmaif_pldif_tx_pma_syncp_hip	=>	int_pmaif_pldif_tx_pma_syncp_hip,
		int_pmaif_pldif_tx_qpi_pulldn	=>	int_pmaif_pldif_tx_qpi_pulldn,
		int_pmaif_pldif_tx_qpi_pullup	=>	int_pmaif_pldif_tx_qpi_pullup,
		int_pmaif_pldif_txdetectrx	=>	int_pmaif_pldif_txdetectrx,
		int_pmaif_scan_mode_n	=>	int_pmaif_scan_mode_n,
		int_rx_dft_obsrv_clk	=>	int_rx_dft_obsrv_clk,
		int_tx_dft_obsrv_clk	=>	int_tx_dft_obsrv_clk,
		iocsr_clk	=>	iocsr_clk,
		iocsr_config	=>	iocsr_config,
		iocsr_rdy	=>	iocsr_rdy,
		iocsr_rdy_dly	=>	iocsr_rdy_dly,
		pma_adapt_done	=>	pma_adapt_done,
		pma_clklow	=>	pma_clklow,
		pma_fref	=>	pma_fref,
		pma_hclk	=>	pma_hclk,
		pma_pcie_sw_done	=>	pma_pcie_sw_done,
		pma_pfdmode_lock	=>	pma_pfdmode_lock,
		pma_reserved_in	=>	pma_reserved_in,
		pma_signal_det	=>	pma_signal_det,
		pma_testbus	=>	pma_testbus,
		pmaif_bundling_in_down	=>	pmaif_bundling_in_down,
		pmaif_bundling_in_up	=>	pmaif_bundling_in_up,
		rx_pmaif_test_out	=>	rx_pmaif_test_out,
		rx_prbs_ver_test	=>	rx_prbs_ver_test,
		tx_prbs_gen_test	=>	tx_prbs_gen_test,
		uhsif_test_out_1	=>	uhsif_test_out_1,
		uhsif_test_out_2	=>	uhsif_test_out_2,
		uhsif_test_out_3	=>	uhsif_test_out_3,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		sta_pma_hclk_by2	=>	sta_pma_hclk_by2,
		int_pmaif_8g_asn_bundling_in	=>	int_pmaif_8g_asn_bundling_in,
		int_pmaif_8g_eios_detected	=>	int_pmaif_8g_eios_detected,
		int_pmaif_8g_inferred_rxvalid	=>	int_pmaif_8g_inferred_rxvalid,
		int_pmaif_8g_power_state_transition_done	=>	int_pmaif_8g_power_state_transition_done,
		int_pmaif_avmm_iocsr_clk	=>	int_pmaif_avmm_iocsr_clk,
		int_pmaif_avmm_iocsr_config	=>	int_pmaif_avmm_iocsr_config,
		int_pmaif_avmm_iocsr_rdy	=>	int_pmaif_avmm_iocsr_rdy,
		int_pmaif_avmm_iocsr_rdy_dly	=>	int_pmaif_avmm_iocsr_rdy_dly,
		int_pmaif_g3_data_sel	=>	int_pmaif_g3_data_sel,
		int_pmaif_g3_inferred_rxvalid	=>	int_pmaif_g3_inferred_rxvalid,
		int_pmaif_g3_pcs_asn_bundling_in	=>	int_pmaif_g3_pcs_asn_bundling_in,
		int_pmaif_pldif_adapt_done	=>	int_pmaif_pldif_adapt_done,
		int_pmaif_pldif_dft_obsrv_clk	=>	int_pmaif_pldif_dft_obsrv_clk,
		int_pmaif_pldif_mask_tx_pll	=>	int_pmaif_pldif_mask_tx_pll,
		int_pmaif_pldif_pcie_sw_done	=>	int_pmaif_pldif_pcie_sw_done,
		int_pmaif_pldif_pfdmode_lock	=>	int_pmaif_pldif_pfdmode_lock,
		int_pmaif_pldif_pma_clklow	=>	int_pmaif_pldif_pma_clklow,
		int_pmaif_pldif_pma_fref	=>	int_pmaif_pldif_pma_fref,
		int_pmaif_pldif_pma_hclk	=>	int_pmaif_pldif_pma_hclk,
		int_pmaif_pldif_pma_reserved_in	=>	int_pmaif_pldif_pma_reserved_in,
		int_pmaif_pldif_test_out	=>	int_pmaif_pldif_test_out,
		int_pmaif_pldif_testbus	=>	int_pmaif_pldif_testbus,
		pma_adapt_start	=>	pma_adapt_start,
		pma_atpg_los_en_n	=>	pma_atpg_los_en_n,
		pma_csr_test_dis	=>	pma_csr_test_dis,
		pma_current_coeff	=>	pma_current_coeff,
		pma_current_rxpreset	=>	pma_current_rxpreset,
		pma_early_eios	=>	pma_early_eios,
		pma_interface_select	=>	pma_interface_select,
		pma_ltd_b	=>	pma_ltd_b,
		pma_ltr	=>	pma_ltr,
		pma_nfrzdrv	=>	pma_nfrzdrv,
		pma_nrpi_freeze	=>	pma_nrpi_freeze,
		pma_pcie_switch	=>	pma_pcie_switch,
		pma_ppm_lock	=>	pma_ppm_lock,
		pma_reserved_out	=>	pma_reserved_out,
		pma_rs_lpbk_b	=>	pma_rs_lpbk_b,
		pma_rx_qpi_pullup	=>	pma_rx_qpi_pullup,
		pma_scan_mode_n	=>	pma_scan_mode_n,
		pma_scan_shift_n	=>	pma_scan_shift_n,
		pma_tx_bitslip	=>	pma_tx_bitslip,
		pma_tx_bonding_rstb	=>	pma_tx_bonding_rstb,
		pma_tx_pma_syncp	=>	pma_tx_pma_syncp,
		pma_tx_qpi_pulldn	=>	pma_tx_qpi_pulldn,
		pma_tx_qpi_pullup	=>	pma_tx_qpi_pullup,
		pma_tx_txdetectrx	=>	pma_tx_txdetectrx,
		pmaif_bundling_out_down	=>	pmaif_bundling_out_down,
		pmaif_bundling_out_up	=>	pmaif_bundling_out_up
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_common_pld_pcs_interface	is
	generic (
		-- Entity parameters
		dft_clk_out_en	:	string	:=	"dft_clk_out_disable";
		dft_clk_out_sel	:	string	:=	"teng_rx_dft_clk";
		hrdrstctrl_en	:	string	:=	"hrst_dis";
		pcs_testbus_block_sel	:	string	:=	"eightg";
		reconfig_settings	:	string	:=	"{}";
		silicon_rev	:	string	:=	"20nm5es"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		int_pldif_10g_rx_dft_clk_out	:	in	std_logic	:=	'0';
		int_pldif_10g_test_data	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		int_pldif_10g_tx_dft_clk_out	:	in	std_logic	:=	'0';
		int_pldif_8g_chnl_test_bus_out	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		int_pldif_8g_rx_clk_to_observation_ff_in_pld_if	:	in	std_logic	:=	'0';
		int_pldif_8g_tx_clk_to_observation_ff_in_pld_if	:	in	std_logic	:=	'0';
		int_pldif_avmm_refclk_dig_en	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		int_pldif_g3_test_out	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		int_pldif_krfec_test_data	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		int_pldif_pmaif_adapt_done	:	in	std_logic	:=	'0';
		int_pldif_pmaif_mask_tx_pll	:	in	std_logic	:=	'0';
		int_pldif_pmaif_pcie_sw_done	:	in	std_logic_vector(1 downto 0)	:=	"00";
		int_pldif_pmaif_pfdmode_lock	:	in	std_logic	:=	'0';
		int_pldif_pmaif_pma_clklow	:	in	std_logic	:=	'0';
		int_pldif_pmaif_pma_fref	:	in	std_logic	:=	'0';
		int_pldif_pmaif_pma_hclk	:	in	std_logic	:=	'0';
		int_pldif_pmaif_pma_reserved_in	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		int_pldif_pmaif_rx_detect_valid	:	in	std_logic	:=	'0';
		int_pldif_pmaif_rx_found	:	in	std_logic	:=	'0';
		int_pldif_pmaif_rxpll_lock	:	in	std_logic	:=	'0';
		int_pldif_pmaif_test_out	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		int_pldif_pmaif_testbus	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		int_pldif_pmaif_uhsif_lock	:	in	std_logic	:=	'0';
		int_pmaif_pldif_dft_obsrv_clk	:	in	std_logic	:=	'0';
		int_pmaif_pldif_uhsif_scan_chain_out	:	in	std_logic	:=	'0';
		pld_8g_eidleinfersel	:	in	std_logic_vector(2 downto 0)	:=	"000";
		pld_8g_refclk_dig2	:	in	std_logic	:=	'0';
		pld_atpg_los_en_n	:	in	std_logic	:=	'0';
		pld_g3_current_coeff	:	in	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		pld_g3_current_rxpreset	:	in	std_logic_vector(2 downto 0)	:=	"000";
		pld_ltr	:	in	std_logic	:=	'0';
		pld_mem_krfec_atpg_rst_n	:	in	std_logic	:=	'0';
		pld_partial_reconfig	:	in	std_logic	:=	'0';
		pld_pcs_refclk_dig	:	in	std_logic	:=	'0';
		pld_pma_adapt_start	:	in	std_logic	:=	'0';
		pld_pma_csr_test_dis	:	in	std_logic	:=	'0';
		pld_pma_early_eios	:	in	std_logic	:=	'0';
		pld_pma_eye_monitor	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		pld_pma_ltd_b	:	in	std_logic	:=	'0';
		pld_pma_nrpi_freeze	:	in	std_logic	:=	'0';
		pld_pma_pcie_switch	:	in	std_logic_vector(1 downto 0)	:=	"00";
		pld_pma_ppm_lock	:	in	std_logic	:=	'0';
		pld_pma_reserved_out	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		pld_pma_rs_lpbk_b	:	in	std_logic	:=	'0';
		pld_pma_rx_qpi_pullup	:	in	std_logic	:=	'0';
		pld_pma_tx_bitslip	:	in	std_logic	:=	'0';
		pld_pma_tx_bonding_rstb	:	in	std_logic	:=	'0';
		pld_pma_tx_qpi_pulldn	:	in	std_logic	:=	'0';
		pld_pma_tx_qpi_pullup	:	in	std_logic	:=	'0';
		pld_pma_txdetectrx	:	in	std_logic	:=	'0';
		pld_rate	:	in	std_logic_vector(1 downto 0)	:=	"00";
		pld_reserved_in	:	in	std_logic_vector(9 downto 0)	:=	"0000000000";
		pld_scan_mode_n	:	in	std_logic	:=	'0';
		pld_scan_shift_n	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		pld_8g_eidleinfersel_fifo	:	out	std_logic	:=	'0';
		pld_8g_eidleinfersel_reg	:	out	std_logic	:=	'0';
		pld_partial_reconfig_fifo	:	out	std_logic	:=	'0';
		pld_partial_reconfig_rx_div_by_2_rxclk_wire	:	out	std_logic	:=	'0';
		pld_partial_reconfig_rx_div_by_2_txclk_wire	:	out	std_logic	:=	'0';
		pld_partial_reconfig_rxclk_reg	:	out	std_logic	:=	'0';
		pld_partial_reconfig_tx_div_by_2_wire	:	out	std_logic	:=	'0';
		pld_partial_reconfig_txclk_reg	:	out	std_logic	:=	'0';
		pld_rate_reg	:	out	std_logic	:=	'0';
		pld_test_data_reg	:	out	std_logic	:=	'0';
		hip_cmn_clk	:	out	std_logic_vector(1 downto 0)	:=	"00";
		hip_cmn_ctrl	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		hip_iocsr_rdy	:	out	std_logic	:=	'0';
		hip_iocsr_rdy_dly	:	out	std_logic	:=	'0';
		hip_nfrzdrv	:	out	std_logic	:=	'0';
		hip_npor	:	out	std_logic	:=	'0';
		hip_usermode	:	out	std_logic	:=	'0';
		int_pldif_10g_refclk_dig	:	out	std_logic	:=	'0';
		int_pldif_10g_scan_mode_n	:	out	std_logic	:=	'0';
		int_pldif_8g_eidleinfersel	:	out	std_logic_vector(2 downto 0)	:=	"000";
		int_pldif_8g_ltr	:	out	std_logic	:=	'0';
		int_pldif_8g_refclk_dig	:	out	std_logic	:=	'0';
		int_pldif_8g_refclk_dig2	:	out	std_logic	:=	'0';
		int_pldif_8g_scan_mode_n	:	out	std_logic	:=	'0';
		int_pldif_avmm_pld_avmm1_request	:	out	std_logic	:=	'0';
		int_pldif_avmm_pld_avmm2_request	:	out	std_logic	:=	'0';
		int_pldif_g3_current_coeff	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		int_pldif_g3_current_rxpreset	:	out	std_logic_vector(2 downto 0)	:=	"000";
		int_pldif_g3_scan_mode_n	:	out	std_logic	:=	'0';
		int_pldif_krfec_refclk_dig	:	out	std_logic	:=	'0';
		int_pldif_krfec_scan_mode_n	:	out	std_logic	:=	'0';
		int_pldif_krfec_scan_rst_n	:	out	std_logic	:=	'0';
		int_pldif_mem_atpg_rst_n	:	out	std_logic	:=	'0';
		int_pldif_mem_scan_mode_n	:	out	std_logic	:=	'0';
		int_pldif_pmaif_adapt_start	:	out	std_logic	:=	'0';
		int_pldif_pmaif_atpg_los_en_n	:	out	std_logic	:=	'0';
		int_pldif_pmaif_csr_test_dis	:	out	std_logic	:=	'0';
		int_pldif_pmaif_early_eios	:	out	std_logic	:=	'0';
		int_pldif_pmaif_eye_monitor	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		int_pldif_pmaif_ltd_b	:	out	std_logic	:=	'0';
		int_pldif_pmaif_ltr	:	out	std_logic	:=	'0';
		int_pldif_pmaif_nfrzdrv	:	out	std_logic	:=	'0';
		int_pldif_pmaif_nrpi_freeze	:	out	std_logic	:=	'0';
		int_pldif_pmaif_pcie_switch	:	out	std_logic_vector(1 downto 0)	:=	"00";
		int_pldif_pmaif_pma_reserved_out	:	out	std_logic_vector(4 downto 0)	:=	"00000";
		int_pldif_pmaif_pma_scan_mode_n	:	out	std_logic	:=	'0';
		int_pldif_pmaif_pma_scan_shift_n	:	out	std_logic	:=	'0';
		int_pldif_pmaif_ppm_lock	:	out	std_logic	:=	'0';
		int_pldif_pmaif_rate	:	out	std_logic_vector(1 downto 0)	:=	"00";
		int_pldif_pmaif_refclk_dig	:	out	std_logic	:=	'0';
		int_pldif_pmaif_rs_lpbk_b	:	out	std_logic	:=	'0';
		int_pldif_pmaif_rx_qpi_pullup	:	out	std_logic	:=	'0';
		int_pldif_pmaif_scan_mode_n	:	out	std_logic	:=	'0';
		int_pldif_pmaif_tx_bitslip	:	out	std_logic	:=	'0';
		int_pldif_pmaif_tx_bonding_rstb	:	out	std_logic	:=	'0';
		int_pldif_pmaif_tx_pma_syncp_hip	:	out	std_logic	:=	'0';
		int_pldif_pmaif_tx_qpi_pulldn	:	out	std_logic	:=	'0';
		int_pldif_pmaif_tx_qpi_pullup	:	out	std_logic	:=	'0';
		int_pldif_pmaif_txdetectrx	:	out	std_logic	:=	'0';
		int_pldif_pmaif_uhsif_refclk_dig	:	out	std_logic	:=	'0';
		int_pldif_usr_rst_sel	:	out	std_logic	:=	'0';
		int_pmaif_pldif_uhsif_scan_chain_in	:	out	std_logic	:=	'0';
		pld_pma_adapt_done	:	out	std_logic	:=	'0';
		pld_pma_clklow	:	out	std_logic	:=	'0';
		pld_pma_fref	:	out	std_logic	:=	'0';
		pld_pma_hclk	:	out	std_logic	:=	'0';
		pld_pma_pcie_sw_done	:	out	std_logic_vector(1 downto 0)	:=	"00";
		pld_pma_pfdmode_lock	:	out	std_logic	:=	'0';
		pld_pma_reserved_in	:	out	std_logic_vector(4 downto 0)	:=	"00000";
		pld_pma_rx_detect_valid	:	out	std_logic	:=	'0';
		pld_pma_rx_found	:	out	std_logic	:=	'0';
		pld_pma_rxpll_lock	:	out	std_logic	:=	'0';
		pld_pma_testbus	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		pld_pmaif_mask_tx_pll	:	out	std_logic	:=	'0';
		pld_reserved_out	:	out	std_logic_vector(9 downto 0)	:=	"0000000000";
		pld_test_data	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		pld_uhsif_lock	:	out	std_logic	:=	'0';
		scan_mode_n	:	out	std_logic	:=	'0'
	);
end twentynm_hssi_common_pld_pcs_interface;

architecture behavior of twentynm_hssi_common_pld_pcs_interface	is




component	twentynm_hssi_common_pld_pcs_interface_encrypted
	generic (
		-- Architecture parameters
		dft_clk_out_en	:	string	:=	"dft_clk_out_disable";
		dft_clk_out_sel	:	string	:=	"teng_rx_dft_clk";
		hrdrstctrl_en	:	string	:=	"hrst_dis";
		pcs_testbus_block_sel	:	string	:=	"eightg";
		reconfig_settings	:	string	:=	"{}";
		silicon_rev	:	string	:=	"20nm5es"
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		int_pldif_10g_rx_dft_clk_out	:	in	std_logic	:=	'0';
		int_pldif_10g_test_data	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		int_pldif_10g_tx_dft_clk_out	:	in	std_logic	:=	'0';
		int_pldif_8g_chnl_test_bus_out	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		int_pldif_8g_rx_clk_to_observation_ff_in_pld_if	:	in	std_logic	:=	'0';
		int_pldif_8g_tx_clk_to_observation_ff_in_pld_if	:	in	std_logic	:=	'0';
		int_pldif_avmm_refclk_dig_en	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		int_pldif_g3_test_out	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		int_pldif_krfec_test_data	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		int_pldif_pmaif_adapt_done	:	in	std_logic	:=	'0';
		int_pldif_pmaif_mask_tx_pll	:	in	std_logic	:=	'0';
		int_pldif_pmaif_pcie_sw_done	:	in	std_logic_vector(1 downto 0)	:=	"00";
		int_pldif_pmaif_pfdmode_lock	:	in	std_logic	:=	'0';
		int_pldif_pmaif_pma_clklow	:	in	std_logic	:=	'0';
		int_pldif_pmaif_pma_fref	:	in	std_logic	:=	'0';
		int_pldif_pmaif_pma_hclk	:	in	std_logic	:=	'0';
		int_pldif_pmaif_pma_reserved_in	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		int_pldif_pmaif_rx_detect_valid	:	in	std_logic	:=	'0';
		int_pldif_pmaif_rx_found	:	in	std_logic	:=	'0';
		int_pldif_pmaif_rxpll_lock	:	in	std_logic	:=	'0';
		int_pldif_pmaif_test_out	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		int_pldif_pmaif_testbus	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		int_pldif_pmaif_uhsif_lock	:	in	std_logic	:=	'0';
		int_pmaif_pldif_dft_obsrv_clk	:	in	std_logic	:=	'0';
		int_pmaif_pldif_uhsif_scan_chain_out	:	in	std_logic	:=	'0';
		pld_8g_eidleinfersel	:	in	std_logic_vector(2 downto 0)	:=	"000";
		pld_8g_refclk_dig2	:	in	std_logic	:=	'0';
		pld_atpg_los_en_n	:	in	std_logic	:=	'0';
		pld_g3_current_coeff	:	in	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		pld_g3_current_rxpreset	:	in	std_logic_vector(2 downto 0)	:=	"000";
		pld_ltr	:	in	std_logic	:=	'0';
		pld_mem_krfec_atpg_rst_n	:	in	std_logic	:=	'0';
		pld_partial_reconfig	:	in	std_logic	:=	'0';
		pld_pcs_refclk_dig	:	in	std_logic	:=	'0';
		pld_pma_adapt_start	:	in	std_logic	:=	'0';
		pld_pma_csr_test_dis	:	in	std_logic	:=	'0';
		pld_pma_early_eios	:	in	std_logic	:=	'0';
		pld_pma_eye_monitor	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		pld_pma_ltd_b	:	in	std_logic	:=	'0';
		pld_pma_nrpi_freeze	:	in	std_logic	:=	'0';
		pld_pma_pcie_switch	:	in	std_logic_vector(1 downto 0)	:=	"00";
		pld_pma_ppm_lock	:	in	std_logic	:=	'0';
		pld_pma_reserved_out	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		pld_pma_rs_lpbk_b	:	in	std_logic	:=	'0';
		pld_pma_rx_qpi_pullup	:	in	std_logic	:=	'0';
		pld_pma_tx_bitslip	:	in	std_logic	:=	'0';
		pld_pma_tx_bonding_rstb	:	in	std_logic	:=	'0';
		pld_pma_tx_qpi_pulldn	:	in	std_logic	:=	'0';
		pld_pma_tx_qpi_pullup	:	in	std_logic	:=	'0';
		pld_pma_txdetectrx	:	in	std_logic	:=	'0';
		pld_rate	:	in	std_logic_vector(1 downto 0)	:=	"00";
		pld_reserved_in	:	in	std_logic_vector(9 downto 0)	:=	"0000000000";
		pld_scan_mode_n	:	in	std_logic	:=	'0';
		pld_scan_shift_n	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		pld_8g_eidleinfersel_fifo	:	out	std_logic	:=	'0';
		pld_8g_eidleinfersel_reg	:	out	std_logic	:=	'0';
		pld_partial_reconfig_fifo	:	out	std_logic	:=	'0';
		pld_partial_reconfig_rx_div_by_2_rxclk_wire	:	out	std_logic	:=	'0';
		pld_partial_reconfig_rx_div_by_2_txclk_wire	:	out	std_logic	:=	'0';
		pld_partial_reconfig_rxclk_reg	:	out	std_logic	:=	'0';
		pld_partial_reconfig_tx_div_by_2_wire	:	out	std_logic	:=	'0';
		pld_partial_reconfig_txclk_reg	:	out	std_logic	:=	'0';
		pld_rate_reg	:	out	std_logic	:=	'0';
		pld_test_data_reg	:	out	std_logic	:=	'0';
		hip_cmn_clk	:	out	std_logic_vector(1 downto 0)	:=	"00";
		hip_cmn_ctrl	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		hip_iocsr_rdy	:	out	std_logic	:=	'0';
		hip_iocsr_rdy_dly	:	out	std_logic	:=	'0';
		hip_nfrzdrv	:	out	std_logic	:=	'0';
		hip_npor	:	out	std_logic	:=	'0';
		hip_usermode	:	out	std_logic	:=	'0';
		int_pldif_10g_refclk_dig	:	out	std_logic	:=	'0';
		int_pldif_10g_scan_mode_n	:	out	std_logic	:=	'0';
		int_pldif_8g_eidleinfersel	:	out	std_logic_vector(2 downto 0)	:=	"000";
		int_pldif_8g_ltr	:	out	std_logic	:=	'0';
		int_pldif_8g_refclk_dig	:	out	std_logic	:=	'0';
		int_pldif_8g_refclk_dig2	:	out	std_logic	:=	'0';
		int_pldif_8g_scan_mode_n	:	out	std_logic	:=	'0';
		int_pldif_avmm_pld_avmm1_request	:	out	std_logic	:=	'0';
		int_pldif_avmm_pld_avmm2_request	:	out	std_logic	:=	'0';
		int_pldif_g3_current_coeff	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		int_pldif_g3_current_rxpreset	:	out	std_logic_vector(2 downto 0)	:=	"000";
		int_pldif_g3_scan_mode_n	:	out	std_logic	:=	'0';
		int_pldif_krfec_refclk_dig	:	out	std_logic	:=	'0';
		int_pldif_krfec_scan_mode_n	:	out	std_logic	:=	'0';
		int_pldif_krfec_scan_rst_n	:	out	std_logic	:=	'0';
		int_pldif_mem_atpg_rst_n	:	out	std_logic	:=	'0';
		int_pldif_mem_scan_mode_n	:	out	std_logic	:=	'0';
		int_pldif_pmaif_adapt_start	:	out	std_logic	:=	'0';
		int_pldif_pmaif_atpg_los_en_n	:	out	std_logic	:=	'0';
		int_pldif_pmaif_csr_test_dis	:	out	std_logic	:=	'0';
		int_pldif_pmaif_early_eios	:	out	std_logic	:=	'0';
		int_pldif_pmaif_eye_monitor	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		int_pldif_pmaif_ltd_b	:	out	std_logic	:=	'0';
		int_pldif_pmaif_ltr	:	out	std_logic	:=	'0';
		int_pldif_pmaif_nfrzdrv	:	out	std_logic	:=	'0';
		int_pldif_pmaif_nrpi_freeze	:	out	std_logic	:=	'0';
		int_pldif_pmaif_pcie_switch	:	out	std_logic_vector(1 downto 0)	:=	"00";
		int_pldif_pmaif_pma_reserved_out	:	out	std_logic_vector(4 downto 0)	:=	"00000";
		int_pldif_pmaif_pma_scan_mode_n	:	out	std_logic	:=	'0';
		int_pldif_pmaif_pma_scan_shift_n	:	out	std_logic	:=	'0';
		int_pldif_pmaif_ppm_lock	:	out	std_logic	:=	'0';
		int_pldif_pmaif_rate	:	out	std_logic_vector(1 downto 0)	:=	"00";
		int_pldif_pmaif_refclk_dig	:	out	std_logic	:=	'0';
		int_pldif_pmaif_rs_lpbk_b	:	out	std_logic	:=	'0';
		int_pldif_pmaif_rx_qpi_pullup	:	out	std_logic	:=	'0';
		int_pldif_pmaif_scan_mode_n	:	out	std_logic	:=	'0';
		int_pldif_pmaif_tx_bitslip	:	out	std_logic	:=	'0';
		int_pldif_pmaif_tx_bonding_rstb	:	out	std_logic	:=	'0';
		int_pldif_pmaif_tx_pma_syncp_hip	:	out	std_logic	:=	'0';
		int_pldif_pmaif_tx_qpi_pulldn	:	out	std_logic	:=	'0';
		int_pldif_pmaif_tx_qpi_pullup	:	out	std_logic	:=	'0';
		int_pldif_pmaif_txdetectrx	:	out	std_logic	:=	'0';
		int_pldif_pmaif_uhsif_refclk_dig	:	out	std_logic	:=	'0';
		int_pldif_usr_rst_sel	:	out	std_logic	:=	'0';
		int_pmaif_pldif_uhsif_scan_chain_in	:	out	std_logic	:=	'0';
		pld_pma_adapt_done	:	out	std_logic	:=	'0';
		pld_pma_clklow	:	out	std_logic	:=	'0';
		pld_pma_fref	:	out	std_logic	:=	'0';
		pld_pma_hclk	:	out	std_logic	:=	'0';
		pld_pma_pcie_sw_done	:	out	std_logic_vector(1 downto 0)	:=	"00";
		pld_pma_pfdmode_lock	:	out	std_logic	:=	'0';
		pld_pma_reserved_in	:	out	std_logic_vector(4 downto 0)	:=	"00000";
		pld_pma_rx_detect_valid	:	out	std_logic	:=	'0';
		pld_pma_rx_found	:	out	std_logic	:=	'0';
		pld_pma_rxpll_lock	:	out	std_logic	:=	'0';
		pld_pma_testbus	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		pld_pmaif_mask_tx_pll	:	out	std_logic	:=	'0';
		pld_reserved_out	:	out	std_logic_vector(9 downto 0)	:=	"0000000000";
		pld_test_data	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		pld_uhsif_lock	:	out	std_logic	:=	'0';
		scan_mode_n	:	out	std_logic	:=	'0'
	);
end component;

begin



inst : twentynm_hssi_common_pld_pcs_interface_encrypted
	generic map (
		-- Instance parameters
		dft_clk_out_en	=>	dft_clk_out_en,
		dft_clk_out_sel	=>	dft_clk_out_sel,
		hrdrstctrl_en	=>	hrdrstctrl_en,
		pcs_testbus_block_sel	=>	pcs_testbus_block_sel,
		reconfig_settings	=>	reconfig_settings,
		silicon_rev	=>	silicon_rev
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		int_pldif_10g_rx_dft_clk_out	=>	int_pldif_10g_rx_dft_clk_out,
		int_pldif_10g_test_data	=>	int_pldif_10g_test_data,
		int_pldif_10g_tx_dft_clk_out	=>	int_pldif_10g_tx_dft_clk_out,
		int_pldif_8g_chnl_test_bus_out	=>	int_pldif_8g_chnl_test_bus_out,
		int_pldif_8g_rx_clk_to_observation_ff_in_pld_if	=>	int_pldif_8g_rx_clk_to_observation_ff_in_pld_if,
		int_pldif_8g_tx_clk_to_observation_ff_in_pld_if	=>	int_pldif_8g_tx_clk_to_observation_ff_in_pld_if,
		int_pldif_avmm_refclk_dig_en	=>	int_pldif_avmm_refclk_dig_en,
		int_pldif_g3_test_out	=>	int_pldif_g3_test_out,
		int_pldif_krfec_test_data	=>	int_pldif_krfec_test_data,
		int_pldif_pmaif_adapt_done	=>	int_pldif_pmaif_adapt_done,
		int_pldif_pmaif_mask_tx_pll	=>	int_pldif_pmaif_mask_tx_pll,
		int_pldif_pmaif_pcie_sw_done	=>	int_pldif_pmaif_pcie_sw_done,
		int_pldif_pmaif_pfdmode_lock	=>	int_pldif_pmaif_pfdmode_lock,
		int_pldif_pmaif_pma_clklow	=>	int_pldif_pmaif_pma_clklow,
		int_pldif_pmaif_pma_fref	=>	int_pldif_pmaif_pma_fref,
		int_pldif_pmaif_pma_hclk	=>	int_pldif_pmaif_pma_hclk,
		int_pldif_pmaif_pma_reserved_in	=>	int_pldif_pmaif_pma_reserved_in,
		int_pldif_pmaif_rx_detect_valid	=>	int_pldif_pmaif_rx_detect_valid,
		int_pldif_pmaif_rx_found	=>	int_pldif_pmaif_rx_found,
		int_pldif_pmaif_rxpll_lock	=>	int_pldif_pmaif_rxpll_lock,
		int_pldif_pmaif_test_out	=>	int_pldif_pmaif_test_out,
		int_pldif_pmaif_testbus	=>	int_pldif_pmaif_testbus,
		int_pldif_pmaif_uhsif_lock	=>	int_pldif_pmaif_uhsif_lock,
		int_pmaif_pldif_dft_obsrv_clk	=>	int_pmaif_pldif_dft_obsrv_clk,
		int_pmaif_pldif_uhsif_scan_chain_out	=>	int_pmaif_pldif_uhsif_scan_chain_out,
		pld_8g_eidleinfersel	=>	pld_8g_eidleinfersel,
		pld_8g_refclk_dig2	=>	pld_8g_refclk_dig2,
		pld_atpg_los_en_n	=>	pld_atpg_los_en_n,
		pld_g3_current_coeff	=>	pld_g3_current_coeff,
		pld_g3_current_rxpreset	=>	pld_g3_current_rxpreset,
		pld_ltr	=>	pld_ltr,
		pld_mem_krfec_atpg_rst_n	=>	pld_mem_krfec_atpg_rst_n,
		pld_partial_reconfig	=>	pld_partial_reconfig,
		pld_pcs_refclk_dig	=>	pld_pcs_refclk_dig,
		pld_pma_adapt_start	=>	pld_pma_adapt_start,
		pld_pma_csr_test_dis	=>	pld_pma_csr_test_dis,
		pld_pma_early_eios	=>	pld_pma_early_eios,
		pld_pma_eye_monitor	=>	pld_pma_eye_monitor,
		pld_pma_ltd_b	=>	pld_pma_ltd_b,
		pld_pma_nrpi_freeze	=>	pld_pma_nrpi_freeze,
		pld_pma_pcie_switch	=>	pld_pma_pcie_switch,
		pld_pma_ppm_lock	=>	pld_pma_ppm_lock,
		pld_pma_reserved_out	=>	pld_pma_reserved_out,
		pld_pma_rs_lpbk_b	=>	pld_pma_rs_lpbk_b,
		pld_pma_rx_qpi_pullup	=>	pld_pma_rx_qpi_pullup,
		pld_pma_tx_bitslip	=>	pld_pma_tx_bitslip,
		pld_pma_tx_bonding_rstb	=>	pld_pma_tx_bonding_rstb,
		pld_pma_tx_qpi_pulldn	=>	pld_pma_tx_qpi_pulldn,
		pld_pma_tx_qpi_pullup	=>	pld_pma_tx_qpi_pullup,
		pld_pma_txdetectrx	=>	pld_pma_txdetectrx,
		pld_rate	=>	pld_rate,
		pld_reserved_in	=>	pld_reserved_in,
		pld_scan_mode_n	=>	pld_scan_mode_n,
		pld_scan_shift_n	=>	pld_scan_shift_n,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		pld_8g_eidleinfersel_fifo	=>	pld_8g_eidleinfersel_fifo,
		pld_8g_eidleinfersel_reg	=>	pld_8g_eidleinfersel_reg,
		pld_partial_reconfig_fifo	=>	pld_partial_reconfig_fifo,
		pld_partial_reconfig_rx_div_by_2_rxclk_wire	=>	pld_partial_reconfig_rx_div_by_2_rxclk_wire,
		pld_partial_reconfig_rx_div_by_2_txclk_wire	=>	pld_partial_reconfig_rx_div_by_2_txclk_wire,
		pld_partial_reconfig_rxclk_reg	=>	pld_partial_reconfig_rxclk_reg,
		pld_partial_reconfig_tx_div_by_2_wire	=>	pld_partial_reconfig_tx_div_by_2_wire,
		pld_partial_reconfig_txclk_reg	=>	pld_partial_reconfig_txclk_reg,
		pld_rate_reg	=>	pld_rate_reg,
		pld_test_data_reg	=>	pld_test_data_reg,
		hip_cmn_clk	=>	hip_cmn_clk,
		hip_cmn_ctrl	=>	hip_cmn_ctrl,
		hip_iocsr_rdy	=>	hip_iocsr_rdy,
		hip_iocsr_rdy_dly	=>	hip_iocsr_rdy_dly,
		hip_nfrzdrv	=>	hip_nfrzdrv,
		hip_npor	=>	hip_npor,
		hip_usermode	=>	hip_usermode,
		int_pldif_10g_refclk_dig	=>	int_pldif_10g_refclk_dig,
		int_pldif_10g_scan_mode_n	=>	int_pldif_10g_scan_mode_n,
		int_pldif_8g_eidleinfersel	=>	int_pldif_8g_eidleinfersel,
		int_pldif_8g_ltr	=>	int_pldif_8g_ltr,
		int_pldif_8g_refclk_dig	=>	int_pldif_8g_refclk_dig,
		int_pldif_8g_refclk_dig2	=>	int_pldif_8g_refclk_dig2,
		int_pldif_8g_scan_mode_n	=>	int_pldif_8g_scan_mode_n,
		int_pldif_avmm_pld_avmm1_request	=>	int_pldif_avmm_pld_avmm1_request,
		int_pldif_avmm_pld_avmm2_request	=>	int_pldif_avmm_pld_avmm2_request,
		int_pldif_g3_current_coeff	=>	int_pldif_g3_current_coeff,
		int_pldif_g3_current_rxpreset	=>	int_pldif_g3_current_rxpreset,
		int_pldif_g3_scan_mode_n	=>	int_pldif_g3_scan_mode_n,
		int_pldif_krfec_refclk_dig	=>	int_pldif_krfec_refclk_dig,
		int_pldif_krfec_scan_mode_n	=>	int_pldif_krfec_scan_mode_n,
		int_pldif_krfec_scan_rst_n	=>	int_pldif_krfec_scan_rst_n,
		int_pldif_mem_atpg_rst_n	=>	int_pldif_mem_atpg_rst_n,
		int_pldif_mem_scan_mode_n	=>	int_pldif_mem_scan_mode_n,
		int_pldif_pmaif_adapt_start	=>	int_pldif_pmaif_adapt_start,
		int_pldif_pmaif_atpg_los_en_n	=>	int_pldif_pmaif_atpg_los_en_n,
		int_pldif_pmaif_csr_test_dis	=>	int_pldif_pmaif_csr_test_dis,
		int_pldif_pmaif_early_eios	=>	int_pldif_pmaif_early_eios,
		int_pldif_pmaif_eye_monitor	=>	int_pldif_pmaif_eye_monitor,
		int_pldif_pmaif_ltd_b	=>	int_pldif_pmaif_ltd_b,
		int_pldif_pmaif_ltr	=>	int_pldif_pmaif_ltr,
		int_pldif_pmaif_nfrzdrv	=>	int_pldif_pmaif_nfrzdrv,
		int_pldif_pmaif_nrpi_freeze	=>	int_pldif_pmaif_nrpi_freeze,
		int_pldif_pmaif_pcie_switch	=>	int_pldif_pmaif_pcie_switch,
		int_pldif_pmaif_pma_reserved_out	=>	int_pldif_pmaif_pma_reserved_out,
		int_pldif_pmaif_pma_scan_mode_n	=>	int_pldif_pmaif_pma_scan_mode_n,
		int_pldif_pmaif_pma_scan_shift_n	=>	int_pldif_pmaif_pma_scan_shift_n,
		int_pldif_pmaif_ppm_lock	=>	int_pldif_pmaif_ppm_lock,
		int_pldif_pmaif_rate	=>	int_pldif_pmaif_rate,
		int_pldif_pmaif_refclk_dig	=>	int_pldif_pmaif_refclk_dig,
		int_pldif_pmaif_rs_lpbk_b	=>	int_pldif_pmaif_rs_lpbk_b,
		int_pldif_pmaif_rx_qpi_pullup	=>	int_pldif_pmaif_rx_qpi_pullup,
		int_pldif_pmaif_scan_mode_n	=>	int_pldif_pmaif_scan_mode_n,
		int_pldif_pmaif_tx_bitslip	=>	int_pldif_pmaif_tx_bitslip,
		int_pldif_pmaif_tx_bonding_rstb	=>	int_pldif_pmaif_tx_bonding_rstb,
		int_pldif_pmaif_tx_pma_syncp_hip	=>	int_pldif_pmaif_tx_pma_syncp_hip,
		int_pldif_pmaif_tx_qpi_pulldn	=>	int_pldif_pmaif_tx_qpi_pulldn,
		int_pldif_pmaif_tx_qpi_pullup	=>	int_pldif_pmaif_tx_qpi_pullup,
		int_pldif_pmaif_txdetectrx	=>	int_pldif_pmaif_txdetectrx,
		int_pldif_pmaif_uhsif_refclk_dig	=>	int_pldif_pmaif_uhsif_refclk_dig,
		int_pldif_usr_rst_sel	=>	int_pldif_usr_rst_sel,
		int_pmaif_pldif_uhsif_scan_chain_in	=>	int_pmaif_pldif_uhsif_scan_chain_in,
		pld_pma_adapt_done	=>	pld_pma_adapt_done,
		pld_pma_clklow	=>	pld_pma_clklow,
		pld_pma_fref	=>	pld_pma_fref,
		pld_pma_hclk	=>	pld_pma_hclk,
		pld_pma_pcie_sw_done	=>	pld_pma_pcie_sw_done,
		pld_pma_pfdmode_lock	=>	pld_pma_pfdmode_lock,
		pld_pma_reserved_in	=>	pld_pma_reserved_in,
		pld_pma_rx_detect_valid	=>	pld_pma_rx_detect_valid,
		pld_pma_rx_found	=>	pld_pma_rx_found,
		pld_pma_rxpll_lock	=>	pld_pma_rxpll_lock,
		pld_pma_testbus	=>	pld_pma_testbus,
		pld_pmaif_mask_tx_pll	=>	pld_pmaif_mask_tx_pll,
		pld_reserved_out	=>	pld_reserved_out,
		pld_test_data	=>	pld_test_data,
		pld_uhsif_lock	=>	pld_uhsif_lock,
		scan_mode_n	=>	scan_mode_n
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_fifo_rx_pcs	is
	generic (
		-- Entity parameters
		double_read_mode	:	string	:=	"double_read_dis";
		prot_mode	:	string	:=	"teng_mode";
		silicon_rev	:	string	:=	"20nm5es"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		atpg_rst_n	:	in	std_logic	:=	'0';
		data_in_10g	:	in	std_logic_vector(73 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000";
		data_in_8g_clock_comp	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		data_in_8g_phase_comp	:	in	std_logic_vector(79 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
		data_in_gen3	:	in	std_logic_vector(39 downto 0)	:=	"0000000000000000000000000000000000000000";
		hard_reset_n	:	in	std_logic	:=	'0';
		rd_ptr2_10g	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rd_ptr2_8g_clock_comp	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		rd_ptr_10g	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rd_ptr_8g_clock_comp	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		rd_ptr_8g_phase_comp	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		rd_ptr_gen3	:	in	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		scan_mode_n	:	in	std_logic	:=	'0';
		wr_clk_10g	:	in	std_logic	:=	'0';
		wr_clk_8g_clock_comp_dw	:	in	std_logic	:=	'0';
		wr_clk_8g_clock_comp_sw	:	in	std_logic	:=	'0';
		wr_clk_8g_phase_comp_dw	:	in	std_logic	:=	'0';
		wr_clk_8g_phase_comp_sw	:	in	std_logic	:=	'0';
		wr_clk_gen3	:	in	std_logic	:=	'0';
		wr_en_10g	:	in	std_logic	:=	'0';
		wr_en_8g_clock_comp	:	in	std_logic	:=	'0';
		wr_en_8g_phase_comp	:	in	std_logic	:=	'0';
		wr_en_gen3	:	in	std_logic	:=	'0';
		wr_ptr_10g	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		wr_ptr_8g_clock_comp	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		wr_ptr_8g_phase_comp	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		wr_ptr_gen3	:	in	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		wr_rst_n_10g	:	in	std_logic	:=	'0';
		wr_rst_n_8g_clock_comp	:	in	std_logic	:=	'0';
		wr_rst_n_8g_phase_comp	:	in	std_logic	:=	'0';
		wr_rst_n_gen3	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		data_out2_10g	:	out	std_logic_vector(73 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000";
		data_out2_8g_clock_comp	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		data_out_10g	:	out	std_logic_vector(73 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000";
		data_out_8g_clock_comp	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		data_out_8g_phase_comp	:	out	std_logic_vector(79 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
		data_out_gen3	:	out	std_logic_vector(39 downto 0)	:=	"0000000000000000000000000000000000000000"
	);
end twentynm_hssi_fifo_rx_pcs;

architecture behavior of twentynm_hssi_fifo_rx_pcs	is




component	twentynm_hssi_fifo_rx_pcs_encrypted
	generic (
		-- Architecture parameters
		double_read_mode	:	string	:=	"double_read_dis";
		prot_mode	:	string	:=	"teng_mode";
		silicon_rev	:	string	:=	"20nm5es"
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		atpg_rst_n	:	in	std_logic	:=	'0';
		data_in_10g	:	in	std_logic_vector(73 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000";
		data_in_8g_clock_comp	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		data_in_8g_phase_comp	:	in	std_logic_vector(79 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
		data_in_gen3	:	in	std_logic_vector(39 downto 0)	:=	"0000000000000000000000000000000000000000";
		hard_reset_n	:	in	std_logic	:=	'0';
		rd_ptr2_10g	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rd_ptr2_8g_clock_comp	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		rd_ptr_10g	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rd_ptr_8g_clock_comp	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		rd_ptr_8g_phase_comp	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		rd_ptr_gen3	:	in	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		scan_mode_n	:	in	std_logic	:=	'0';
		wr_clk_10g	:	in	std_logic	:=	'0';
		wr_clk_8g_clock_comp_dw	:	in	std_logic	:=	'0';
		wr_clk_8g_clock_comp_sw	:	in	std_logic	:=	'0';
		wr_clk_8g_phase_comp_dw	:	in	std_logic	:=	'0';
		wr_clk_8g_phase_comp_sw	:	in	std_logic	:=	'0';
		wr_clk_gen3	:	in	std_logic	:=	'0';
		wr_en_10g	:	in	std_logic	:=	'0';
		wr_en_8g_clock_comp	:	in	std_logic	:=	'0';
		wr_en_8g_phase_comp	:	in	std_logic	:=	'0';
		wr_en_gen3	:	in	std_logic	:=	'0';
		wr_ptr_10g	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		wr_ptr_8g_clock_comp	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		wr_ptr_8g_phase_comp	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		wr_ptr_gen3	:	in	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		wr_rst_n_10g	:	in	std_logic	:=	'0';
		wr_rst_n_8g_clock_comp	:	in	std_logic	:=	'0';
		wr_rst_n_8g_phase_comp	:	in	std_logic	:=	'0';
		wr_rst_n_gen3	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		data_out2_10g	:	out	std_logic_vector(73 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000";
		data_out2_8g_clock_comp	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		data_out_10g	:	out	std_logic_vector(73 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000";
		data_out_8g_clock_comp	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		data_out_8g_phase_comp	:	out	std_logic_vector(79 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000000000";
		data_out_gen3	:	out	std_logic_vector(39 downto 0)	:=	"0000000000000000000000000000000000000000"
	);
end component;

begin



inst : twentynm_hssi_fifo_rx_pcs_encrypted
	generic map (
		-- Instance parameters
		double_read_mode	=>	double_read_mode,
		prot_mode	=>	prot_mode,
		silicon_rev	=>	silicon_rev
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		atpg_rst_n	=>	atpg_rst_n,
		data_in_10g	=>	data_in_10g,
		data_in_8g_clock_comp	=>	data_in_8g_clock_comp,
		data_in_8g_phase_comp	=>	data_in_8g_phase_comp,
		data_in_gen3	=>	data_in_gen3,
		hard_reset_n	=>	hard_reset_n,
		rd_ptr2_10g	=>	rd_ptr2_10g,
		rd_ptr2_8g_clock_comp	=>	rd_ptr2_8g_clock_comp,
		rd_ptr_10g	=>	rd_ptr_10g,
		rd_ptr_8g_clock_comp	=>	rd_ptr_8g_clock_comp,
		rd_ptr_8g_phase_comp	=>	rd_ptr_8g_phase_comp,
		rd_ptr_gen3	=>	rd_ptr_gen3,
		scan_mode_n	=>	scan_mode_n,
		wr_clk_10g	=>	wr_clk_10g,
		wr_clk_8g_clock_comp_dw	=>	wr_clk_8g_clock_comp_dw,
		wr_clk_8g_clock_comp_sw	=>	wr_clk_8g_clock_comp_sw,
		wr_clk_8g_phase_comp_dw	=>	wr_clk_8g_phase_comp_dw,
		wr_clk_8g_phase_comp_sw	=>	wr_clk_8g_phase_comp_sw,
		wr_clk_gen3	=>	wr_clk_gen3,
		wr_en_10g	=>	wr_en_10g,
		wr_en_8g_clock_comp	=>	wr_en_8g_clock_comp,
		wr_en_8g_phase_comp	=>	wr_en_8g_phase_comp,
		wr_en_gen3	=>	wr_en_gen3,
		wr_ptr_10g	=>	wr_ptr_10g,
		wr_ptr_8g_clock_comp	=>	wr_ptr_8g_clock_comp,
		wr_ptr_8g_phase_comp	=>	wr_ptr_8g_phase_comp,
		wr_ptr_gen3	=>	wr_ptr_gen3,
		wr_rst_n_10g	=>	wr_rst_n_10g,
		wr_rst_n_8g_clock_comp	=>	wr_rst_n_8g_clock_comp,
		wr_rst_n_8g_phase_comp	=>	wr_rst_n_8g_phase_comp,
		wr_rst_n_gen3	=>	wr_rst_n_gen3,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		data_out2_10g	=>	data_out2_10g,
		data_out2_8g_clock_comp	=>	data_out2_8g_clock_comp,
		data_out_10g	=>	data_out_10g,
		data_out_8g_clock_comp	=>	data_out_8g_clock_comp,
		data_out_8g_phase_comp	=>	data_out_8g_phase_comp,
		data_out_gen3	=>	data_out_gen3
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_fifo_tx_pcs	is
	generic (
		-- Entity parameters
		double_write_mode	:	string	:=	"double_write_dis";
		prot_mode	:	string	:=	"teng_mode";
		silicon_rev	:	string	:=	"20nm5es"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		atpg_rst_n	:	in	std_logic	:=	'0';
		data_in2_10g	:	in	std_logic_vector(72 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000000000000";
		data_in_10g	:	in	std_logic_vector(72 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000000000000";
		data_in_8g_phase_comp	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		hard_reset_n	:	in	std_logic	:=	'0';
		rd_ptr_10g	:	in	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		rd_ptr_8g_phase_comp	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		scan_mode_n	:	in	std_logic	:=	'0';
		wr_clk_10g	:	in	std_logic	:=	'0';
		wr_clk_8g_phase_comp_dw	:	in	std_logic	:=	'0';
		wr_clk_8g_phase_comp_sw	:	in	std_logic	:=	'0';
		wr_en_10g	:	in	std_logic	:=	'0';
		wr_en_8g_phase_comp	:	in	std_logic	:=	'0';
		wr_ptr_10g	:	in	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		wr_ptr_8g_phase_comp	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		wr_rst_n_10g	:	in	std_logic	:=	'0';
		wr_rst_n_8g_phase_comp	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		data_out_10g	:	out	std_logic_vector(72 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000000000000";
		data_out_8g_phase_comp	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000"
	);
end twentynm_hssi_fifo_tx_pcs;

architecture behavior of twentynm_hssi_fifo_tx_pcs	is




component	twentynm_hssi_fifo_tx_pcs_encrypted
	generic (
		-- Architecture parameters
		double_write_mode	:	string	:=	"double_write_dis";
		prot_mode	:	string	:=	"teng_mode";
		silicon_rev	:	string	:=	"20nm5es"
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		atpg_rst_n	:	in	std_logic	:=	'0';
		data_in2_10g	:	in	std_logic_vector(72 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000000000000";
		data_in_10g	:	in	std_logic_vector(72 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000000000000";
		data_in_8g_phase_comp	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		hard_reset_n	:	in	std_logic	:=	'0';
		rd_ptr_10g	:	in	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		rd_ptr_8g_phase_comp	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		scan_mode_n	:	in	std_logic	:=	'0';
		wr_clk_10g	:	in	std_logic	:=	'0';
		wr_clk_8g_phase_comp_dw	:	in	std_logic	:=	'0';
		wr_clk_8g_phase_comp_sw	:	in	std_logic	:=	'0';
		wr_en_10g	:	in	std_logic	:=	'0';
		wr_en_8g_phase_comp	:	in	std_logic	:=	'0';
		wr_ptr_10g	:	in	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		wr_ptr_8g_phase_comp	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		wr_rst_n_10g	:	in	std_logic	:=	'0';
		wr_rst_n_8g_phase_comp	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		data_out_10g	:	out	std_logic_vector(72 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000000000000";
		data_out_8g_phase_comp	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000"
	);
end component;

begin



inst : twentynm_hssi_fifo_tx_pcs_encrypted
	generic map (
		-- Instance parameters
		double_write_mode	=>	double_write_mode,
		prot_mode	=>	prot_mode,
		silicon_rev	=>	silicon_rev
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		atpg_rst_n	=>	atpg_rst_n,
		data_in2_10g	=>	data_in2_10g,
		data_in_10g	=>	data_in_10g,
		data_in_8g_phase_comp	=>	data_in_8g_phase_comp,
		hard_reset_n	=>	hard_reset_n,
		rd_ptr_10g	=>	rd_ptr_10g,
		rd_ptr_8g_phase_comp	=>	rd_ptr_8g_phase_comp,
		scan_mode_n	=>	scan_mode_n,
		wr_clk_10g	=>	wr_clk_10g,
		wr_clk_8g_phase_comp_dw	=>	wr_clk_8g_phase_comp_dw,
		wr_clk_8g_phase_comp_sw	=>	wr_clk_8g_phase_comp_sw,
		wr_en_10g	=>	wr_en_10g,
		wr_en_8g_phase_comp	=>	wr_en_8g_phase_comp,
		wr_ptr_10g	=>	wr_ptr_10g,
		wr_ptr_8g_phase_comp	=>	wr_ptr_8g_phase_comp,
		wr_rst_n_10g	=>	wr_rst_n_10g,
		wr_rst_n_8g_phase_comp	=>	wr_rst_n_8g_phase_comp,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		data_out_10g	=>	data_out_10g,
		data_out_8g_phase_comp	=>	data_out_8g_phase_comp
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_gen3_rx_pcs	is
	generic (
		-- Entity parameters
		block_sync	:	string	:=	"enable_block_sync";
		block_sync_sm	:	string	:=	"enable_blk_sync_sm";
		cdr_ctrl_force_unalgn	:	string	:=	"enable";
		lpbk_force	:	string	:=	"lpbk_frce_dis";
		mode	:	string	:=	"gen3_func";
		rate_match_fifo	:	string	:=	"enable_rm_fifo_600ppm";
		rate_match_fifo_latency	:	string	:=	"regular_latency";
		reconfig_settings	:	string	:=	"{}";
		reverse_lpbk	:	string	:=	"rev_lpbk_en";
		rx_b4gb_par_lpbk	:	string	:=	"b4gb_par_lpbk_dis";
		rx_force_balign	:	string	:=	"en_force_balign";
		rx_ins_del_one_skip	:	string	:=	"ins_del_one_skip_en";
		rx_num_fixed_pat	:	bit_vector	:=	B"1000";
		rx_test_out_sel	:	string	:=	"rx_test_out0";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		data_in	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		gen3_clk_sel	:	in	std_logic	:=	'0';
		inferred_rxvalid	:	in	std_logic	:=	'0';
		lpbk_en	:	in	std_logic	:=	'0';
		mem_rx_fifo_rd_data	:	in	std_logic_vector(39 downto 0)	:=	"0000000000000000000000000000000000000000";
		par_lpbk_b4gb_in	:	in	std_logic_vector(35 downto 0)	:=	"000000000000000000000000000000000000";
		par_lpbk_in	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		pcs_rst	:	in	std_logic	:=	'0';
		rcvd_clk	:	in	std_logic	:=	'0';
		rx_pma_clk	:	in	std_logic	:=	'0';
		rx_pma_rstn	:	in	std_logic	:=	'0';
		rx_rcvd_rstn	:	in	std_logic	:=	'0';
		rxpolarity	:	in	std_logic	:=	'0';
		shutdown_clk	:	in	std_logic	:=	'0';
		sync_sm_en	:	in	std_logic	:=	'0';
		txdatak_in	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		blk_algnd_int	:	out	std_logic	:=	'0';
		blk_lockd_int	:	out	std_logic	:=	'0';
		blk_start	:	out	std_logic	:=	'0';
		clkcomp_delete_int	:	out	std_logic	:=	'0';
		clkcomp_insert_int	:	out	std_logic	:=	'0';
		clkcomp_overfl_int	:	out	std_logic	:=	'0';
		clkcomp_undfl_int	:	out	std_logic	:=	'0';
		data_out	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		data_valid	:	out	std_logic	:=	'0';
		ei_det_int	:	out	std_logic	:=	'0';
		ei_partial_det_int	:	out	std_logic	:=	'0';
		err_decode_int	:	out	std_logic	:=	'0';
		i_det_int	:	out	std_logic	:=	'0';
		lpbk_blk_start	:	out	std_logic	:=	'0';
		lpbk_data	:	out	std_logic_vector(33 downto 0)	:=	"0000000000000000000000000000000000";
		lpbk_data_valid	:	out	std_logic	:=	'0';
		mem_rx_fifo_rd_ptr	:	out	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		mem_rx_fifo_wr_clk	:	out	std_logic	:=	'0';
		mem_rx_fifo_wr_data	:	out	std_logic_vector(39 downto 0)	:=	"0000000000000000000000000000000000000000";
		mem_rx_fifo_wr_en	:	out	std_logic	:=	'0';
		mem_rx_fifo_wr_ptr	:	out	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		mem_rx_fifo_wr_rst_n	:	out	std_logic	:=	'0';
		rcv_lfsr_chk_int	:	out	std_logic	:=	'0';
		rx_test_out	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		skp_det_int	:	out	std_logic	:=	'0';
		sync_hdr	:	out	std_logic_vector(1 downto 0)	:=	"00"
	);
end twentynm_hssi_gen3_rx_pcs;

architecture behavior of twentynm_hssi_gen3_rx_pcs	is

constant rx_num_fixed_pat_int	:	integer	:=	bin2int(rx_num_fixed_pat);



component	twentynm_hssi_gen3_rx_pcs_encrypted
	generic (
		-- Architecture parameters
		block_sync	:	string	:=	"enable_block_sync";
		block_sync_sm	:	string	:=	"enable_blk_sync_sm";
		cdr_ctrl_force_unalgn	:	string	:=	"enable";
		lpbk_force	:	string	:=	"lpbk_frce_dis";
		mode	:	string	:=	"gen3_func";
		rate_match_fifo	:	string	:=	"enable_rm_fifo_600ppm";
		rate_match_fifo_latency	:	string	:=	"regular_latency";
		reconfig_settings	:	string	:=	"{}";
		reverse_lpbk	:	string	:=	"rev_lpbk_en";
		rx_b4gb_par_lpbk	:	string	:=	"b4gb_par_lpbk_dis";
		rx_force_balign	:	string	:=	"en_force_balign";
		rx_ins_del_one_skip	:	string	:=	"ins_del_one_skip_en";
		rx_num_fixed_pat	:	integer	:=	8;
		rx_test_out_sel	:	string	:=	"rx_test_out0";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode"
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		data_in	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		gen3_clk_sel	:	in	std_logic	:=	'0';
		inferred_rxvalid	:	in	std_logic	:=	'0';
		lpbk_en	:	in	std_logic	:=	'0';
		mem_rx_fifo_rd_data	:	in	std_logic_vector(39 downto 0)	:=	"0000000000000000000000000000000000000000";
		par_lpbk_b4gb_in	:	in	std_logic_vector(35 downto 0)	:=	"000000000000000000000000000000000000";
		par_lpbk_in	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		pcs_rst	:	in	std_logic	:=	'0';
		rcvd_clk	:	in	std_logic	:=	'0';
		rx_pma_clk	:	in	std_logic	:=	'0';
		rx_pma_rstn	:	in	std_logic	:=	'0';
		rx_rcvd_rstn	:	in	std_logic	:=	'0';
		rxpolarity	:	in	std_logic	:=	'0';
		shutdown_clk	:	in	std_logic	:=	'0';
		sync_sm_en	:	in	std_logic	:=	'0';
		txdatak_in	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		blk_algnd_int	:	out	std_logic	:=	'0';
		blk_lockd_int	:	out	std_logic	:=	'0';
		blk_start	:	out	std_logic	:=	'0';
		clkcomp_delete_int	:	out	std_logic	:=	'0';
		clkcomp_insert_int	:	out	std_logic	:=	'0';
		clkcomp_overfl_int	:	out	std_logic	:=	'0';
		clkcomp_undfl_int	:	out	std_logic	:=	'0';
		data_out	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		data_valid	:	out	std_logic	:=	'0';
		ei_det_int	:	out	std_logic	:=	'0';
		ei_partial_det_int	:	out	std_logic	:=	'0';
		err_decode_int	:	out	std_logic	:=	'0';
		i_det_int	:	out	std_logic	:=	'0';
		lpbk_blk_start	:	out	std_logic	:=	'0';
		lpbk_data	:	out	std_logic_vector(33 downto 0)	:=	"0000000000000000000000000000000000";
		lpbk_data_valid	:	out	std_logic	:=	'0';
		mem_rx_fifo_rd_ptr	:	out	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		mem_rx_fifo_wr_clk	:	out	std_logic	:=	'0';
		mem_rx_fifo_wr_data	:	out	std_logic_vector(39 downto 0)	:=	"0000000000000000000000000000000000000000";
		mem_rx_fifo_wr_en	:	out	std_logic	:=	'0';
		mem_rx_fifo_wr_ptr	:	out	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		mem_rx_fifo_wr_rst_n	:	out	std_logic	:=	'0';
		rcv_lfsr_chk_int	:	out	std_logic	:=	'0';
		rx_test_out	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		skp_det_int	:	out	std_logic	:=	'0';
		sync_hdr	:	out	std_logic_vector(1 downto 0)	:=	"00"
	);
end component;

begin



inst : twentynm_hssi_gen3_rx_pcs_encrypted
	generic map (
		-- Instance parameters
		block_sync	=>	block_sync,
		block_sync_sm	=>	block_sync_sm,
		cdr_ctrl_force_unalgn	=>	cdr_ctrl_force_unalgn,
		lpbk_force	=>	lpbk_force,
		mode	=>	mode,
		rate_match_fifo	=>	rate_match_fifo,
		rate_match_fifo_latency	=>	rate_match_fifo_latency,
		reconfig_settings	=>	reconfig_settings,
		reverse_lpbk	=>	reverse_lpbk,
		rx_b4gb_par_lpbk	=>	rx_b4gb_par_lpbk,
		rx_force_balign	=>	rx_force_balign,
		rx_ins_del_one_skip	=>	rx_ins_del_one_skip,
		rx_num_fixed_pat	=>	rx_num_fixed_pat_int,
		rx_test_out_sel	=>	rx_test_out_sel,
		silicon_rev	=>	silicon_rev,
		sup_mode	=>	sup_mode
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		data_in	=>	data_in,
		gen3_clk_sel	=>	gen3_clk_sel,
		inferred_rxvalid	=>	inferred_rxvalid,
		lpbk_en	=>	lpbk_en,
		mem_rx_fifo_rd_data	=>	mem_rx_fifo_rd_data,
		par_lpbk_b4gb_in	=>	par_lpbk_b4gb_in,
		par_lpbk_in	=>	par_lpbk_in,
		pcs_rst	=>	pcs_rst,
		rcvd_clk	=>	rcvd_clk,
		rx_pma_clk	=>	rx_pma_clk,
		rx_pma_rstn	=>	rx_pma_rstn,
		rx_rcvd_rstn	=>	rx_rcvd_rstn,
		rxpolarity	=>	rxpolarity,
		shutdown_clk	=>	shutdown_clk,
		sync_sm_en	=>	sync_sm_en,
		txdatak_in	=>	txdatak_in,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		blk_algnd_int	=>	blk_algnd_int,
		blk_lockd_int	=>	blk_lockd_int,
		blk_start	=>	blk_start,
		clkcomp_delete_int	=>	clkcomp_delete_int,
		clkcomp_insert_int	=>	clkcomp_insert_int,
		clkcomp_overfl_int	=>	clkcomp_overfl_int,
		clkcomp_undfl_int	=>	clkcomp_undfl_int,
		data_out	=>	data_out,
		data_valid	=>	data_valid,
		ei_det_int	=>	ei_det_int,
		ei_partial_det_int	=>	ei_partial_det_int,
		err_decode_int	=>	err_decode_int,
		i_det_int	=>	i_det_int,
		lpbk_blk_start	=>	lpbk_blk_start,
		lpbk_data	=>	lpbk_data,
		lpbk_data_valid	=>	lpbk_data_valid,
		mem_rx_fifo_rd_ptr	=>	mem_rx_fifo_rd_ptr,
		mem_rx_fifo_wr_clk	=>	mem_rx_fifo_wr_clk,
		mem_rx_fifo_wr_data	=>	mem_rx_fifo_wr_data,
		mem_rx_fifo_wr_en	=>	mem_rx_fifo_wr_en,
		mem_rx_fifo_wr_ptr	=>	mem_rx_fifo_wr_ptr,
		mem_rx_fifo_wr_rst_n	=>	mem_rx_fifo_wr_rst_n,
		rcv_lfsr_chk_int	=>	rcv_lfsr_chk_int,
		rx_test_out	=>	rx_test_out,
		skp_det_int	=>	skp_det_int,
		sync_hdr	=>	sync_hdr
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_gen3_tx_pcs	is
	generic (
		-- Entity parameters
		mode	:	string	:=	"gen3_func";
		reverse_lpbk	:	string	:=	"rev_lpbk_en";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode";
		tx_bitslip	:	bit_vector	:=	B"00000";
		tx_gbox_byp	:	string	:=	"bypass_gbox"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		blk_start_in	:	in	std_logic	:=	'0';
		data_in	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		data_valid	:	in	std_logic	:=	'0';
		lpbk_blk_start	:	in	std_logic	:=	'0';
		lpbk_data_in	:	in	std_logic_vector(33 downto 0)	:=	"0000000000000000000000000000000000";
		lpbk_data_valid	:	in	std_logic	:=	'0';
		lpbk_en	:	in	std_logic	:=	'0';
		sync_in	:	in	std_logic_vector(1 downto 0)	:=	"00";
		tx_pma_clk	:	in	std_logic	:=	'0';
		tx_rstn	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		data_out	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		par_lpbk_b4gb_out	:	out	std_logic_vector(35 downto 0)	:=	"000000000000000000000000000000000000";
		par_lpbk_out	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		tx_test_out	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000"
	);
end twentynm_hssi_gen3_tx_pcs;

architecture behavior of twentynm_hssi_gen3_tx_pcs	is

constant tx_bitslip_int	:	integer	:=	bin2int(tx_bitslip);



component	twentynm_hssi_gen3_tx_pcs_encrypted
	generic (
		-- Architecture parameters
		mode	:	string	:=	"gen3_func";
		reverse_lpbk	:	string	:=	"rev_lpbk_en";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode";
		tx_bitslip	:	integer	:=	0;
		tx_gbox_byp	:	string	:=	"bypass_gbox"
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		blk_start_in	:	in	std_logic	:=	'0';
		data_in	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		data_valid	:	in	std_logic	:=	'0';
		lpbk_blk_start	:	in	std_logic	:=	'0';
		lpbk_data_in	:	in	std_logic_vector(33 downto 0)	:=	"0000000000000000000000000000000000";
		lpbk_data_valid	:	in	std_logic	:=	'0';
		lpbk_en	:	in	std_logic	:=	'0';
		sync_in	:	in	std_logic_vector(1 downto 0)	:=	"00";
		tx_pma_clk	:	in	std_logic	:=	'0';
		tx_rstn	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		data_out	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		par_lpbk_b4gb_out	:	out	std_logic_vector(35 downto 0)	:=	"000000000000000000000000000000000000";
		par_lpbk_out	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		tx_test_out	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000"
	);
end component;

begin



inst : twentynm_hssi_gen3_tx_pcs_encrypted
	generic map (
		-- Instance parameters
		mode	=>	mode,
		reverse_lpbk	=>	reverse_lpbk,
		silicon_rev	=>	silicon_rev,
		sup_mode	=>	sup_mode,
		tx_bitslip	=>	tx_bitslip_int,
		tx_gbox_byp	=>	tx_gbox_byp
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		blk_start_in	=>	blk_start_in,
		data_in	=>	data_in,
		data_valid	=>	data_valid,
		lpbk_blk_start	=>	lpbk_blk_start,
		lpbk_data_in	=>	lpbk_data_in,
		lpbk_data_valid	=>	lpbk_data_valid,
		lpbk_en	=>	lpbk_en,
		sync_in	=>	sync_in,
		tx_pma_clk	=>	tx_pma_clk,
		tx_rstn	=>	tx_rstn,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		data_out	=>	data_out,
		par_lpbk_b4gb_out	=>	par_lpbk_b4gb_out,
		par_lpbk_out	=>	par_lpbk_out,
		tx_test_out	=>	tx_test_out
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_gen3_x8_pcie_hip	is
	generic (
		-- Entity parameters
		acknack_base	:	bit_vector	:=	B"0000000000000";
		acknack_set	:	string	:=	"false";
		advance_error_reporting	:	string	:=	"disable";
		app_interface_width	:	string	:=	"avst_64bit";
		arb_upfc_30us_counter	:	bit_vector	:=	B"0000";
		arb_upfc_30us_en	:	string	:=	"enable";
		aspm_config_management	:	string	:=	"true";
		aspm_patch_disable	:	string	:=	"enable_both";
		ast_width_rx	:	string	:=	"rx_64";
		ast_width_tx	:	string	:=	"tx_64";
		atomic_malformed	:	string	:=	"false";
		atomic_op_completer_32bit	:	string	:=	"false";
		atomic_op_completer_64bit	:	string	:=	"false";
		atomic_op_routing	:	string	:=	"false";
		auto_msg_drop_enable	:	string	:=	"false";
		avmm_cvp_inter_sel_csr_ctrl	:	string	:=	"disable";
		avmm_dprio_broadcast_en_csr_ctrl	:	string	:=	"disable";
		avmm_force_inter_sel_csr_ctrl	:	string	:=	"disable";
		avmm_power_iso_en_csr_ctrl	:	string	:=	"disable";
		bar0_size_mask	:	bit_vector	:=	B"1111111111111111111111111111";
		bar0_type	:	string	:=	"bar0_64bit_prefetch_mem";
		bar1_size_mask	:	bit_vector	:=	B"0000000000000000000000000000";
		bar1_type	:	string	:=	"bar1_disable";
		bar2_size_mask	:	bit_vector	:=	B"0000000000000000000000000000";
		bar2_type	:	string	:=	"bar2_disable";
		bar3_size_mask	:	bit_vector	:=	B"0000000000000000000000000000";
		bar3_type	:	string	:=	"bar3_disable";
		bar4_size_mask	:	bit_vector	:=	B"0000000000000000000000000000";
		bar4_type	:	string	:=	"bar4_disable";
		bar5_size_mask	:	bit_vector	:=	B"0000000000000000000000000000";
		bar5_type	:	string	:=	"bar5_disable";
		base_counter_sel	:	string	:=	"count_clk_62p5";
		bist_memory_settings	:	string	:=	"000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		bridge_port_ssid_support	:	string	:=	"false";
		bridge_port_vga_enable	:	string	:=	"false";
		bypass_cdc	:	string	:=	"false";
		bypass_clk_switch	:	string	:=	"false";
		bypass_tl	:	string	:=	"false";
		capab_rate_rxcfg_en	:	string	:=	"disable";
		cas_completer_128bit	:	string	:=	"false";
		cdc_clk_relation	:	string	:=	"plesiochronous";
		cdc_dummy_insert_limit	:	bit_vector	:=	B"1011";
		cfg_parchk_ena	:	string	:=	"disable";
		cfgbp_req_recov_disable	:	string	:=	"false";
		class_code	:	bit_vector	:=	B"111111110000000000000000";
		clock_pwr_management	:	string	:=	"false";
		completion_timeout	:	string	:=	"abcd";
		core_clk_divider	:	string	:=	"div_1";
		core_clk_freq_mhz	:	string	:=	"core_clk_250mhz";
		core_clk_out_sel	:	string	:=	"core_clk_out_div_1";
		core_clk_sel	:	string	:=	"pld_clk";
		core_clk_source	:	string	:=	"pll_fixed_clk";
		cseb_bar_match_checking	:	string	:=	"enable";
		cseb_config_bypass	:	string	:=	"disable";
		cseb_cpl_status_during_cvp	:	string	:=	"completer_abort";
		cseb_cpl_tag_checking	:	string	:=	"enable";
		cseb_disable_auto_crs	:	string	:=	"false";
		cseb_extend_pci	:	string	:=	"false";
		cseb_extend_pcie	:	string	:=	"false";
		cseb_min_error_checking	:	string	:=	"false";
		cseb_route_to_avl_rx_st	:	string	:=	"cseb";
		cseb_temp_busy_crs	:	string	:=	"completer_abort_tmp_busy";
		cvp_clk_reset	:	string	:=	"false";
		cvp_data_compressed	:	string	:=	"false";
		cvp_data_encrypted	:	string	:=	"false";
		cvp_enable	:	string	:=	"cvp_dis";
		cvp_mode_reset	:	string	:=	"false";
		cvp_rate_sel	:	string	:=	"full_rate";
		d0_pme	:	string	:=	"false";
		d1_pme	:	string	:=	"false";
		d1_support	:	string	:=	"false";
		d2_pme	:	string	:=	"false";
		d2_support	:	string	:=	"false";
		d3_cold_pme	:	string	:=	"false";
		d3_hot_pme	:	string	:=	"false";
		data_pack_rx	:	string	:=	"disable";
		deemphasis_enable	:	string	:=	"false";
		deskew_comma	:	string	:=	"skp_eieos_deskw";
		device_id	:	bit_vector	:=	B"1110000000000001";
		device_number	:	bit_vector	:=	B"00000";
		device_specific_init	:	string	:=	"false";
		dft_clock_obsrv_en	:	string	:=	"disable";
		dft_clock_obsrv_sel	:	string	:=	"dft_pclk";
		diffclock_nfts_count	:	bit_vector	:=	B"00000000";
		dis_cplovf	:	string	:=	"disable";
		dis_paritychk	:	string	:=	"enable";
		disable_link_x2_support	:	string	:=	"false";
		disable_snoop_packet	:	string	:=	"false";
		dl_tx_check_parity_edb	:	string	:=	"disable";
		dll_active_report_support	:	string	:=	"false";
		early_dl_up	:	string	:=	"true";
		eco_fb332688_dis	:	string	:=	"true";
		ecrc_check_capable	:	string	:=	"true";
		ecrc_gen_capable	:	string	:=	"true";
		egress_block_err_report_ena	:	string	:=	"false";
		ei_delay_powerdown_count	:	bit_vector	:=	B"00001010";
		eie_before_nfts_count	:	bit_vector	:=	B"0100";
		electromech_interlock	:	string	:=	"false";
		en_ieiupdatefc	:	string	:=	"false";
		en_lane_errchk	:	string	:=	"false";
		en_phystatus_dly	:	string	:=	"false";
		ena_ido_cpl	:	string	:=	"false";
		ena_ido_req	:	string	:=	"false";
		enable_adapter_half_rate_mode	:	string	:=	"false";
		enable_ch01_pclk_out	:	string	:=	"pclk_ch0";
		enable_ch0_pclk_out	:	string	:=	"pclk_ch01";
		enable_completion_timeout_disable	:	string	:=	"true";
		enable_directed_spd_chng	:	string	:=	"false";
		enable_function_msix_support	:	string	:=	"true";
		enable_l0s_aspm	:	string	:=	"false";
		enable_l1_aspm	:	string	:=	"false";
		enable_rx_buffer_checking	:	string	:=	"false";
		enable_rx_reordering	:	string	:=	"true";
		enable_slot_register	:	string	:=	"false";
		endpoint_l0_latency	:	bit_vector	:=	B"000";
		endpoint_l1_latency	:	bit_vector	:=	B"000";
		eql_rq_int_en_number	:	bit_vector	:=	B"000000";
		errmgt_fcpe_patch_dis	:	string	:=	"enable";
		errmgt_fep_patch_dis	:	string	:=	"enable";
		expansion_base_address_register	:	string	:=	"00000000000000000000000000000000";
		extend_tag_field	:	string	:=	"false";
		extended_format_field	:	string	:=	"true";
		extended_tag_reset	:	string	:=	"false";
		fc_init_timer	:	bit_vector	:=	B"10000000000";
		flow_control_timeout_count	:	bit_vector	:=	B"11001000";
		flow_control_update_count	:	bit_vector	:=	B"11110";
		flr_capability	:	string	:=	"true";
		force_dis_to_det	:	string	:=	"false";
		force_gen1_dis	:	string	:=	"false";
		force_tx_coeff_preset_lpbk	:	string	:=	"false";
		frame_err_patch_dis	:	string	:=	"enable";
		func_mode	:	string	:=	"disable";
		g3_bypass_equlz	:	string	:=	"false";
		g3_coeff_done_tmout	:	string	:=	"enable";
		g3_deskew_char	:	string	:=	"default_sdsos";
		g3_dis_be_frm_err	:	string	:=	"false";
		g3_dn_rx_hint_eqlz_0	:	bit_vector	:=	B"000";
		g3_dn_rx_hint_eqlz_1	:	bit_vector	:=	B"000";
		g3_dn_rx_hint_eqlz_2	:	bit_vector	:=	B"000";
		g3_dn_rx_hint_eqlz_3	:	bit_vector	:=	B"000";
		g3_dn_rx_hint_eqlz_4	:	bit_vector	:=	B"000";
		g3_dn_rx_hint_eqlz_5	:	bit_vector	:=	B"000";
		g3_dn_rx_hint_eqlz_6	:	bit_vector	:=	B"000";
		g3_dn_rx_hint_eqlz_7	:	bit_vector	:=	B"000";
		g3_dn_tx_preset_eqlz_0	:	bit_vector	:=	B"0000";
		g3_dn_tx_preset_eqlz_1	:	bit_vector	:=	B"0000";
		g3_dn_tx_preset_eqlz_2	:	bit_vector	:=	B"0000";
		g3_dn_tx_preset_eqlz_3	:	bit_vector	:=	B"0000";
		g3_dn_tx_preset_eqlz_4	:	bit_vector	:=	B"0000";
		g3_dn_tx_preset_eqlz_5	:	bit_vector	:=	B"0000";
		g3_dn_tx_preset_eqlz_6	:	bit_vector	:=	B"0000";
		g3_dn_tx_preset_eqlz_7	:	bit_vector	:=	B"0000";
		g3_force_ber_max	:	string	:=	"false";
		g3_force_ber_min	:	string	:=	"false";
		g3_lnk_trn_rx_ts	:	string	:=	"false";
		g3_ltssm_eq_dbg	:	string	:=	"false";
		g3_ltssm_rec_dbg	:	string	:=	"false";
		g3_pause_ltssm_rec_en	:	string	:=	"disable";
		g3_quiesce_guarant	:	string	:=	"false";
		g3_redo_equlz_dis	:	string	:=	"false";
		g3_redo_equlz_en	:	string	:=	"false";
		g3_up_rx_hint_eqlz_0	:	bit_vector	:=	B"000";
		g3_up_rx_hint_eqlz_1	:	bit_vector	:=	B"000";
		g3_up_rx_hint_eqlz_2	:	bit_vector	:=	B"000";
		g3_up_rx_hint_eqlz_3	:	bit_vector	:=	B"000";
		g3_up_rx_hint_eqlz_4	:	bit_vector	:=	B"000";
		g3_up_rx_hint_eqlz_5	:	bit_vector	:=	B"000";
		g3_up_rx_hint_eqlz_6	:	bit_vector	:=	B"000";
		g3_up_rx_hint_eqlz_7	:	bit_vector	:=	B"000";
		g3_up_tx_preset_eqlz_0	:	bit_vector	:=	B"0000";
		g3_up_tx_preset_eqlz_1	:	bit_vector	:=	B"0000";
		g3_up_tx_preset_eqlz_2	:	bit_vector	:=	B"0000";
		g3_up_tx_preset_eqlz_3	:	bit_vector	:=	B"0000";
		g3_up_tx_preset_eqlz_4	:	bit_vector	:=	B"0000";
		g3_up_tx_preset_eqlz_5	:	bit_vector	:=	B"0000";
		g3_up_tx_preset_eqlz_6	:	bit_vector	:=	B"0000";
		g3_up_tx_preset_eqlz_7	:	bit_vector	:=	B"0000";
		gen123_lane_rate_mode	:	string	:=	"gen1_rate";
		gen2_diffclock_nfts_count	:	bit_vector	:=	B"11111111";
		gen2_pma_pll_usage	:	string	:=	"not_applicaple";
		gen2_sameclock_nfts_count	:	bit_vector	:=	B"11111111";
		gen3_coeff_1	:	bit_vector	:=	B"000000000000000100";
		gen3_coeff_10	:	bit_vector	:=	B"000000000000000111";
		gen3_coeff_10_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_10_nxtber_less	:	bit_vector	:=	B"1111";
		gen3_coeff_10_nxtber_more	:	bit_vector	:=	B"1010";
		gen3_coeff_10_preset_hint	:	bit_vector	:=	B"011";
		gen3_coeff_10_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_10_sel	:	string	:=	"preset_10";
		gen3_coeff_11	:	bit_vector	:=	B"000000000000000111";
		gen3_coeff_11_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_11_nxtber_less	:	bit_vector	:=	B"1111";
		gen3_coeff_11_nxtber_more	:	bit_vector	:=	B"1111";
		gen3_coeff_11_preset_hint	:	bit_vector	:=	B"100";
		gen3_coeff_11_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_11_sel	:	string	:=	"preset_11";
		gen3_coeff_12	:	bit_vector	:=	B"000000000000000111";
		gen3_coeff_12_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_12_nxtber_less	:	bit_vector	:=	B"1111";
		gen3_coeff_12_nxtber_more	:	bit_vector	:=	B"1111";
		gen3_coeff_12_preset_hint	:	bit_vector	:=	B"010";
		gen3_coeff_12_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_12_sel	:	string	:=	"preset_12";
		gen3_coeff_13	:	bit_vector	:=	B"000000000000000100";
		gen3_coeff_13_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_13_nxtber_less	:	bit_vector	:=	B"1101";
		gen3_coeff_13_nxtber_more	:	bit_vector	:=	B"0001";
		gen3_coeff_13_preset_hint	:	bit_vector	:=	B"100";
		gen3_coeff_13_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_13_sel	:	string	:=	"preset_13";
		gen3_coeff_14	:	bit_vector	:=	B"000000000000000100";
		gen3_coeff_14_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_14_nxtber_less	:	bit_vector	:=	B"1111";
		gen3_coeff_14_nxtber_more	:	bit_vector	:=	B"0010";
		gen3_coeff_14_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_14_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_14_sel	:	string	:=	"preset_14";
		gen3_coeff_15	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_15_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_15_nxtber_less	:	bit_vector	:=	B"0000";
		gen3_coeff_15_nxtber_more	:	bit_vector	:=	B"0000";
		gen3_coeff_15_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_15_reqber	:	bit_vector	:=	B"00000";
		gen3_coeff_15_sel	:	string	:=	"coeff_15";
		gen3_coeff_16	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_16_ber_meas	:	bit_vector	:=	B"000000";
		gen3_coeff_16_nxtber_less	:	bit_vector	:=	B"0000";
		gen3_coeff_16_nxtber_more	:	bit_vector	:=	B"0000";
		gen3_coeff_16_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_16_reqber	:	bit_vector	:=	B"00000";
		gen3_coeff_16_sel	:	string	:=	"coeff_16";
		gen3_coeff_17	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_17_ber_meas	:	bit_vector	:=	B"000000";
		gen3_coeff_17_nxtber_less	:	bit_vector	:=	B"0000";
		gen3_coeff_17_nxtber_more	:	bit_vector	:=	B"0000";
		gen3_coeff_17_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_17_reqber	:	bit_vector	:=	B"00000";
		gen3_coeff_17_sel	:	string	:=	"coeff_17";
		gen3_coeff_18	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_18_ber_meas	:	bit_vector	:=	B"000000";
		gen3_coeff_18_nxtber_less	:	bit_vector	:=	B"0000";
		gen3_coeff_18_nxtber_more	:	bit_vector	:=	B"0000";
		gen3_coeff_18_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_18_reqber	:	bit_vector	:=	B"00000";
		gen3_coeff_18_sel	:	string	:=	"coeff_18";
		gen3_coeff_19	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_19_ber_meas	:	bit_vector	:=	B"000000";
		gen3_coeff_19_nxtber_less	:	bit_vector	:=	B"0000";
		gen3_coeff_19_nxtber_more	:	bit_vector	:=	B"0000";
		gen3_coeff_19_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_19_reqber	:	bit_vector	:=	B"00000";
		gen3_coeff_19_sel	:	string	:=	"coeff_19";
		gen3_coeff_1_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_1_nxtber_less	:	bit_vector	:=	B"1100";
		gen3_coeff_1_nxtber_more	:	bit_vector	:=	B"0110";
		gen3_coeff_1_preset_hint	:	bit_vector	:=	B"010";
		gen3_coeff_1_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_1_sel	:	string	:=	"preset_1";
		gen3_coeff_2	:	bit_vector	:=	B"000000000000000001";
		gen3_coeff_20	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_20_ber_meas	:	bit_vector	:=	B"000000";
		gen3_coeff_20_nxtber_less	:	bit_vector	:=	B"0000";
		gen3_coeff_20_nxtber_more	:	bit_vector	:=	B"0000";
		gen3_coeff_20_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_20_reqber	:	bit_vector	:=	B"00000";
		gen3_coeff_20_sel	:	string	:=	"coeff_20";
		gen3_coeff_21	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_21_ber_meas	:	bit_vector	:=	B"000000";
		gen3_coeff_21_nxtber_less	:	bit_vector	:=	B"0000";
		gen3_coeff_21_nxtber_more	:	bit_vector	:=	B"0000";
		gen3_coeff_21_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_21_reqber	:	bit_vector	:=	B"00000";
		gen3_coeff_21_sel	:	string	:=	"coeff_21";
		gen3_coeff_22	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_22_ber_meas	:	bit_vector	:=	B"000000";
		gen3_coeff_22_nxtber_less	:	bit_vector	:=	B"0000";
		gen3_coeff_22_nxtber_more	:	bit_vector	:=	B"0000";
		gen3_coeff_22_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_22_reqber	:	bit_vector	:=	B"00000";
		gen3_coeff_22_sel	:	string	:=	"coeff_22";
		gen3_coeff_23	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_23_ber_meas	:	bit_vector	:=	B"000000";
		gen3_coeff_23_nxtber_less	:	bit_vector	:=	B"0000";
		gen3_coeff_23_nxtber_more	:	bit_vector	:=	B"0000";
		gen3_coeff_23_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_23_reqber	:	bit_vector	:=	B"00000";
		gen3_coeff_23_sel	:	string	:=	"coeff_23";
		gen3_coeff_24	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_24_ber_meas	:	bit_vector	:=	B"000000";
		gen3_coeff_24_nxtber_less	:	bit_vector	:=	B"0000";
		gen3_coeff_24_nxtber_more	:	bit_vector	:=	B"0000";
		gen3_coeff_24_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_24_reqber	:	bit_vector	:=	B"00000";
		gen3_coeff_24_sel	:	string	:=	"coeff_24";
		gen3_coeff_2_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_2_nxtber_less	:	bit_vector	:=	B"0010";
		gen3_coeff_2_nxtber_more	:	bit_vector	:=	B"0100";
		gen3_coeff_2_preset_hint	:	bit_vector	:=	B"100";
		gen3_coeff_2_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_2_sel	:	string	:=	"preset_2";
		gen3_coeff_3	:	bit_vector	:=	B"000000000000000001";
		gen3_coeff_3_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_3_nxtber_less	:	bit_vector	:=	B"1111";
		gen3_coeff_3_nxtber_more	:	bit_vector	:=	B"0011";
		gen3_coeff_3_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_3_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_3_sel	:	string	:=	"preset_3";
		gen3_coeff_4	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_4_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_4_nxtber_less	:	bit_vector	:=	B"1111";
		gen3_coeff_4_nxtber_more	:	bit_vector	:=	B"0100";
		gen3_coeff_4_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_4_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_4_sel	:	string	:=	"preset_4";
		gen3_coeff_5	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_5_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_5_nxtber_less	:	bit_vector	:=	B"1111";
		gen3_coeff_5_nxtber_more	:	bit_vector	:=	B"0101";
		gen3_coeff_5_preset_hint	:	bit_vector	:=	B"100";
		gen3_coeff_5_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_5_sel	:	string	:=	"preset_5";
		gen3_coeff_6	:	bit_vector	:=	B"000000000000000111";
		gen3_coeff_6_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_6_nxtber_less	:	bit_vector	:=	B"1111";
		gen3_coeff_6_nxtber_more	:	bit_vector	:=	B"1111";
		gen3_coeff_6_preset_hint	:	bit_vector	:=	B"100";
		gen3_coeff_6_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_6_sel	:	string	:=	"preset_6";
		gen3_coeff_7	:	bit_vector	:=	B"000000000000000001";
		gen3_coeff_7_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_7_nxtber_less	:	bit_vector	:=	B"0001";
		gen3_coeff_7_nxtber_more	:	bit_vector	:=	B"0111";
		gen3_coeff_7_preset_hint	:	bit_vector	:=	B"010";
		gen3_coeff_7_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_7_sel	:	string	:=	"preset_7";
		gen3_coeff_8	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_8_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_8_nxtber_less	:	bit_vector	:=	B"0100";
		gen3_coeff_8_nxtber_more	:	bit_vector	:=	B"1000";
		gen3_coeff_8_preset_hint	:	bit_vector	:=	B"010";
		gen3_coeff_8_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_8_sel	:	string	:=	"preset_8";
		gen3_coeff_9	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_9_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_9_nxtber_less	:	bit_vector	:=	B"1011";
		gen3_coeff_9_nxtber_more	:	bit_vector	:=	B"1001";
		gen3_coeff_9_preset_hint	:	bit_vector	:=	B"011";
		gen3_coeff_9_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_9_sel	:	string	:=	"preset_9";
		gen3_coeff_delay_count	:	bit_vector	:=	B"1111101";
		gen3_coeff_errchk	:	string	:=	"enable";
		gen3_dcbal_en	:	string	:=	"true";
		gen3_diffclock_nfts_count	:	bit_vector	:=	B"10000000";
		gen3_force_local_coeff	:	string	:=	"false";
		gen3_full_swing	:	bit_vector	:=	B"111111";
		gen3_half_swing	:	string	:=	"false";
		gen3_low_freq	:	bit_vector	:=	B"000001";
		gen3_paritychk	:	string	:=	"enable";
		gen3_pl_framing_err_dis	:	string	:=	"enable";
		gen3_preset_coeff_1	:	bit_vector	:=	B"000000110101001010";
		gen3_preset_coeff_10	:	bit_vector	:=	B"001011110100000000";
		gen3_preset_coeff_11	:	bit_vector	:=	B"011110100001000000";
		gen3_preset_coeff_2	:	bit_vector	:=	B"000000110100001011";
		gen3_preset_coeff_3	:	bit_vector	:=	B"000000110010001101";
		gen3_preset_coeff_4	:	bit_vector	:=	B"000000110111001000";
		gen3_preset_coeff_5	:	bit_vector	:=	B"000000111111000000";
		gen3_preset_coeff_6	:	bit_vector	:=	B"000110111001000000";
		gen3_preset_coeff_7	:	bit_vector	:=	B"001000110111000000";
		gen3_preset_coeff_8	:	bit_vector	:=	B"000110101100001101";
		gen3_preset_coeff_9	:	bit_vector	:=	B"001000101111001000";
		gen3_reset_eieos_cnt_bit	:	string	:=	"false";
		gen3_rxfreqlock_counter	:	bit_vector	:=	B"00000000000000000000";
		gen3_sameclock_nfts_count	:	bit_vector	:=	B"10000000";
		gen3_scrdscr_bypass	:	string	:=	"false";
		gen3_skip_ph2_ph3	:	string	:=	"false";
		hard_reset_bypass	:	string	:=	"false";
		hard_rst_sig_chnl_en	:	string	:=	"disable_hrc_sig";
		hard_rst_tx_pll_rst_chnl_en	:	string	:=	"disable_hrc_txpll_rst";
		hip_ac_pwr_clk_freq_in_hz	:	bit_vector	:=	B"000000000000000000000000000000";
		hip_ac_pwr_uw_per_mhz	:	bit_vector	:=	B"000000000000000000000000000000";
		hip_base_address	:	bit_vector	:=	B"0000000000";
		hip_clock_dis	:	string	:=	"enable_hip_clk";
		hip_hard_reset	:	string	:=	"enable";
		hip_pcs_sig_chnl_en	:	string	:=	"disable_hip_pcs_sig";
		hot_plug_support	:	bit_vector	:=	B"0000000";
		hrc_chnl_txpll_master_cgb_rst_select	:	string	:=	"disable_master_cgb_sel";
		hrdrstctrl_en	:	string	:=	"hrdrstctrl_dis";
		iei_enable_settings	:	string	:=	"gen3gen2_infei_infsd_gen1_infei_sd";
		indicator	:	bit_vector	:=	B"111";
		intel_id_access	:	string	:=	"false";
		interrupt_pin	:	string	:=	"inta";
		io_window_addr_width	:	string	:=	"window_32_bit";
		jtag_id	:	string	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		ko_compl_data	:	bit_vector	:=	B"000000000000";
		ko_compl_header	:	bit_vector	:=	B"000000000000";
		l01_entry_latency	:	bit_vector	:=	B"11111";
		l0_exit_latency_diffclock	:	bit_vector	:=	B"110";
		l0_exit_latency_sameclock	:	bit_vector	:=	B"110";
		l0s_adj_rply_timer_dis	:	string	:=	"enable";
		l1_exit_latency_diffclock	:	bit_vector	:=	B"000";
		l1_exit_latency_sameclock	:	bit_vector	:=	B"000";
		l2_async_logic	:	string	:=	"enable";
		lane_mask	:	string	:=	"ln_mask_x4";
		lane_rate	:	string	:=	"gen1";
		link_width	:	string	:=	"x1";
		lmi_hold_off_cfg_timer_en	:	string	:=	"disable";
		low_priority_vc	:	string	:=	"single_vc_low_pr";
		ltr_mechanism	:	string	:=	"false";
		ltssm_1ms_timeout	:	string	:=	"disable";
		ltssm_freqlocked_check	:	string	:=	"disable";
		malformed_tlp_truncate_en	:	string	:=	"disable";
		max_link_width	:	string	:=	"x4_link_width";
		max_payload_size	:	string	:=	"payload_512";
		maximum_current	:	bit_vector	:=	B"000";
		millisecond_cycle_count	:	bit_vector	:=	B"00000000000000000000";
		msi_64bit_addressing_capable	:	string	:=	"true";
		msi_masking_capable	:	string	:=	"false";
		msi_multi_message_capable	:	string	:=	"count_4";
		msi_support	:	string	:=	"true";
		msix_pba_bir	:	bit_vector	:=	B"000";
		msix_pba_offset	:	bit_vector	:=	B"00000000000000000000000000000";
		msix_table_bir	:	bit_vector	:=	B"000";
		msix_table_offset	:	bit_vector	:=	B"00000000000000000000000000000";
		msix_table_size	:	bit_vector	:=	B"00000000000";
		national_inst_thru_enhance	:	string	:=	"true";
		no_command_completed	:	string	:=	"true";
		no_soft_reset	:	string	:=	"false";
		not_use_k_gbl_bits	:	string	:=	"not_used_k_gbl";
		operating_voltage	:	string	:=	"standard";
		pcie_base_spec	:	string	:=	"pcie_2p1";
		pcie_mode	:	string	:=	"shared_mode";
		pcie_spec_1p0_compliance	:	string	:=	"spec_1p1";
		pcie_spec_version	:	string	:=	"v2";
		pclk_out_sel	:	string	:=	"pclk";
		pld_in_use_reg	:	string	:=	"false";
		pm_latency_patch_dis	:	string	:=	"enable";
		pm_txdl_patch_dis	:	string	:=	"enable";
		pme_clock	:	string	:=	"false";
		port_link_number	:	bit_vector	:=	B"00000001";
		port_type	:	string	:=	"native_ep";
		powerdown_mode	:	string	:=	"powerup";
		prefetchable_mem_window_addr_width	:	string	:=	"prefetch_32";
		r2c_mask_easy	:	string	:=	"false";
		r2c_mask_enable	:	string	:=	"false";
		rec_frqlk_mon_en	:	string	:=	"disable";
		register_pipe_signals	:	string	:=	"true";
		retry_buffer_last_active_address	:	bit_vector	:=	B"1111111111";
		retry_buffer_memory_settings	:	string	:=	"000000000000000000000000000000000000";
		retry_ecc_corr_mask_dis	:	string	:=	"enable";
		revision_id	:	bit_vector	:=	B"00000001";
		role_based_error_reporting	:	string	:=	"false";
		rp_bug_fix_pri_sec_stat_reg	:	bit_vector	:=	B"1111111";
		rpltim_base	:	bit_vector	:=	B"00000000000000";
		rpltim_set	:	string	:=	"false";
		rstctl_ltssm_dis	:	string	:=	"false";
		rstctrl_1ms_count_fref_clk	:	bit_vector	:=	B"00001111010000100100";
		rstctrl_1us_count_fref_clk	:	bit_vector	:=	B"00000000000000111111";
		rstctrl_altpe3_crst_n_inv	:	string	:=	"false";
		rstctrl_altpe3_rst_n_inv	:	string	:=	"false";
		rstctrl_altpe3_srst_n_inv	:	string	:=	"false";
		rstctrl_chnl_cal_done_select	:	string	:=	"not_active_chnl_cal_done";
		rstctrl_debug_en	:	string	:=	"false";
		rstctrl_force_inactive_rst	:	string	:=	"false";
		rstctrl_fref_clk_select	:	string	:=	"ch0_sel";
		rstctrl_hard_block_enable	:	string	:=	"hard_rst_ctl";
		rstctrl_hip_ep	:	string	:=	"hip_ep";
		rstctrl_mask_tx_pll_lock_select	:	string	:=	"not_active_mask_tx_pll_lock";
		rstctrl_perst_enable	:	string	:=	"level";
		rstctrl_perstn_select	:	string	:=	"perstn_pin";
		rstctrl_pld_clr	:	string	:=	"false";
		rstctrl_pll_cal_done_select	:	string	:=	"not_active_pll_cal_done";
		rstctrl_rx_pcs_rst_n_inv	:	string	:=	"false";
		rstctrl_rx_pcs_rst_n_select	:	string	:=	"not_active_rx_pcs_rst";
		rstctrl_rx_pll_freq_lock_select	:	string	:=	"not_active_rx_pll_f_lock";
		rstctrl_rx_pll_lock_select	:	string	:=	"not_active_rx_pll_lock";
		rstctrl_rx_pma_rstb_inv	:	string	:=	"false";
		rstctrl_rx_pma_rstb_select	:	string	:=	"not_active_rx_pma_rstb";
		rstctrl_timer_a	:	bit_vector	:=	B"00001010";
		rstctrl_timer_a_type	:	string	:=	"a_timer_milli_secs";
		rstctrl_timer_b	:	bit_vector	:=	B"00001010";
		rstctrl_timer_b_type	:	string	:=	"b_timer_milli_secs";
		rstctrl_timer_c	:	bit_vector	:=	B"00001010";
		rstctrl_timer_c_type	:	string	:=	"c_timer_milli_secs";
		rstctrl_timer_d	:	bit_vector	:=	B"00010100";
		rstctrl_timer_d_type	:	string	:=	"d_timer_milli_secs";
		rstctrl_timer_e	:	bit_vector	:=	B"00000001";
		rstctrl_timer_e_type	:	string	:=	"e_timer_milli_secs";
		rstctrl_timer_f	:	bit_vector	:=	B"00001010";
		rstctrl_timer_f_type	:	string	:=	"f_timer_milli_secs";
		rstctrl_timer_g	:	bit_vector	:=	B"00001010";
		rstctrl_timer_g_type	:	string	:=	"g_timer_milli_secs";
		rstctrl_timer_h	:	bit_vector	:=	B"00000100";
		rstctrl_timer_h_type	:	string	:=	"h_timer_milli_secs";
		rstctrl_timer_i	:	bit_vector	:=	B"00010100";
		rstctrl_timer_i_type	:	string	:=	"i_timer_milli_secs";
		rstctrl_timer_j	:	bit_vector	:=	B"00010100";
		rstctrl_timer_j_type	:	string	:=	"j_timer_milli_secs";
		rstctrl_tx_lcff_pll_lock_select	:	string	:=	"not_active_lcff_pll_lock";
		rstctrl_tx_lcff_pll_rstb_select	:	string	:=	"not_active_lcff_pll_rstb";
		rstctrl_tx_pcs_rst_n_inv	:	string	:=	"false";
		rstctrl_tx_pcs_rst_n_select	:	string	:=	"not_active_tx_pcs_rst";
		rstctrl_tx_pma_rstb_inv	:	string	:=	"false";
		rstctrl_tx_pma_syncp_inv	:	string	:=	"false";
		rstctrl_tx_pma_syncp_select	:	string	:=	"not_active_tx_pma_syncp";
		rx_ast_parity	:	string	:=	"disable";
		rx_buffer_credit_alloc	:	string	:=	"balance";
		rx_buffer_fc_protect	:	bit_vector	:=	B"00000000000001000100";
		rx_buffer_protect	:	bit_vector	:=	B"00001000100";
		rx_cdc_almost_empty	:	bit_vector	:=	B"0011";
		rx_cdc_almost_full	:	bit_vector	:=	B"1100";
		rx_cred_ctl_param	:	string	:=	"disable";
		rx_ei_l0s	:	string	:=	"disable";
		rx_l0s_count_idl	:	bit_vector	:=	B"00000000";
		rx_ptr0_nonposted_dpram_max	:	bit_vector	:=	B"00000000000";
		rx_ptr0_nonposted_dpram_min	:	bit_vector	:=	B"00000000000";
		rx_ptr0_posted_dpram_max	:	bit_vector	:=	B"00000000000";
		rx_ptr0_posted_dpram_min	:	bit_vector	:=	B"00000000000";
		rx_runt_patch_dis	:	string	:=	"enable";
		rx_sop_ctrl	:	string	:=	"rx_sop_boundary_64";
		rx_trunc_patch_dis	:	string	:=	"enable";
		rx_use_prst	:	string	:=	"false";
		rx_use_prst_ep	:	string	:=	"true";
		rxbuf_ecc_corr_mask_dis	:	string	:=	"enable";
		rxdl_bad_sop_eop_filter_dis	:	string	:=	"rxdlbug1_enable_both";
		rxdl_bad_tlp_patch_dis	:	string	:=	"rxdlbug2_enable_both";
		rxdl_lcrc_patch_dis	:	string	:=	"rxdlbug3_enable_both";
		sameclock_nfts_count	:	bit_vector	:=	B"00000000";
		sel_enable_pcs_rx_fifo_err	:	string	:=	"disable_sel";
		silicon_rev	:	string	:=	"20nm5es";
		sim_mode	:	string	:=	"disable";
		simple_ro_fifo_control_en	:	string	:=	"disable";
		single_rx_detect	:	string	:=	"detect_all_lanes";
		skp_os_gen3_count	:	bit_vector	:=	B"00000000000";
		skp_os_schedule_count	:	bit_vector	:=	B"00000000000";
		slot_number	:	bit_vector	:=	B"0000000000000";
		slot_power_limit	:	bit_vector	:=	B"00000000";
		slot_power_scale	:	bit_vector	:=	B"00";
		slotclk_cfg	:	string	:=	"static_slotclkcfgon";
		ssid	:	bit_vector	:=	B"0000000000000000";
		ssvid	:	bit_vector	:=	B"0000000000000000";
		subsystem_device_id	:	bit_vector	:=	B"1110000000000001";
		subsystem_vendor_id	:	bit_vector	:=	B"0001000101110010";
		sup_mode	:	string	:=	"user_mode";
		surprise_down_error_support	:	string	:=	"false";
		tl_cfg_div	:	string	:=	"cfg_clk_div_7";
		tl_tx_check_parity_msg	:	string	:=	"disable";
		tph_completer	:	string	:=	"false";
		tx_ast_parity	:	string	:=	"disable";
		tx_cdc_almost_empty	:	bit_vector	:=	B"0101";
		tx_cdc_almost_full	:	bit_vector	:=	B"1100";
		tx_sop_ctrl	:	string	:=	"boundary_64";
		tx_swing	:	bit_vector	:=	B"00000000";
		txdl_fair_arbiter_counter	:	bit_vector	:=	B"0000";
		txdl_fair_arbiter_en	:	string	:=	"enable";
		txrate_adv	:	string	:=	"capability";
		uc_calibration_en	:	string	:=	"uc_calibration_dis";
		use_aer	:	string	:=	"false";
		use_crc_forwarding	:	string	:=	"false";
		user_id	:	bit_vector	:=	B"0000000000000000";
		vc0_clk_enable	:	string	:=	"true";
		vc0_rx_buffer_memory_settings	:	string	:=	"000000000000000000000000000000000000";
		vc0_rx_flow_ctrl_compl_data	:	bit_vector	:=	B"000111000000";
		vc0_rx_flow_ctrl_compl_header	:	bit_vector	:=	B"01110000";
		vc0_rx_flow_ctrl_nonposted_data	:	bit_vector	:=	B"00000000";
		vc0_rx_flow_ctrl_nonposted_header	:	bit_vector	:=	B"00110110";
		vc0_rx_flow_ctrl_posted_data	:	bit_vector	:=	B"000101101000";
		vc0_rx_flow_ctrl_posted_header	:	bit_vector	:=	B"00110010";
		vc1_clk_enable	:	string	:=	"false";
		vc_arbitration	:	string	:=	"single_vc_arb";
		vc_enable	:	string	:=	"single_vc";
		vendor_id	:	bit_vector	:=	B"0001000101110010";
		vsec_cap	:	bit_vector	:=	B"0000";
		vsec_id	:	bit_vector	:=	B"0001000101110010";
		wrong_device_id	:	string	:=	"disable"
	);
	port (
		-- Entity ports
		aer_msi_num	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		app_int_err	:	in	std_logic_vector(1 downto 0)	:=	"00";
		app_inta_sts	:	in	std_logic	:=	'0';
		app_msi_num	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		app_msi_req	:	in	std_logic	:=	'0';
		app_msi_tc	:	in	std_logic_vector(2 downto 0)	:=	"000";
		atpg_los_en_n	:	in	std_logic	:=	'0';
		avmm_address	:	in	std_logic_vector(9 downto 0)	:=	"0000000000";
		avmm_byte_en	:	in	std_logic_vector(1 downto 0)	:=	"00";
		avmm_clk	:	in	std_logic	:=	'0';
		avmm_read	:	in	std_logic	:=	'0';
		avmm_rst_n	:	in	std_logic	:=	'0';
		avmm_write	:	in	std_logic	:=	'0';
		avmm_writedata	:	in	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		bist_scanen	:	in	std_logic	:=	'0';
		bist_scanin	:	in	std_logic	:=	'0';
		bisten_rcv_n	:	in	std_logic	:=	'0';
		bisten_rpl_n	:	in	std_logic	:=	'0';
		bistmode_n	:	in	std_logic	:=	'0';
		cfg_link2csr_pld	:	in	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		cfg_prmbus_pld	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		chnl_cal_done0	:	in	std_logic	:=	'0';
		chnl_cal_done1	:	in	std_logic	:=	'0';
		chnl_cal_done2	:	in	std_logic	:=	'0';
		chnl_cal_done3	:	in	std_logic	:=	'0';
		chnl_cal_done4	:	in	std_logic	:=	'0';
		chnl_cal_done5	:	in	std_logic	:=	'0';
		chnl_cal_done6	:	in	std_logic	:=	'0';
		chnl_cal_done7	:	in	std_logic	:=	'0';
		core_clk_in	:	in	std_logic	:=	'0';
		core_crst	:	in	std_logic	:=	'0';
		core_por	:	in	std_logic	:=	'0';
		core_rst	:	in	std_logic	:=	'0';
		core_srst	:	in	std_logic	:=	'0';
		cpl_err	:	in	std_logic_vector(6 downto 0)	:=	"0000000";
		cpl_pending	:	in	std_logic	:=	'0';
		cseb_rddata	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		cseb_rddata_parity	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		cseb_rdresponse	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		cseb_waitrequest	:	in	std_logic	:=	'0';
		cseb_wrresp_valid	:	in	std_logic	:=	'0';
		cseb_wrresponse	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		csr_cbdin	:	in	std_logic	:=	'0';
		csr_clk	:	in	std_logic	:=	'0';
		csr_din	:	in	std_logic	:=	'0';
		csr_en	:	in	std_logic	:=	'0';
		csr_enscan	:	in	std_logic	:=	'0';
		csr_entest	:	in	std_logic	:=	'0';
		csr_in	:	in	std_logic	:=	'0';
		csr_load_csr	:	in	std_logic	:=	'0';
		csr_pipe_in	:	in	std_logic	:=	'0';
		csr_seg	:	in	std_logic	:=	'0';
		csr_tcsrin	:	in	std_logic	:=	'0';
		csr_tverify	:	in	std_logic	:=	'0';
		cvp_config_done	:	in	std_logic	:=	'0';
		cvp_config_error	:	in	std_logic	:=	'0';
		cvp_config_ready	:	in	std_logic	:=	'0';
		cvp_en	:	in	std_logic	:=	'0';
		egress_blk_err	:	in	std_logic	:=	'0';
		entest	:	in	std_logic	:=	'0';
		flr_reset	:	in	std_logic	:=	'0';
		force_tx_eidle	:	in	std_logic	:=	'0';
		fref_clk0	:	in	std_logic	:=	'0';
		fref_clk1	:	in	std_logic	:=	'0';
		fref_clk2	:	in	std_logic	:=	'0';
		fref_clk3	:	in	std_logic	:=	'0';
		fref_clk4	:	in	std_logic	:=	'0';
		fref_clk5	:	in	std_logic	:=	'0';
		fref_clk6	:	in	std_logic	:=	'0';
		fref_clk7	:	in	std_logic	:=	'0';
		frzlogic	:	in	std_logic	:=	'0';
		frzreg	:	in	std_logic	:=	'0';
		hold_ltssm_rec	:	in	std_logic	:=	'0';
		hpg_ctrler	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		iocsrrdy_dly	:	in	std_logic	:=	'0';
		lmi_addr	:	in	std_logic_vector(11 downto 0)	:=	"000000000000";
		lmi_din	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		lmi_rden	:	in	std_logic	:=	'0';
		lmi_wren	:	in	std_logic	:=	'0';
		m10k_select	:	in	std_logic_vector(2 downto 0)	:=	"000";
		mask_tx_pll_lock0	:	in	std_logic	:=	'0';
		mask_tx_pll_lock1	:	in	std_logic	:=	'0';
		mask_tx_pll_lock2	:	in	std_logic	:=	'0';
		mask_tx_pll_lock3	:	in	std_logic	:=	'0';
		mask_tx_pll_lock4	:	in	std_logic	:=	'0';
		mask_tx_pll_lock5	:	in	std_logic	:=	'0';
		mask_tx_pll_lock6	:	in	std_logic	:=	'0';
		mask_tx_pll_lock7	:	in	std_logic	:=	'0';
		mem_hip_test_enable	:	in	std_logic	:=	'0';
		mem_regscanen_n	:	in	std_logic	:=	'0';
		mem_rscin_rcv_bot	:	in	std_logic	:=	'0';
		mem_rscin_rcv_top	:	in	std_logic	:=	'0';
		mem_rscin_rtry	:	in	std_logic	:=	'0';
		nfrzdrv	:	in	std_logic	:=	'0';
		npor	:	in	std_logic	:=	'0';
		pclk_central	:	in	std_logic	:=	'0';
		pclk_ch0	:	in	std_logic	:=	'0';
		pclk_ch1	:	in	std_logic	:=	'0';
		pex_msi_num	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		phy_rst	:	in	std_logic	:=	'0';
		phy_srst	:	in	std_logic	:=	'0';
		phystatus0	:	in	std_logic	:=	'0';
		phystatus1	:	in	std_logic	:=	'0';
		phystatus2	:	in	std_logic	:=	'0';
		phystatus3	:	in	std_logic	:=	'0';
		phystatus4	:	in	std_logic	:=	'0';
		phystatus5	:	in	std_logic	:=	'0';
		phystatus6	:	in	std_logic	:=	'0';
		phystatus7	:	in	std_logic	:=	'0';
		pin_perst_n	:	in	std_logic	:=	'0';
		pld_clk	:	in	std_logic	:=	'0';
		pld_clrhip_n	:	in	std_logic	:=	'0';
		pld_clrpcship_n	:	in	std_logic	:=	'0';
		pld_clrpmapcship_n	:	in	std_logic	:=	'0';
		pld_core_ready	:	in	std_logic	:=	'0';
		pld_gp_status	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		pld_perst_n	:	in	std_logic	:=	'0';
		pll_cal_done0	:	in	std_logic	:=	'0';
		pll_cal_done1	:	in	std_logic	:=	'0';
		pll_cal_done2	:	in	std_logic	:=	'0';
		pll_cal_done3	:	in	std_logic	:=	'0';
		pll_cal_done4	:	in	std_logic	:=	'0';
		pll_cal_done5	:	in	std_logic	:=	'0';
		pll_cal_done6	:	in	std_logic	:=	'0';
		pll_cal_done7	:	in	std_logic	:=	'0';
		pll_fixed_clk_central	:	in	std_logic	:=	'0';
		pll_fixed_clk_ch0	:	in	std_logic	:=	'0';
		pll_fixed_clk_ch1	:	in	std_logic	:=	'0';
		plniotri	:	in	std_logic	:=	'0';
		pm_auxpwr	:	in	std_logic	:=	'0';
		pm_data	:	in	std_logic_vector(9 downto 0)	:=	"0000000000";
		pm_event	:	in	std_logic	:=	'0';
		pm_exit_d0_ack	:	in	std_logic	:=	'0';
		pme_to_cr	:	in	std_logic	:=	'0';
		reserved_clk_in	:	in	std_logic	:=	'0';
		reserved_in	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		rx_cred_ctl	:	in	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		rx_pll_freq_lock0	:	in	std_logic	:=	'0';
		rx_pll_freq_lock1	:	in	std_logic	:=	'0';
		rx_pll_freq_lock2	:	in	std_logic	:=	'0';
		rx_pll_freq_lock3	:	in	std_logic	:=	'0';
		rx_pll_freq_lock4	:	in	std_logic	:=	'0';
		rx_pll_freq_lock5	:	in	std_logic	:=	'0';
		rx_pll_freq_lock6	:	in	std_logic	:=	'0';
		rx_pll_freq_lock7	:	in	std_logic	:=	'0';
		rx_pll_phase_lock0	:	in	std_logic	:=	'0';
		rx_pll_phase_lock1	:	in	std_logic	:=	'0';
		rx_pll_phase_lock2	:	in	std_logic	:=	'0';
		rx_pll_phase_lock3	:	in	std_logic	:=	'0';
		rx_pll_phase_lock4	:	in	std_logic	:=	'0';
		rx_pll_phase_lock5	:	in	std_logic	:=	'0';
		rx_pll_phase_lock6	:	in	std_logic	:=	'0';
		rx_pll_phase_lock7	:	in	std_logic	:=	'0';
		rx_st_mask	:	in	std_logic	:=	'0';
		rx_st_ready	:	in	std_logic	:=	'0';
		rxblkst0	:	in	std_logic	:=	'0';
		rxblkst1	:	in	std_logic	:=	'0';
		rxblkst2	:	in	std_logic	:=	'0';
		rxblkst3	:	in	std_logic	:=	'0';
		rxblkst4	:	in	std_logic	:=	'0';
		rxblkst5	:	in	std_logic	:=	'0';
		rxblkst6	:	in	std_logic	:=	'0';
		rxblkst7	:	in	std_logic	:=	'0';
		rxdata0	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata1	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata2	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata3	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata4	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata5	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata6	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata7	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdatak0	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak1	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak2	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak3	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak4	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak5	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak6	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak7	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdataskip0	:	in	std_logic	:=	'0';
		rxdataskip1	:	in	std_logic	:=	'0';
		rxdataskip2	:	in	std_logic	:=	'0';
		rxdataskip3	:	in	std_logic	:=	'0';
		rxdataskip4	:	in	std_logic	:=	'0';
		rxdataskip5	:	in	std_logic	:=	'0';
		rxdataskip6	:	in	std_logic	:=	'0';
		rxdataskip7	:	in	std_logic	:=	'0';
		rxelecidle0	:	in	std_logic	:=	'0';
		rxelecidle1	:	in	std_logic	:=	'0';
		rxelecidle2	:	in	std_logic	:=	'0';
		rxelecidle3	:	in	std_logic	:=	'0';
		rxelecidle4	:	in	std_logic	:=	'0';
		rxelecidle5	:	in	std_logic	:=	'0';
		rxelecidle6	:	in	std_logic	:=	'0';
		rxelecidle7	:	in	std_logic	:=	'0';
		rxfreqlocked0	:	in	std_logic	:=	'0';
		rxfreqlocked1	:	in	std_logic	:=	'0';
		rxfreqlocked2	:	in	std_logic	:=	'0';
		rxfreqlocked3	:	in	std_logic	:=	'0';
		rxfreqlocked4	:	in	std_logic	:=	'0';
		rxfreqlocked5	:	in	std_logic	:=	'0';
		rxfreqlocked6	:	in	std_logic	:=	'0';
		rxfreqlocked7	:	in	std_logic	:=	'0';
		rxstatus0	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus1	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus2	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus3	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus4	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus5	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus6	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus7	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxsynchd0	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd1	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd2	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd3	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd4	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd5	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd6	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd7	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxvalid0	:	in	std_logic	:=	'0';
		rxvalid1	:	in	std_logic	:=	'0';
		rxvalid2	:	in	std_logic	:=	'0';
		rxvalid3	:	in	std_logic	:=	'0';
		rxvalid4	:	in	std_logic	:=	'0';
		rxvalid5	:	in	std_logic	:=	'0';
		rxvalid6	:	in	std_logic	:=	'0';
		rxvalid7	:	in	std_logic	:=	'0';
		scan_mode_n	:	in	std_logic	:=	'0';
		scan_shift_n	:	in	std_logic	:=	'0';
		sw_ctmod	:	in	std_logic_vector(1 downto 0)	:=	"00";
		swdn_in	:	in	std_logic_vector(2 downto 0)	:=	"000";
		swup_in	:	in	std_logic_vector(6 downto 0)	:=	"0000000";
		test_in_1_hip	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		test_in_hip	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		test_pl_dbg_eqin	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		tx_cred_cons_select	:	in	std_logic	:=	'0';
		tx_cred_fc_sel	:	in	std_logic_vector(1 downto 0)	:=	"00";
		tx_lcff_pll_lock0	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock1	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock2	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock3	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock4	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock5	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock6	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock7	:	in	std_logic	:=	'0';
		tx_st_data	:	in	std_logic_vector(255 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		tx_st_empty	:	in	std_logic_vector(1 downto 0)	:=	"00";
		tx_st_eop	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		tx_st_err	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		tx_st_parity	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		tx_st_sop	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		tx_st_valid	:	in	std_logic	:=	'0';
		user_mode	:	in	std_logic	:=	'0';
		sta_hd_altpe3_hip_core_top_hd_altpe3_hip_core_u_clkmux_core_clk_cnt_reg_0_0_Q	:	out	std_logic	:=	'0';
		sta_hd_altpe3_hip_core_top_hd_altpe3_hip_core_u_clkmux_core_clk_cnt_reg_1_0_Q	:	out	std_logic	:=	'0';
		sta_hd_altpe3_hip_core_top_hd_altpe3_hip_core_u_clkmux_core_clk_cnt_reg_2_0_Q	:	out	std_logic	:=	'0';
		app_inta_ack	:	out	std_logic	:=	'0';
		app_msi_ack	:	out	std_logic	:=	'0';
		avmm_readdata	:	out	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		cfg_par_err	:	out	std_logic	:=	'0';
		core_clk_out	:	out	std_logic	:=	'0';
		cseb_addr	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		cseb_addr_parity	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		cseb_be	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		cseb_is_shadow	:	out	std_logic	:=	'0';
		cseb_rden	:	out	std_logic	:=	'0';
		cseb_wrdata	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		cseb_wrdata_parity	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		cseb_wren	:	out	std_logic	:=	'0';
		cseb_wrresp_req	:	out	std_logic	:=	'0';
		csr_dout	:	out	std_logic	:=	'0';
		csr_out	:	out	std_logic	:=	'0';
		csr_pipe_out	:	out	std_logic	:=	'0';
		current_coeff0	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff1	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff2	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff3	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff4	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff5	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff6	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff7	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_rxpreset0	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset1	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset2	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset3	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset4	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset5	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset6	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset7	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_speed	:	out	std_logic_vector(1 downto 0)	:=	"00";
		cvp_clk	:	out	std_logic	:=	'0';
		cvp_config	:	out	std_logic	:=	'0';
		cvp_data	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		cvp_full_config	:	out	std_logic	:=	'0';
		cvp_start_xfer	:	out	std_logic	:=	'0';
		dl_up	:	out	std_logic	:=	'0';
		dlup_exit	:	out	std_logic	:=	'0';
		eidle_infer_sel0	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel1	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel2	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel3	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel4	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel5	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel6	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel7	:	out	std_logic_vector(2 downto 0)	:=	"000";
		ev_128ns	:	out	std_logic	:=	'0';
		ev_1us	:	out	std_logic	:=	'0';
		flr_sts	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n0	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n1	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n2	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n3	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n4	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n5	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n6	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n7	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n0	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n1	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n2	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n3	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n4	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n5	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n6	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n7	:	out	std_logic	:=	'0';
		hotrst_exit	:	out	std_logic	:=	'0';
		int_status	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		k_hip_pcs_chnl_en	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		k_hrc_chnl_en	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		k_hrc_chnl_txpll_master_cgb_rst_en	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		k_hrc_chnl_txpll_rst_en	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		l2_exit	:	out	std_logic	:=	'0';
		lane_act	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		lmi_ack	:	out	std_logic	:=	'0';
		lmi_dout	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		ltssm_state	:	out	std_logic_vector(4 downto 0)	:=	"00000";
		mem_rscout_rcv_bot	:	out	std_logic	:=	'0';
		mem_rscout_rcv_top	:	out	std_logic	:=	'0';
		mem_rscout_rtry	:	out	std_logic	:=	'0';
		pld_clk_in_use	:	out	std_logic	:=	'0';
		pld_gp_ctrl	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		pm_exit_d0_req	:	out	std_logic	:=	'0';
		pme_to_sr	:	out	std_logic	:=	'0';
		powerdown0	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown1	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown2	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown3	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown4	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown5	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown6	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown7	:	out	std_logic_vector(1 downto 0)	:=	"00";
		r2c_unc_ecc	:	out	std_logic	:=	'0';
		rate0	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate1	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate2	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate3	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate4	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate5	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate6	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate7	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate_ctrl	:	out	std_logic_vector(1 downto 0)	:=	"00";
		reserved_clk_out	:	out	std_logic	:=	'0';
		reserved_out	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		reset_status	:	out	std_logic	:=	'0';
		retry_corr_ecc	:	out	std_logic	:=	'0';
		retry_unc_ecc	:	out	std_logic	:=	'0';
		rx_corr_ecc	:	out	std_logic	:=	'0';
		rx_cred_status	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		rx_par_err	:	out	std_logic	:=	'0';
		rx_pcs_rst_n0	:	out	std_logic	:=	'0';
		rx_pcs_rst_n1	:	out	std_logic	:=	'0';
		rx_pcs_rst_n2	:	out	std_logic	:=	'0';
		rx_pcs_rst_n3	:	out	std_logic	:=	'0';
		rx_pcs_rst_n4	:	out	std_logic	:=	'0';
		rx_pcs_rst_n5	:	out	std_logic	:=	'0';
		rx_pcs_rst_n6	:	out	std_logic	:=	'0';
		rx_pcs_rst_n7	:	out	std_logic	:=	'0';
		rx_pma_rstb0	:	out	std_logic	:=	'0';
		rx_pma_rstb1	:	out	std_logic	:=	'0';
		rx_pma_rstb2	:	out	std_logic	:=	'0';
		rx_pma_rstb3	:	out	std_logic	:=	'0';
		rx_pma_rstb4	:	out	std_logic	:=	'0';
		rx_pma_rstb5	:	out	std_logic	:=	'0';
		rx_pma_rstb6	:	out	std_logic	:=	'0';
		rx_pma_rstb7	:	out	std_logic	:=	'0';
		rx_st_bardec1	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		rx_st_bardec2	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		rx_st_be	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rx_st_data	:	out	std_logic_vector(255 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		rx_st_empty	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rx_st_eop	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		rx_st_err	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		rx_st_parity	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rx_st_sop	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		rx_st_valid	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		rxfc_cplbuf_ovf	:	out	std_logic	:=	'0';
		rxfc_cplovf_tag	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		rxpolarity0	:	out	std_logic	:=	'0';
		rxpolarity1	:	out	std_logic	:=	'0';
		rxpolarity2	:	out	std_logic	:=	'0';
		rxpolarity3	:	out	std_logic	:=	'0';
		rxpolarity4	:	out	std_logic	:=	'0';
		rxpolarity5	:	out	std_logic	:=	'0';
		rxpolarity6	:	out	std_logic	:=	'0';
		rxpolarity7	:	out	std_logic	:=	'0';
		serr_out	:	out	std_logic	:=	'0';
		swdn_out	:	out	std_logic_vector(6 downto 0)	:=	"0000000";
		swup_out	:	out	std_logic_vector(2 downto 0)	:=	"000";
		test_fref_clk	:	out	std_logic	:=	'0';
		test_out_1_hip	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		test_out_hip	:	out	std_logic_vector(255 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		tl_cfg_add	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		tl_cfg_ctl	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		tl_cfg_sts	:	out	std_logic_vector(52 downto 0)	:=	"00000000000000000000000000000000000000000000000000000";
		tl_cfg_sts_wr	:	out	std_logic	:=	'0';
		tx_cred_data_fc	:	out	std_logic_vector(11 downto 0)	:=	"000000000000";
		tx_cred_fc_hip_cons	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		tx_cred_fc_infinite	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		tx_cred_hdr_fc	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		tx_deemph0	:	out	std_logic	:=	'0';
		tx_deemph1	:	out	std_logic	:=	'0';
		tx_deemph2	:	out	std_logic	:=	'0';
		tx_deemph3	:	out	std_logic	:=	'0';
		tx_deemph4	:	out	std_logic	:=	'0';
		tx_deemph5	:	out	std_logic	:=	'0';
		tx_deemph6	:	out	std_logic	:=	'0';
		tx_deemph7	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb0	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb1	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb2	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb3	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb4	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb5	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb6	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb7	:	out	std_logic	:=	'0';
		tx_margin0	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin1	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin2	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin3	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin4	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin5	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin6	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin7	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_par_err	:	out	std_logic_vector(1 downto 0)	:=	"00";
		tx_pcs_rst_n0	:	out	std_logic	:=	'0';
		tx_pcs_rst_n1	:	out	std_logic	:=	'0';
		tx_pcs_rst_n2	:	out	std_logic	:=	'0';
		tx_pcs_rst_n3	:	out	std_logic	:=	'0';
		tx_pcs_rst_n4	:	out	std_logic	:=	'0';
		tx_pcs_rst_n5	:	out	std_logic	:=	'0';
		tx_pcs_rst_n6	:	out	std_logic	:=	'0';
		tx_pcs_rst_n7	:	out	std_logic	:=	'0';
		tx_pma_syncp0	:	out	std_logic	:=	'0';
		tx_pma_syncp1	:	out	std_logic	:=	'0';
		tx_pma_syncp2	:	out	std_logic	:=	'0';
		tx_pma_syncp3	:	out	std_logic	:=	'0';
		tx_pma_syncp4	:	out	std_logic	:=	'0';
		tx_pma_syncp5	:	out	std_logic	:=	'0';
		tx_pma_syncp6	:	out	std_logic	:=	'0';
		tx_pma_syncp7	:	out	std_logic	:=	'0';
		tx_st_ready	:	out	std_logic	:=	'0';
		txblkst0	:	out	std_logic	:=	'0';
		txblkst1	:	out	std_logic	:=	'0';
		txblkst2	:	out	std_logic	:=	'0';
		txblkst3	:	out	std_logic	:=	'0';
		txblkst4	:	out	std_logic	:=	'0';
		txblkst5	:	out	std_logic	:=	'0';
		txblkst6	:	out	std_logic	:=	'0';
		txblkst7	:	out	std_logic	:=	'0';
		txcompl0	:	out	std_logic	:=	'0';
		txcompl1	:	out	std_logic	:=	'0';
		txcompl2	:	out	std_logic	:=	'0';
		txcompl3	:	out	std_logic	:=	'0';
		txcompl4	:	out	std_logic	:=	'0';
		txcompl5	:	out	std_logic	:=	'0';
		txcompl6	:	out	std_logic	:=	'0';
		txcompl7	:	out	std_logic	:=	'0';
		txdata0	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata1	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata2	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata3	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata4	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata5	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata6	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata7	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdatak0	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak1	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak2	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak3	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak4	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak5	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak6	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak7	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdataskip0	:	out	std_logic	:=	'0';
		txdataskip1	:	out	std_logic	:=	'0';
		txdataskip2	:	out	std_logic	:=	'0';
		txdataskip3	:	out	std_logic	:=	'0';
		txdataskip4	:	out	std_logic	:=	'0';
		txdataskip5	:	out	std_logic	:=	'0';
		txdataskip6	:	out	std_logic	:=	'0';
		txdataskip7	:	out	std_logic	:=	'0';
		txdetectrx0	:	out	std_logic	:=	'0';
		txdetectrx1	:	out	std_logic	:=	'0';
		txdetectrx2	:	out	std_logic	:=	'0';
		txdetectrx3	:	out	std_logic	:=	'0';
		txdetectrx4	:	out	std_logic	:=	'0';
		txdetectrx5	:	out	std_logic	:=	'0';
		txdetectrx6	:	out	std_logic	:=	'0';
		txdetectrx7	:	out	std_logic	:=	'0';
		txelecidle0	:	out	std_logic	:=	'0';
		txelecidle1	:	out	std_logic	:=	'0';
		txelecidle2	:	out	std_logic	:=	'0';
		txelecidle3	:	out	std_logic	:=	'0';
		txelecidle4	:	out	std_logic	:=	'0';
		txelecidle5	:	out	std_logic	:=	'0';
		txelecidle6	:	out	std_logic	:=	'0';
		txelecidle7	:	out	std_logic	:=	'0';
		txst_prot_err	:	out	std_logic	:=	'0';
		txswing0	:	out	std_logic	:=	'0';
		txswing1	:	out	std_logic	:=	'0';
		txswing2	:	out	std_logic	:=	'0';
		txswing3	:	out	std_logic	:=	'0';
		txswing4	:	out	std_logic	:=	'0';
		txswing5	:	out	std_logic	:=	'0';
		txswing6	:	out	std_logic	:=	'0';
		txswing7	:	out	std_logic	:=	'0';
		txsynchd0	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd1	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd2	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd3	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd4	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd5	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd6	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd7	:	out	std_logic_vector(1 downto 0)	:=	"00";
		wake_oen	:	out	std_logic	:=	'0'
	);
end twentynm_hssi_gen3_x8_pcie_hip;

architecture behavior of twentynm_hssi_gen3_x8_pcie_hip	is

constant acknack_base_int	:	integer	:=	bin2int(acknack_base);
constant arb_upfc_30us_counter_int	:	integer	:=	bin2int(arb_upfc_30us_counter);
constant bar0_size_mask_int	:	integer	:=	bin2int(bar0_size_mask);
constant bar1_size_mask_int	:	integer	:=	bin2int(bar1_size_mask);
constant bar2_size_mask_int	:	integer	:=	bin2int(bar2_size_mask);
constant bar3_size_mask_int	:	integer	:=	bin2int(bar3_size_mask);
constant bar4_size_mask_int	:	integer	:=	bin2int(bar4_size_mask);
constant bar5_size_mask_int	:	integer	:=	bin2int(bar5_size_mask);
constant cdc_dummy_insert_limit_int	:	integer	:=	bin2int(cdc_dummy_insert_limit);
constant class_code_int	:	integer	:=	bin2int(class_code);
constant device_id_int	:	integer	:=	bin2int(device_id);
constant device_number_int	:	integer	:=	bin2int(device_number);
constant diffclock_nfts_count_int	:	integer	:=	bin2int(diffclock_nfts_count);
constant ei_delay_powerdown_count_int	:	integer	:=	bin2int(ei_delay_powerdown_count);
constant eie_before_nfts_count_int	:	integer	:=	bin2int(eie_before_nfts_count);
constant endpoint_l0_latency_int	:	integer	:=	bin2int(endpoint_l0_latency);
constant endpoint_l1_latency_int	:	integer	:=	bin2int(endpoint_l1_latency);
constant eql_rq_int_en_number_int	:	integer	:=	bin2int(eql_rq_int_en_number);
constant fc_init_timer_int	:	integer	:=	bin2int(fc_init_timer);
constant flow_control_timeout_count_int	:	integer	:=	bin2int(flow_control_timeout_count);
constant flow_control_update_count_int	:	integer	:=	bin2int(flow_control_update_count);
constant g3_dn_rx_hint_eqlz_0_int	:	integer	:=	bin2int(g3_dn_rx_hint_eqlz_0);
constant g3_dn_rx_hint_eqlz_1_int	:	integer	:=	bin2int(g3_dn_rx_hint_eqlz_1);
constant g3_dn_rx_hint_eqlz_2_int	:	integer	:=	bin2int(g3_dn_rx_hint_eqlz_2);
constant g3_dn_rx_hint_eqlz_3_int	:	integer	:=	bin2int(g3_dn_rx_hint_eqlz_3);
constant g3_dn_rx_hint_eqlz_4_int	:	integer	:=	bin2int(g3_dn_rx_hint_eqlz_4);
constant g3_dn_rx_hint_eqlz_5_int	:	integer	:=	bin2int(g3_dn_rx_hint_eqlz_5);
constant g3_dn_rx_hint_eqlz_6_int	:	integer	:=	bin2int(g3_dn_rx_hint_eqlz_6);
constant g3_dn_rx_hint_eqlz_7_int	:	integer	:=	bin2int(g3_dn_rx_hint_eqlz_7);
constant g3_dn_tx_preset_eqlz_0_int	:	integer	:=	bin2int(g3_dn_tx_preset_eqlz_0);
constant g3_dn_tx_preset_eqlz_1_int	:	integer	:=	bin2int(g3_dn_tx_preset_eqlz_1);
constant g3_dn_tx_preset_eqlz_2_int	:	integer	:=	bin2int(g3_dn_tx_preset_eqlz_2);
constant g3_dn_tx_preset_eqlz_3_int	:	integer	:=	bin2int(g3_dn_tx_preset_eqlz_3);
constant g3_dn_tx_preset_eqlz_4_int	:	integer	:=	bin2int(g3_dn_tx_preset_eqlz_4);
constant g3_dn_tx_preset_eqlz_5_int	:	integer	:=	bin2int(g3_dn_tx_preset_eqlz_5);
constant g3_dn_tx_preset_eqlz_6_int	:	integer	:=	bin2int(g3_dn_tx_preset_eqlz_6);
constant g3_dn_tx_preset_eqlz_7_int	:	integer	:=	bin2int(g3_dn_tx_preset_eqlz_7);
constant g3_up_rx_hint_eqlz_0_int	:	integer	:=	bin2int(g3_up_rx_hint_eqlz_0);
constant g3_up_rx_hint_eqlz_1_int	:	integer	:=	bin2int(g3_up_rx_hint_eqlz_1);
constant g3_up_rx_hint_eqlz_2_int	:	integer	:=	bin2int(g3_up_rx_hint_eqlz_2);
constant g3_up_rx_hint_eqlz_3_int	:	integer	:=	bin2int(g3_up_rx_hint_eqlz_3);
constant g3_up_rx_hint_eqlz_4_int	:	integer	:=	bin2int(g3_up_rx_hint_eqlz_4);
constant g3_up_rx_hint_eqlz_5_int	:	integer	:=	bin2int(g3_up_rx_hint_eqlz_5);
constant g3_up_rx_hint_eqlz_6_int	:	integer	:=	bin2int(g3_up_rx_hint_eqlz_6);
constant g3_up_rx_hint_eqlz_7_int	:	integer	:=	bin2int(g3_up_rx_hint_eqlz_7);
constant g3_up_tx_preset_eqlz_0_int	:	integer	:=	bin2int(g3_up_tx_preset_eqlz_0);
constant g3_up_tx_preset_eqlz_1_int	:	integer	:=	bin2int(g3_up_tx_preset_eqlz_1);
constant g3_up_tx_preset_eqlz_2_int	:	integer	:=	bin2int(g3_up_tx_preset_eqlz_2);
constant g3_up_tx_preset_eqlz_3_int	:	integer	:=	bin2int(g3_up_tx_preset_eqlz_3);
constant g3_up_tx_preset_eqlz_4_int	:	integer	:=	bin2int(g3_up_tx_preset_eqlz_4);
constant g3_up_tx_preset_eqlz_5_int	:	integer	:=	bin2int(g3_up_tx_preset_eqlz_5);
constant g3_up_tx_preset_eqlz_6_int	:	integer	:=	bin2int(g3_up_tx_preset_eqlz_6);
constant g3_up_tx_preset_eqlz_7_int	:	integer	:=	bin2int(g3_up_tx_preset_eqlz_7);
constant gen2_diffclock_nfts_count_int	:	integer	:=	bin2int(gen2_diffclock_nfts_count);
constant gen2_sameclock_nfts_count_int	:	integer	:=	bin2int(gen2_sameclock_nfts_count);
constant gen3_coeff_1_int	:	integer	:=	bin2int(gen3_coeff_1);
constant gen3_coeff_10_int	:	integer	:=	bin2int(gen3_coeff_10);
constant gen3_coeff_10_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_10_ber_meas);
constant gen3_coeff_10_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_10_nxtber_less);
constant gen3_coeff_10_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_10_nxtber_more);
constant gen3_coeff_10_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_10_preset_hint);
constant gen3_coeff_10_reqber_int	:	integer	:=	bin2int(gen3_coeff_10_reqber);
constant gen3_coeff_11_int	:	integer	:=	bin2int(gen3_coeff_11);
constant gen3_coeff_11_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_11_ber_meas);
constant gen3_coeff_11_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_11_nxtber_less);
constant gen3_coeff_11_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_11_nxtber_more);
constant gen3_coeff_11_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_11_preset_hint);
constant gen3_coeff_11_reqber_int	:	integer	:=	bin2int(gen3_coeff_11_reqber);
constant gen3_coeff_12_int	:	integer	:=	bin2int(gen3_coeff_12);
constant gen3_coeff_12_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_12_ber_meas);
constant gen3_coeff_12_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_12_nxtber_less);
constant gen3_coeff_12_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_12_nxtber_more);
constant gen3_coeff_12_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_12_preset_hint);
constant gen3_coeff_12_reqber_int	:	integer	:=	bin2int(gen3_coeff_12_reqber);
constant gen3_coeff_13_int	:	integer	:=	bin2int(gen3_coeff_13);
constant gen3_coeff_13_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_13_ber_meas);
constant gen3_coeff_13_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_13_nxtber_less);
constant gen3_coeff_13_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_13_nxtber_more);
constant gen3_coeff_13_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_13_preset_hint);
constant gen3_coeff_13_reqber_int	:	integer	:=	bin2int(gen3_coeff_13_reqber);
constant gen3_coeff_14_int	:	integer	:=	bin2int(gen3_coeff_14);
constant gen3_coeff_14_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_14_ber_meas);
constant gen3_coeff_14_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_14_nxtber_less);
constant gen3_coeff_14_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_14_nxtber_more);
constant gen3_coeff_14_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_14_preset_hint);
constant gen3_coeff_14_reqber_int	:	integer	:=	bin2int(gen3_coeff_14_reqber);
constant gen3_coeff_15_int	:	integer	:=	bin2int(gen3_coeff_15);
constant gen3_coeff_15_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_15_ber_meas);
constant gen3_coeff_15_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_15_nxtber_less);
constant gen3_coeff_15_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_15_nxtber_more);
constant gen3_coeff_15_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_15_preset_hint);
constant gen3_coeff_15_reqber_int	:	integer	:=	bin2int(gen3_coeff_15_reqber);
constant gen3_coeff_16_int	:	integer	:=	bin2int(gen3_coeff_16);
constant gen3_coeff_16_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_16_ber_meas);
constant gen3_coeff_16_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_16_nxtber_less);
constant gen3_coeff_16_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_16_nxtber_more);
constant gen3_coeff_16_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_16_preset_hint);
constant gen3_coeff_16_reqber_int	:	integer	:=	bin2int(gen3_coeff_16_reqber);
constant gen3_coeff_17_int	:	integer	:=	bin2int(gen3_coeff_17);
constant gen3_coeff_17_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_17_ber_meas);
constant gen3_coeff_17_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_17_nxtber_less);
constant gen3_coeff_17_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_17_nxtber_more);
constant gen3_coeff_17_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_17_preset_hint);
constant gen3_coeff_17_reqber_int	:	integer	:=	bin2int(gen3_coeff_17_reqber);
constant gen3_coeff_18_int	:	integer	:=	bin2int(gen3_coeff_18);
constant gen3_coeff_18_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_18_ber_meas);
constant gen3_coeff_18_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_18_nxtber_less);
constant gen3_coeff_18_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_18_nxtber_more);
constant gen3_coeff_18_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_18_preset_hint);
constant gen3_coeff_18_reqber_int	:	integer	:=	bin2int(gen3_coeff_18_reqber);
constant gen3_coeff_19_int	:	integer	:=	bin2int(gen3_coeff_19);
constant gen3_coeff_19_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_19_ber_meas);
constant gen3_coeff_19_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_19_nxtber_less);
constant gen3_coeff_19_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_19_nxtber_more);
constant gen3_coeff_19_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_19_preset_hint);
constant gen3_coeff_19_reqber_int	:	integer	:=	bin2int(gen3_coeff_19_reqber);
constant gen3_coeff_1_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_1_ber_meas);
constant gen3_coeff_1_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_1_nxtber_less);
constant gen3_coeff_1_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_1_nxtber_more);
constant gen3_coeff_1_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_1_preset_hint);
constant gen3_coeff_1_reqber_int	:	integer	:=	bin2int(gen3_coeff_1_reqber);
constant gen3_coeff_2_int	:	integer	:=	bin2int(gen3_coeff_2);
constant gen3_coeff_20_int	:	integer	:=	bin2int(gen3_coeff_20);
constant gen3_coeff_20_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_20_ber_meas);
constant gen3_coeff_20_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_20_nxtber_less);
constant gen3_coeff_20_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_20_nxtber_more);
constant gen3_coeff_20_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_20_preset_hint);
constant gen3_coeff_20_reqber_int	:	integer	:=	bin2int(gen3_coeff_20_reqber);
constant gen3_coeff_21_int	:	integer	:=	bin2int(gen3_coeff_21);
constant gen3_coeff_21_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_21_ber_meas);
constant gen3_coeff_21_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_21_nxtber_less);
constant gen3_coeff_21_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_21_nxtber_more);
constant gen3_coeff_21_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_21_preset_hint);
constant gen3_coeff_21_reqber_int	:	integer	:=	bin2int(gen3_coeff_21_reqber);
constant gen3_coeff_22_int	:	integer	:=	bin2int(gen3_coeff_22);
constant gen3_coeff_22_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_22_ber_meas);
constant gen3_coeff_22_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_22_nxtber_less);
constant gen3_coeff_22_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_22_nxtber_more);
constant gen3_coeff_22_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_22_preset_hint);
constant gen3_coeff_22_reqber_int	:	integer	:=	bin2int(gen3_coeff_22_reqber);
constant gen3_coeff_23_int	:	integer	:=	bin2int(gen3_coeff_23);
constant gen3_coeff_23_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_23_ber_meas);
constant gen3_coeff_23_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_23_nxtber_less);
constant gen3_coeff_23_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_23_nxtber_more);
constant gen3_coeff_23_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_23_preset_hint);
constant gen3_coeff_23_reqber_int	:	integer	:=	bin2int(gen3_coeff_23_reqber);
constant gen3_coeff_24_int	:	integer	:=	bin2int(gen3_coeff_24);
constant gen3_coeff_24_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_24_ber_meas);
constant gen3_coeff_24_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_24_nxtber_less);
constant gen3_coeff_24_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_24_nxtber_more);
constant gen3_coeff_24_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_24_preset_hint);
constant gen3_coeff_24_reqber_int	:	integer	:=	bin2int(gen3_coeff_24_reqber);
constant gen3_coeff_2_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_2_ber_meas);
constant gen3_coeff_2_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_2_nxtber_less);
constant gen3_coeff_2_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_2_nxtber_more);
constant gen3_coeff_2_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_2_preset_hint);
constant gen3_coeff_2_reqber_int	:	integer	:=	bin2int(gen3_coeff_2_reqber);
constant gen3_coeff_3_int	:	integer	:=	bin2int(gen3_coeff_3);
constant gen3_coeff_3_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_3_ber_meas);
constant gen3_coeff_3_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_3_nxtber_less);
constant gen3_coeff_3_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_3_nxtber_more);
constant gen3_coeff_3_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_3_preset_hint);
constant gen3_coeff_3_reqber_int	:	integer	:=	bin2int(gen3_coeff_3_reqber);
constant gen3_coeff_4_int	:	integer	:=	bin2int(gen3_coeff_4);
constant gen3_coeff_4_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_4_ber_meas);
constant gen3_coeff_4_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_4_nxtber_less);
constant gen3_coeff_4_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_4_nxtber_more);
constant gen3_coeff_4_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_4_preset_hint);
constant gen3_coeff_4_reqber_int	:	integer	:=	bin2int(gen3_coeff_4_reqber);
constant gen3_coeff_5_int	:	integer	:=	bin2int(gen3_coeff_5);
constant gen3_coeff_5_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_5_ber_meas);
constant gen3_coeff_5_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_5_nxtber_less);
constant gen3_coeff_5_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_5_nxtber_more);
constant gen3_coeff_5_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_5_preset_hint);
constant gen3_coeff_5_reqber_int	:	integer	:=	bin2int(gen3_coeff_5_reqber);
constant gen3_coeff_6_int	:	integer	:=	bin2int(gen3_coeff_6);
constant gen3_coeff_6_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_6_ber_meas);
constant gen3_coeff_6_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_6_nxtber_less);
constant gen3_coeff_6_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_6_nxtber_more);
constant gen3_coeff_6_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_6_preset_hint);
constant gen3_coeff_6_reqber_int	:	integer	:=	bin2int(gen3_coeff_6_reqber);
constant gen3_coeff_7_int	:	integer	:=	bin2int(gen3_coeff_7);
constant gen3_coeff_7_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_7_ber_meas);
constant gen3_coeff_7_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_7_nxtber_less);
constant gen3_coeff_7_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_7_nxtber_more);
constant gen3_coeff_7_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_7_preset_hint);
constant gen3_coeff_7_reqber_int	:	integer	:=	bin2int(gen3_coeff_7_reqber);
constant gen3_coeff_8_int	:	integer	:=	bin2int(gen3_coeff_8);
constant gen3_coeff_8_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_8_ber_meas);
constant gen3_coeff_8_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_8_nxtber_less);
constant gen3_coeff_8_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_8_nxtber_more);
constant gen3_coeff_8_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_8_preset_hint);
constant gen3_coeff_8_reqber_int	:	integer	:=	bin2int(gen3_coeff_8_reqber);
constant gen3_coeff_9_int	:	integer	:=	bin2int(gen3_coeff_9);
constant gen3_coeff_9_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_9_ber_meas);
constant gen3_coeff_9_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_9_nxtber_less);
constant gen3_coeff_9_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_9_nxtber_more);
constant gen3_coeff_9_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_9_preset_hint);
constant gen3_coeff_9_reqber_int	:	integer	:=	bin2int(gen3_coeff_9_reqber);
constant gen3_coeff_delay_count_int	:	integer	:=	bin2int(gen3_coeff_delay_count);
constant gen3_diffclock_nfts_count_int	:	integer	:=	bin2int(gen3_diffclock_nfts_count);
constant gen3_full_swing_int	:	integer	:=	bin2int(gen3_full_swing);
constant gen3_low_freq_int	:	integer	:=	bin2int(gen3_low_freq);
constant gen3_preset_coeff_1_int	:	integer	:=	bin2int(gen3_preset_coeff_1);
constant gen3_preset_coeff_10_int	:	integer	:=	bin2int(gen3_preset_coeff_10);
constant gen3_preset_coeff_11_int	:	integer	:=	bin2int(gen3_preset_coeff_11);
constant gen3_preset_coeff_2_int	:	integer	:=	bin2int(gen3_preset_coeff_2);
constant gen3_preset_coeff_3_int	:	integer	:=	bin2int(gen3_preset_coeff_3);
constant gen3_preset_coeff_4_int	:	integer	:=	bin2int(gen3_preset_coeff_4);
constant gen3_preset_coeff_5_int	:	integer	:=	bin2int(gen3_preset_coeff_5);
constant gen3_preset_coeff_6_int	:	integer	:=	bin2int(gen3_preset_coeff_6);
constant gen3_preset_coeff_7_int	:	integer	:=	bin2int(gen3_preset_coeff_7);
constant gen3_preset_coeff_8_int	:	integer	:=	bin2int(gen3_preset_coeff_8);
constant gen3_preset_coeff_9_int	:	integer	:=	bin2int(gen3_preset_coeff_9);
constant gen3_rxfreqlock_counter_int	:	integer	:=	bin2int(gen3_rxfreqlock_counter);
constant gen3_sameclock_nfts_count_int	:	integer	:=	bin2int(gen3_sameclock_nfts_count);
constant hip_ac_pwr_clk_freq_in_hz_int	:	integer	:=	bin2int(hip_ac_pwr_clk_freq_in_hz);
constant hip_ac_pwr_uw_per_mhz_int	:	integer	:=	bin2int(hip_ac_pwr_uw_per_mhz);
constant hip_base_address_int	:	integer	:=	bin2int(hip_base_address);
constant hot_plug_support_int	:	integer	:=	bin2int(hot_plug_support);
constant indicator_int	:	integer	:=	bin2int(indicator);
constant ko_compl_data_int	:	integer	:=	bin2int(ko_compl_data);
constant ko_compl_header_int	:	integer	:=	bin2int(ko_compl_header);
constant l01_entry_latency_int	:	integer	:=	bin2int(l01_entry_latency);
constant l0_exit_latency_diffclock_int	:	integer	:=	bin2int(l0_exit_latency_diffclock);
constant l0_exit_latency_sameclock_int	:	integer	:=	bin2int(l0_exit_latency_sameclock);
constant l1_exit_latency_diffclock_int	:	integer	:=	bin2int(l1_exit_latency_diffclock);
constant l1_exit_latency_sameclock_int	:	integer	:=	bin2int(l1_exit_latency_sameclock);
constant maximum_current_int	:	integer	:=	bin2int(maximum_current);
constant millisecond_cycle_count_int	:	integer	:=	bin2int(millisecond_cycle_count);
constant msix_pba_bir_int	:	integer	:=	bin2int(msix_pba_bir);
constant msix_pba_offset_int	:	integer	:=	bin2int(msix_pba_offset);
constant msix_table_bir_int	:	integer	:=	bin2int(msix_table_bir);
constant msix_table_offset_int	:	integer	:=	bin2int(msix_table_offset);
constant msix_table_size_int	:	integer	:=	bin2int(msix_table_size);
constant port_link_number_int	:	integer	:=	bin2int(port_link_number);
constant retry_buffer_last_active_address_int	:	integer	:=	bin2int(retry_buffer_last_active_address);
constant revision_id_int	:	integer	:=	bin2int(revision_id);
constant rp_bug_fix_pri_sec_stat_reg_int	:	integer	:=	bin2int(rp_bug_fix_pri_sec_stat_reg);
constant rpltim_base_int	:	integer	:=	bin2int(rpltim_base);
constant rstctrl_1ms_count_fref_clk_int	:	integer	:=	bin2int(rstctrl_1ms_count_fref_clk);
constant rstctrl_1us_count_fref_clk_int	:	integer	:=	bin2int(rstctrl_1us_count_fref_clk);
constant rstctrl_timer_a_int	:	integer	:=	bin2int(rstctrl_timer_a);
constant rstctrl_timer_b_int	:	integer	:=	bin2int(rstctrl_timer_b);
constant rstctrl_timer_c_int	:	integer	:=	bin2int(rstctrl_timer_c);
constant rstctrl_timer_d_int	:	integer	:=	bin2int(rstctrl_timer_d);
constant rstctrl_timer_e_int	:	integer	:=	bin2int(rstctrl_timer_e);
constant rstctrl_timer_f_int	:	integer	:=	bin2int(rstctrl_timer_f);
constant rstctrl_timer_g_int	:	integer	:=	bin2int(rstctrl_timer_g);
constant rstctrl_timer_h_int	:	integer	:=	bin2int(rstctrl_timer_h);
constant rstctrl_timer_i_int	:	integer	:=	bin2int(rstctrl_timer_i);
constant rstctrl_timer_j_int	:	integer	:=	bin2int(rstctrl_timer_j);
constant rx_buffer_fc_protect_int	:	integer	:=	bin2int(rx_buffer_fc_protect);
constant rx_buffer_protect_int	:	integer	:=	bin2int(rx_buffer_protect);
constant rx_cdc_almost_empty_int	:	integer	:=	bin2int(rx_cdc_almost_empty);
constant rx_cdc_almost_full_int	:	integer	:=	bin2int(rx_cdc_almost_full);
constant rx_l0s_count_idl_int	:	integer	:=	bin2int(rx_l0s_count_idl);
constant rx_ptr0_nonposted_dpram_max_int	:	integer	:=	bin2int(rx_ptr0_nonposted_dpram_max);
constant rx_ptr0_nonposted_dpram_min_int	:	integer	:=	bin2int(rx_ptr0_nonposted_dpram_min);
constant rx_ptr0_posted_dpram_max_int	:	integer	:=	bin2int(rx_ptr0_posted_dpram_max);
constant rx_ptr0_posted_dpram_min_int	:	integer	:=	bin2int(rx_ptr0_posted_dpram_min);
constant sameclock_nfts_count_int	:	integer	:=	bin2int(sameclock_nfts_count);
constant skp_os_gen3_count_int	:	integer	:=	bin2int(skp_os_gen3_count);
constant skp_os_schedule_count_int	:	integer	:=	bin2int(skp_os_schedule_count);
constant slot_number_int	:	integer	:=	bin2int(slot_number);
constant slot_power_limit_int	:	integer	:=	bin2int(slot_power_limit);
constant slot_power_scale_int	:	integer	:=	bin2int(slot_power_scale);
constant ssid_int	:	integer	:=	bin2int(ssid);
constant ssvid_int	:	integer	:=	bin2int(ssvid);
constant subsystem_device_id_int	:	integer	:=	bin2int(subsystem_device_id);
constant subsystem_vendor_id_int	:	integer	:=	bin2int(subsystem_vendor_id);
constant tx_cdc_almost_empty_int	:	integer	:=	bin2int(tx_cdc_almost_empty);
constant tx_cdc_almost_full_int	:	integer	:=	bin2int(tx_cdc_almost_full);
constant tx_swing_int	:	integer	:=	bin2int(tx_swing);
constant txdl_fair_arbiter_counter_int	:	integer	:=	bin2int(txdl_fair_arbiter_counter);
constant user_id_int	:	integer	:=	bin2int(user_id);
constant vc0_rx_flow_ctrl_compl_data_int	:	integer	:=	bin2int(vc0_rx_flow_ctrl_compl_data);
constant vc0_rx_flow_ctrl_compl_header_int	:	integer	:=	bin2int(vc0_rx_flow_ctrl_compl_header);
constant vc0_rx_flow_ctrl_nonposted_data_int	:	integer	:=	bin2int(vc0_rx_flow_ctrl_nonposted_data);
constant vc0_rx_flow_ctrl_nonposted_header_int	:	integer	:=	bin2int(vc0_rx_flow_ctrl_nonposted_header);
constant vc0_rx_flow_ctrl_posted_data_int	:	integer	:=	bin2int(vc0_rx_flow_ctrl_posted_data);
constant vc0_rx_flow_ctrl_posted_header_int	:	integer	:=	bin2int(vc0_rx_flow_ctrl_posted_header);
constant vendor_id_int	:	integer	:=	bin2int(vendor_id);
constant vsec_cap_int	:	integer	:=	bin2int(vsec_cap);
constant vsec_id_int	:	integer	:=	bin2int(vsec_id);



component	twentynm_hssi_gen3_x8_pcie_hip_encrypted
	generic (
		-- Architecture parameters
		acknack_base	:	integer	:=	0;
		acknack_set	:	string	:=	"false";
		advance_error_reporting	:	string	:=	"disable";
		app_interface_width	:	string	:=	"avst_64bit";
		arb_upfc_30us_counter	:	integer	:=	0;
		arb_upfc_30us_en	:	string	:=	"enable";
		aspm_config_management	:	string	:=	"true";
		aspm_patch_disable	:	string	:=	"enable_both";
		ast_width_rx	:	string	:=	"rx_64";
		ast_width_tx	:	string	:=	"tx_64";
		atomic_malformed	:	string	:=	"false";
		atomic_op_completer_32bit	:	string	:=	"false";
		atomic_op_completer_64bit	:	string	:=	"false";
		atomic_op_routing	:	string	:=	"false";
		auto_msg_drop_enable	:	string	:=	"false";
		avmm_cvp_inter_sel_csr_ctrl	:	string	:=	"disable";
		avmm_dprio_broadcast_en_csr_ctrl	:	string	:=	"disable";
		avmm_force_inter_sel_csr_ctrl	:	string	:=	"disable";
		avmm_power_iso_en_csr_ctrl	:	string	:=	"disable";
		bar0_size_mask	:	integer	:=	268435455;
		bar0_type	:	string	:=	"bar0_64bit_prefetch_mem";
		bar1_size_mask	:	integer	:=	0;
		bar1_type	:	string	:=	"bar1_disable";
		bar2_size_mask	:	integer	:=	0;
		bar2_type	:	string	:=	"bar2_disable";
		bar3_size_mask	:	integer	:=	0;
		bar3_type	:	string	:=	"bar3_disable";
		bar4_size_mask	:	integer	:=	0;
		bar4_type	:	string	:=	"bar4_disable";
		bar5_size_mask	:	integer	:=	0;
		bar5_type	:	string	:=	"bar5_disable";
		base_counter_sel	:	string	:=	"count_clk_62p5";
		bist_memory_settings	:	string	:=	"000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		bridge_port_ssid_support	:	string	:=	"false";
		bridge_port_vga_enable	:	string	:=	"false";
		bypass_cdc	:	string	:=	"false";
		bypass_clk_switch	:	string	:=	"false";
		bypass_tl	:	string	:=	"false";
		capab_rate_rxcfg_en	:	string	:=	"disable";
		cas_completer_128bit	:	string	:=	"false";
		cdc_clk_relation	:	string	:=	"plesiochronous";
		cdc_dummy_insert_limit	:	integer	:=	11;
		cfg_parchk_ena	:	string	:=	"disable";
		cfgbp_req_recov_disable	:	string	:=	"false";
		class_code	:	integer	:=	16711680;
		clock_pwr_management	:	string	:=	"false";
		completion_timeout	:	string	:=	"abcd";
		core_clk_divider	:	string	:=	"div_1";
		core_clk_freq_mhz	:	string	:=	"core_clk_250mhz";
		core_clk_out_sel	:	string	:=	"core_clk_out_div_1";
		core_clk_sel	:	string	:=	"pld_clk";
		core_clk_source	:	string	:=	"pll_fixed_clk";
		cseb_bar_match_checking	:	string	:=	"enable";
		cseb_config_bypass	:	string	:=	"disable";
		cseb_cpl_status_during_cvp	:	string	:=	"completer_abort";
		cseb_cpl_tag_checking	:	string	:=	"enable";
		cseb_disable_auto_crs	:	string	:=	"false";
		cseb_extend_pci	:	string	:=	"false";
		cseb_extend_pcie	:	string	:=	"false";
		cseb_min_error_checking	:	string	:=	"false";
		cseb_route_to_avl_rx_st	:	string	:=	"cseb";
		cseb_temp_busy_crs	:	string	:=	"completer_abort_tmp_busy";
		cvp_clk_reset	:	string	:=	"false";
		cvp_data_compressed	:	string	:=	"false";
		cvp_data_encrypted	:	string	:=	"false";
		cvp_enable	:	string	:=	"cvp_dis";
		cvp_mode_reset	:	string	:=	"false";
		cvp_rate_sel	:	string	:=	"full_rate";
		d0_pme	:	string	:=	"false";
		d1_pme	:	string	:=	"false";
		d1_support	:	string	:=	"false";
		d2_pme	:	string	:=	"false";
		d2_support	:	string	:=	"false";
		d3_cold_pme	:	string	:=	"false";
		d3_hot_pme	:	string	:=	"false";
		data_pack_rx	:	string	:=	"disable";
		deemphasis_enable	:	string	:=	"false";
		deskew_comma	:	string	:=	"skp_eieos_deskw";
		device_id	:	integer	:=	57345;
		device_number	:	integer	:=	0;
		device_specific_init	:	string	:=	"false";
		dft_clock_obsrv_en	:	string	:=	"disable";
		dft_clock_obsrv_sel	:	string	:=	"dft_pclk";
		diffclock_nfts_count	:	integer	:=	0;
		dis_cplovf	:	string	:=	"disable";
		dis_paritychk	:	string	:=	"enable";
		disable_link_x2_support	:	string	:=	"false";
		disable_snoop_packet	:	string	:=	"false";
		dl_tx_check_parity_edb	:	string	:=	"disable";
		dll_active_report_support	:	string	:=	"false";
		early_dl_up	:	string	:=	"true";
		eco_fb332688_dis	:	string	:=	"true";
		ecrc_check_capable	:	string	:=	"true";
		ecrc_gen_capable	:	string	:=	"true";
		egress_block_err_report_ena	:	string	:=	"false";
		ei_delay_powerdown_count	:	integer	:=	10;
		eie_before_nfts_count	:	integer	:=	4;
		electromech_interlock	:	string	:=	"false";
		en_ieiupdatefc	:	string	:=	"false";
		en_lane_errchk	:	string	:=	"false";
		en_phystatus_dly	:	string	:=	"false";
		ena_ido_cpl	:	string	:=	"false";
		ena_ido_req	:	string	:=	"false";
		enable_adapter_half_rate_mode	:	string	:=	"false";
		enable_ch01_pclk_out	:	string	:=	"pclk_ch0";
		enable_ch0_pclk_out	:	string	:=	"pclk_ch01";
		enable_completion_timeout_disable	:	string	:=	"true";
		enable_directed_spd_chng	:	string	:=	"false";
		enable_function_msix_support	:	string	:=	"true";
		enable_l0s_aspm	:	string	:=	"false";
		enable_l1_aspm	:	string	:=	"false";
		enable_rx_buffer_checking	:	string	:=	"false";
		enable_rx_reordering	:	string	:=	"true";
		enable_slot_register	:	string	:=	"false";
		endpoint_l0_latency	:	integer	:=	0;
		endpoint_l1_latency	:	integer	:=	0;
		eql_rq_int_en_number	:	integer	:=	0;
		errmgt_fcpe_patch_dis	:	string	:=	"enable";
		errmgt_fep_patch_dis	:	string	:=	"enable";
		expansion_base_address_register	:	string	:=	"00000000000000000000000000000000";
		extend_tag_field	:	string	:=	"false";
		extended_format_field	:	string	:=	"true";
		extended_tag_reset	:	string	:=	"false";
		fc_init_timer	:	integer	:=	1024;
		flow_control_timeout_count	:	integer	:=	200;
		flow_control_update_count	:	integer	:=	30;
		flr_capability	:	string	:=	"true";
		force_dis_to_det	:	string	:=	"false";
		force_gen1_dis	:	string	:=	"false";
		force_tx_coeff_preset_lpbk	:	string	:=	"false";
		frame_err_patch_dis	:	string	:=	"enable";
		func_mode	:	string	:=	"disable";
		g3_bypass_equlz	:	string	:=	"false";
		g3_coeff_done_tmout	:	string	:=	"enable";
		g3_deskew_char	:	string	:=	"default_sdsos";
		g3_dis_be_frm_err	:	string	:=	"false";
		g3_dn_rx_hint_eqlz_0	:	integer	:=	0;
		g3_dn_rx_hint_eqlz_1	:	integer	:=	0;
		g3_dn_rx_hint_eqlz_2	:	integer	:=	0;
		g3_dn_rx_hint_eqlz_3	:	integer	:=	0;
		g3_dn_rx_hint_eqlz_4	:	integer	:=	0;
		g3_dn_rx_hint_eqlz_5	:	integer	:=	0;
		g3_dn_rx_hint_eqlz_6	:	integer	:=	0;
		g3_dn_rx_hint_eqlz_7	:	integer	:=	0;
		g3_dn_tx_preset_eqlz_0	:	integer	:=	0;
		g3_dn_tx_preset_eqlz_1	:	integer	:=	0;
		g3_dn_tx_preset_eqlz_2	:	integer	:=	0;
		g3_dn_tx_preset_eqlz_3	:	integer	:=	0;
		g3_dn_tx_preset_eqlz_4	:	integer	:=	0;
		g3_dn_tx_preset_eqlz_5	:	integer	:=	0;
		g3_dn_tx_preset_eqlz_6	:	integer	:=	0;
		g3_dn_tx_preset_eqlz_7	:	integer	:=	0;
		g3_force_ber_max	:	string	:=	"false";
		g3_force_ber_min	:	string	:=	"false";
		g3_lnk_trn_rx_ts	:	string	:=	"false";
		g3_ltssm_eq_dbg	:	string	:=	"false";
		g3_ltssm_rec_dbg	:	string	:=	"false";
		g3_pause_ltssm_rec_en	:	string	:=	"disable";
		g3_quiesce_guarant	:	string	:=	"false";
		g3_redo_equlz_dis	:	string	:=	"false";
		g3_redo_equlz_en	:	string	:=	"false";
		g3_up_rx_hint_eqlz_0	:	integer	:=	0;
		g3_up_rx_hint_eqlz_1	:	integer	:=	0;
		g3_up_rx_hint_eqlz_2	:	integer	:=	0;
		g3_up_rx_hint_eqlz_3	:	integer	:=	0;
		g3_up_rx_hint_eqlz_4	:	integer	:=	0;
		g3_up_rx_hint_eqlz_5	:	integer	:=	0;
		g3_up_rx_hint_eqlz_6	:	integer	:=	0;
		g3_up_rx_hint_eqlz_7	:	integer	:=	0;
		g3_up_tx_preset_eqlz_0	:	integer	:=	0;
		g3_up_tx_preset_eqlz_1	:	integer	:=	0;
		g3_up_tx_preset_eqlz_2	:	integer	:=	0;
		g3_up_tx_preset_eqlz_3	:	integer	:=	0;
		g3_up_tx_preset_eqlz_4	:	integer	:=	0;
		g3_up_tx_preset_eqlz_5	:	integer	:=	0;
		g3_up_tx_preset_eqlz_6	:	integer	:=	0;
		g3_up_tx_preset_eqlz_7	:	integer	:=	0;
		gen123_lane_rate_mode	:	string	:=	"gen1_rate";
		gen2_diffclock_nfts_count	:	integer	:=	255;
		gen2_pma_pll_usage	:	string	:=	"not_applicaple";
		gen2_sameclock_nfts_count	:	integer	:=	255;
		gen3_coeff_1	:	integer	:=	4;
		gen3_coeff_10	:	integer	:=	7;
		gen3_coeff_10_ber_meas	:	integer	:=	2;
		gen3_coeff_10_nxtber_less	:	integer	:=	15;
		gen3_coeff_10_nxtber_more	:	integer	:=	10;
		gen3_coeff_10_preset_hint	:	integer	:=	3;
		gen3_coeff_10_reqber	:	integer	:=	8;
		gen3_coeff_10_sel	:	string	:=	"preset_10";
		gen3_coeff_11	:	integer	:=	7;
		gen3_coeff_11_ber_meas	:	integer	:=	2;
		gen3_coeff_11_nxtber_less	:	integer	:=	15;
		gen3_coeff_11_nxtber_more	:	integer	:=	15;
		gen3_coeff_11_preset_hint	:	integer	:=	4;
		gen3_coeff_11_reqber	:	integer	:=	8;
		gen3_coeff_11_sel	:	string	:=	"preset_11";
		gen3_coeff_12	:	integer	:=	7;
		gen3_coeff_12_ber_meas	:	integer	:=	2;
		gen3_coeff_12_nxtber_less	:	integer	:=	15;
		gen3_coeff_12_nxtber_more	:	integer	:=	15;
		gen3_coeff_12_preset_hint	:	integer	:=	2;
		gen3_coeff_12_reqber	:	integer	:=	8;
		gen3_coeff_12_sel	:	string	:=	"preset_12";
		gen3_coeff_13	:	integer	:=	4;
		gen3_coeff_13_ber_meas	:	integer	:=	2;
		gen3_coeff_13_nxtber_less	:	integer	:=	13;
		gen3_coeff_13_nxtber_more	:	integer	:=	1;
		gen3_coeff_13_preset_hint	:	integer	:=	4;
		gen3_coeff_13_reqber	:	integer	:=	8;
		gen3_coeff_13_sel	:	string	:=	"preset_13";
		gen3_coeff_14	:	integer	:=	4;
		gen3_coeff_14_ber_meas	:	integer	:=	2;
		gen3_coeff_14_nxtber_less	:	integer	:=	15;
		gen3_coeff_14_nxtber_more	:	integer	:=	2;
		gen3_coeff_14_preset_hint	:	integer	:=	0;
		gen3_coeff_14_reqber	:	integer	:=	8;
		gen3_coeff_14_sel	:	string	:=	"preset_14";
		gen3_coeff_15	:	integer	:=	0;
		gen3_coeff_15_ber_meas	:	integer	:=	2;
		gen3_coeff_15_nxtber_less	:	integer	:=	0;
		gen3_coeff_15_nxtber_more	:	integer	:=	0;
		gen3_coeff_15_preset_hint	:	integer	:=	0;
		gen3_coeff_15_reqber	:	integer	:=	0;
		gen3_coeff_15_sel	:	string	:=	"coeff_15";
		gen3_coeff_16	:	integer	:=	0;
		gen3_coeff_16_ber_meas	:	integer	:=	0;
		gen3_coeff_16_nxtber_less	:	integer	:=	0;
		gen3_coeff_16_nxtber_more	:	integer	:=	0;
		gen3_coeff_16_preset_hint	:	integer	:=	0;
		gen3_coeff_16_reqber	:	integer	:=	0;
		gen3_coeff_16_sel	:	string	:=	"coeff_16";
		gen3_coeff_17	:	integer	:=	0;
		gen3_coeff_17_ber_meas	:	integer	:=	0;
		gen3_coeff_17_nxtber_less	:	integer	:=	0;
		gen3_coeff_17_nxtber_more	:	integer	:=	0;
		gen3_coeff_17_preset_hint	:	integer	:=	0;
		gen3_coeff_17_reqber	:	integer	:=	0;
		gen3_coeff_17_sel	:	string	:=	"coeff_17";
		gen3_coeff_18	:	integer	:=	0;
		gen3_coeff_18_ber_meas	:	integer	:=	0;
		gen3_coeff_18_nxtber_less	:	integer	:=	0;
		gen3_coeff_18_nxtber_more	:	integer	:=	0;
		gen3_coeff_18_preset_hint	:	integer	:=	0;
		gen3_coeff_18_reqber	:	integer	:=	0;
		gen3_coeff_18_sel	:	string	:=	"coeff_18";
		gen3_coeff_19	:	integer	:=	0;
		gen3_coeff_19_ber_meas	:	integer	:=	0;
		gen3_coeff_19_nxtber_less	:	integer	:=	0;
		gen3_coeff_19_nxtber_more	:	integer	:=	0;
		gen3_coeff_19_preset_hint	:	integer	:=	0;
		gen3_coeff_19_reqber	:	integer	:=	0;
		gen3_coeff_19_sel	:	string	:=	"coeff_19";
		gen3_coeff_1_ber_meas	:	integer	:=	2;
		gen3_coeff_1_nxtber_less	:	integer	:=	12;
		gen3_coeff_1_nxtber_more	:	integer	:=	6;
		gen3_coeff_1_preset_hint	:	integer	:=	2;
		gen3_coeff_1_reqber	:	integer	:=	8;
		gen3_coeff_1_sel	:	string	:=	"preset_1";
		gen3_coeff_2	:	integer	:=	1;
		gen3_coeff_20	:	integer	:=	0;
		gen3_coeff_20_ber_meas	:	integer	:=	0;
		gen3_coeff_20_nxtber_less	:	integer	:=	0;
		gen3_coeff_20_nxtber_more	:	integer	:=	0;
		gen3_coeff_20_preset_hint	:	integer	:=	0;
		gen3_coeff_20_reqber	:	integer	:=	0;
		gen3_coeff_20_sel	:	string	:=	"coeff_20";
		gen3_coeff_21	:	integer	:=	0;
		gen3_coeff_21_ber_meas	:	integer	:=	0;
		gen3_coeff_21_nxtber_less	:	integer	:=	0;
		gen3_coeff_21_nxtber_more	:	integer	:=	0;
		gen3_coeff_21_preset_hint	:	integer	:=	0;
		gen3_coeff_21_reqber	:	integer	:=	0;
		gen3_coeff_21_sel	:	string	:=	"coeff_21";
		gen3_coeff_22	:	integer	:=	0;
		gen3_coeff_22_ber_meas	:	integer	:=	0;
		gen3_coeff_22_nxtber_less	:	integer	:=	0;
		gen3_coeff_22_nxtber_more	:	integer	:=	0;
		gen3_coeff_22_preset_hint	:	integer	:=	0;
		gen3_coeff_22_reqber	:	integer	:=	0;
		gen3_coeff_22_sel	:	string	:=	"coeff_22";
		gen3_coeff_23	:	integer	:=	0;
		gen3_coeff_23_ber_meas	:	integer	:=	0;
		gen3_coeff_23_nxtber_less	:	integer	:=	0;
		gen3_coeff_23_nxtber_more	:	integer	:=	0;
		gen3_coeff_23_preset_hint	:	integer	:=	0;
		gen3_coeff_23_reqber	:	integer	:=	0;
		gen3_coeff_23_sel	:	string	:=	"coeff_23";
		gen3_coeff_24	:	integer	:=	0;
		gen3_coeff_24_ber_meas	:	integer	:=	0;
		gen3_coeff_24_nxtber_less	:	integer	:=	0;
		gen3_coeff_24_nxtber_more	:	integer	:=	0;
		gen3_coeff_24_preset_hint	:	integer	:=	0;
		gen3_coeff_24_reqber	:	integer	:=	0;
		gen3_coeff_24_sel	:	string	:=	"coeff_24";
		gen3_coeff_2_ber_meas	:	integer	:=	2;
		gen3_coeff_2_nxtber_less	:	integer	:=	2;
		gen3_coeff_2_nxtber_more	:	integer	:=	4;
		gen3_coeff_2_preset_hint	:	integer	:=	4;
		gen3_coeff_2_reqber	:	integer	:=	8;
		gen3_coeff_2_sel	:	string	:=	"preset_2";
		gen3_coeff_3	:	integer	:=	1;
		gen3_coeff_3_ber_meas	:	integer	:=	2;
		gen3_coeff_3_nxtber_less	:	integer	:=	15;
		gen3_coeff_3_nxtber_more	:	integer	:=	3;
		gen3_coeff_3_preset_hint	:	integer	:=	0;
		gen3_coeff_3_reqber	:	integer	:=	8;
		gen3_coeff_3_sel	:	string	:=	"preset_3";
		gen3_coeff_4	:	integer	:=	0;
		gen3_coeff_4_ber_meas	:	integer	:=	2;
		gen3_coeff_4_nxtber_less	:	integer	:=	15;
		gen3_coeff_4_nxtber_more	:	integer	:=	4;
		gen3_coeff_4_preset_hint	:	integer	:=	0;
		gen3_coeff_4_reqber	:	integer	:=	8;
		gen3_coeff_4_sel	:	string	:=	"preset_4";
		gen3_coeff_5	:	integer	:=	0;
		gen3_coeff_5_ber_meas	:	integer	:=	2;
		gen3_coeff_5_nxtber_less	:	integer	:=	15;
		gen3_coeff_5_nxtber_more	:	integer	:=	5;
		gen3_coeff_5_preset_hint	:	integer	:=	4;
		gen3_coeff_5_reqber	:	integer	:=	8;
		gen3_coeff_5_sel	:	string	:=	"preset_5";
		gen3_coeff_6	:	integer	:=	7;
		gen3_coeff_6_ber_meas	:	integer	:=	2;
		gen3_coeff_6_nxtber_less	:	integer	:=	15;
		gen3_coeff_6_nxtber_more	:	integer	:=	15;
		gen3_coeff_6_preset_hint	:	integer	:=	4;
		gen3_coeff_6_reqber	:	integer	:=	8;
		gen3_coeff_6_sel	:	string	:=	"preset_6";
		gen3_coeff_7	:	integer	:=	1;
		gen3_coeff_7_ber_meas	:	integer	:=	2;
		gen3_coeff_7_nxtber_less	:	integer	:=	1;
		gen3_coeff_7_nxtber_more	:	integer	:=	7;
		gen3_coeff_7_preset_hint	:	integer	:=	2;
		gen3_coeff_7_reqber	:	integer	:=	8;
		gen3_coeff_7_sel	:	string	:=	"preset_7";
		gen3_coeff_8	:	integer	:=	0;
		gen3_coeff_8_ber_meas	:	integer	:=	2;
		gen3_coeff_8_nxtber_less	:	integer	:=	4;
		gen3_coeff_8_nxtber_more	:	integer	:=	8;
		gen3_coeff_8_preset_hint	:	integer	:=	2;
		gen3_coeff_8_reqber	:	integer	:=	8;
		gen3_coeff_8_sel	:	string	:=	"preset_8";
		gen3_coeff_9	:	integer	:=	0;
		gen3_coeff_9_ber_meas	:	integer	:=	2;
		gen3_coeff_9_nxtber_less	:	integer	:=	11;
		gen3_coeff_9_nxtber_more	:	integer	:=	9;
		gen3_coeff_9_preset_hint	:	integer	:=	3;
		gen3_coeff_9_reqber	:	integer	:=	8;
		gen3_coeff_9_sel	:	string	:=	"preset_9";
		gen3_coeff_delay_count	:	integer	:=	125;
		gen3_coeff_errchk	:	string	:=	"enable";
		gen3_dcbal_en	:	string	:=	"true";
		gen3_diffclock_nfts_count	:	integer	:=	128;
		gen3_force_local_coeff	:	string	:=	"false";
		gen3_full_swing	:	integer	:=	63;
		gen3_half_swing	:	string	:=	"false";
		gen3_low_freq	:	integer	:=	1;
		gen3_paritychk	:	string	:=	"enable";
		gen3_pl_framing_err_dis	:	string	:=	"enable";
		gen3_preset_coeff_1	:	integer	:=	3402;
		gen3_preset_coeff_10	:	integer	:=	48384;
		gen3_preset_coeff_11	:	integer	:=	124992;
		gen3_preset_coeff_2	:	integer	:=	3339;
		gen3_preset_coeff_3	:	integer	:=	3213;
		gen3_preset_coeff_4	:	integer	:=	3528;
		gen3_preset_coeff_5	:	integer	:=	4032;
		gen3_preset_coeff_6	:	integer	:=	28224;
		gen3_preset_coeff_7	:	integer	:=	36288;
		gen3_preset_coeff_8	:	integer	:=	27405;
		gen3_preset_coeff_9	:	integer	:=	35784;
		gen3_reset_eieos_cnt_bit	:	string	:=	"false";
		gen3_rxfreqlock_counter	:	integer	:=	0;
		gen3_sameclock_nfts_count	:	integer	:=	128;
		gen3_scrdscr_bypass	:	string	:=	"false";
		gen3_skip_ph2_ph3	:	string	:=	"false";
		hard_reset_bypass	:	string	:=	"false";
		hard_rst_sig_chnl_en	:	string	:=	"disable_hrc_sig";
		hard_rst_tx_pll_rst_chnl_en	:	string	:=	"disable_hrc_txpll_rst";
		hip_ac_pwr_clk_freq_in_hz	:	integer	:=	0;
		hip_ac_pwr_uw_per_mhz	:	integer	:=	0;
		hip_base_address	:	integer	:=	0;
		hip_clock_dis	:	string	:=	"enable_hip_clk";
		hip_hard_reset	:	string	:=	"enable";
		hip_pcs_sig_chnl_en	:	string	:=	"disable_hip_pcs_sig";
		hot_plug_support	:	integer	:=	0;
		hrc_chnl_txpll_master_cgb_rst_select	:	string	:=	"disable_master_cgb_sel";
		hrdrstctrl_en	:	string	:=	"hrdrstctrl_dis";
		iei_enable_settings	:	string	:=	"gen3gen2_infei_infsd_gen1_infei_sd";
		indicator	:	integer	:=	7;
		intel_id_access	:	string	:=	"false";
		interrupt_pin	:	string	:=	"inta";
		io_window_addr_width	:	string	:=	"window_32_bit";
		jtag_id	:	string	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		ko_compl_data	:	integer	:=	0;
		ko_compl_header	:	integer	:=	0;
		l01_entry_latency	:	integer	:=	31;
		l0_exit_latency_diffclock	:	integer	:=	6;
		l0_exit_latency_sameclock	:	integer	:=	6;
		l0s_adj_rply_timer_dis	:	string	:=	"enable";
		l1_exit_latency_diffclock	:	integer	:=	0;
		l1_exit_latency_sameclock	:	integer	:=	0;
		l2_async_logic	:	string	:=	"enable";
		lane_mask	:	string	:=	"ln_mask_x4";
		lane_rate	:	string	:=	"gen1";
		link_width	:	string	:=	"x1";
		lmi_hold_off_cfg_timer_en	:	string	:=	"disable";
		low_priority_vc	:	string	:=	"single_vc_low_pr";
		ltr_mechanism	:	string	:=	"false";
		ltssm_1ms_timeout	:	string	:=	"disable";
		ltssm_freqlocked_check	:	string	:=	"disable";
		malformed_tlp_truncate_en	:	string	:=	"disable";
		max_link_width	:	string	:=	"x4_link_width";
		max_payload_size	:	string	:=	"payload_512";
		maximum_current	:	integer	:=	0;
		millisecond_cycle_count	:	integer	:=	0;
		msi_64bit_addressing_capable	:	string	:=	"true";
		msi_masking_capable	:	string	:=	"false";
		msi_multi_message_capable	:	string	:=	"count_4";
		msi_support	:	string	:=	"true";
		msix_pba_bir	:	integer	:=	0;
		msix_pba_offset	:	integer	:=	0;
		msix_table_bir	:	integer	:=	0;
		msix_table_offset	:	integer	:=	0;
		msix_table_size	:	integer	:=	0;
		national_inst_thru_enhance	:	string	:=	"true";
		no_command_completed	:	string	:=	"true";
		no_soft_reset	:	string	:=	"false";
		not_use_k_gbl_bits	:	string	:=	"not_used_k_gbl";
		operating_voltage	:	string	:=	"standard";
		pcie_base_spec	:	string	:=	"pcie_2p1";
		pcie_mode	:	string	:=	"shared_mode";
		pcie_spec_1p0_compliance	:	string	:=	"spec_1p1";
		pcie_spec_version	:	string	:=	"v2";
		pclk_out_sel	:	string	:=	"pclk";
		pld_in_use_reg	:	string	:=	"false";
		pm_latency_patch_dis	:	string	:=	"enable";
		pm_txdl_patch_dis	:	string	:=	"enable";
		pme_clock	:	string	:=	"false";
		port_link_number	:	integer	:=	1;
		port_type	:	string	:=	"native_ep";
		powerdown_mode	:	string	:=	"powerup";
		prefetchable_mem_window_addr_width	:	string	:=	"prefetch_32";
		r2c_mask_easy	:	string	:=	"false";
		r2c_mask_enable	:	string	:=	"false";
		rec_frqlk_mon_en	:	string	:=	"disable";
		register_pipe_signals	:	string	:=	"true";
		retry_buffer_last_active_address	:	integer	:=	1023;
		retry_buffer_memory_settings	:	string	:=	"000000000000000000000000000000000000";
		retry_ecc_corr_mask_dis	:	string	:=	"enable";
		revision_id	:	integer	:=	1;
		role_based_error_reporting	:	string	:=	"false";
		rp_bug_fix_pri_sec_stat_reg	:	integer	:=	127;
		rpltim_base	:	integer	:=	0;
		rpltim_set	:	string	:=	"false";
		rstctl_ltssm_dis	:	string	:=	"false";
		rstctrl_1ms_count_fref_clk	:	integer	:=	62500;
		rstctrl_1us_count_fref_clk	:	integer	:=	63;
		rstctrl_altpe3_crst_n_inv	:	string	:=	"false";
		rstctrl_altpe3_rst_n_inv	:	string	:=	"false";
		rstctrl_altpe3_srst_n_inv	:	string	:=	"false";
		rstctrl_chnl_cal_done_select	:	string	:=	"not_active_chnl_cal_done";
		rstctrl_debug_en	:	string	:=	"false";
		rstctrl_force_inactive_rst	:	string	:=	"false";
		rstctrl_fref_clk_select	:	string	:=	"ch0_sel";
		rstctrl_hard_block_enable	:	string	:=	"hard_rst_ctl";
		rstctrl_hip_ep	:	string	:=	"hip_ep";
		rstctrl_mask_tx_pll_lock_select	:	string	:=	"not_active_mask_tx_pll_lock";
		rstctrl_perst_enable	:	string	:=	"level";
		rstctrl_perstn_select	:	string	:=	"perstn_pin";
		rstctrl_pld_clr	:	string	:=	"false";
		rstctrl_pll_cal_done_select	:	string	:=	"not_active_pll_cal_done";
		rstctrl_rx_pcs_rst_n_inv	:	string	:=	"false";
		rstctrl_rx_pcs_rst_n_select	:	string	:=	"not_active_rx_pcs_rst";
		rstctrl_rx_pll_freq_lock_select	:	string	:=	"not_active_rx_pll_f_lock";
		rstctrl_rx_pll_lock_select	:	string	:=	"not_active_rx_pll_lock";
		rstctrl_rx_pma_rstb_inv	:	string	:=	"false";
		rstctrl_rx_pma_rstb_select	:	string	:=	"not_active_rx_pma_rstb";
		rstctrl_timer_a	:	integer	:=	10;
		rstctrl_timer_a_type	:	string	:=	"a_timer_milli_secs";
		rstctrl_timer_b	:	integer	:=	10;
		rstctrl_timer_b_type	:	string	:=	"b_timer_milli_secs";
		rstctrl_timer_c	:	integer	:=	10;
		rstctrl_timer_c_type	:	string	:=	"c_timer_milli_secs";
		rstctrl_timer_d	:	integer	:=	20;
		rstctrl_timer_d_type	:	string	:=	"d_timer_milli_secs";
		rstctrl_timer_e	:	integer	:=	1;
		rstctrl_timer_e_type	:	string	:=	"e_timer_milli_secs";
		rstctrl_timer_f	:	integer	:=	10;
		rstctrl_timer_f_type	:	string	:=	"f_timer_milli_secs";
		rstctrl_timer_g	:	integer	:=	10;
		rstctrl_timer_g_type	:	string	:=	"g_timer_milli_secs";
		rstctrl_timer_h	:	integer	:=	4;
		rstctrl_timer_h_type	:	string	:=	"h_timer_milli_secs";
		rstctrl_timer_i	:	integer	:=	20;
		rstctrl_timer_i_type	:	string	:=	"i_timer_milli_secs";
		rstctrl_timer_j	:	integer	:=	20;
		rstctrl_timer_j_type	:	string	:=	"j_timer_milli_secs";
		rstctrl_tx_lcff_pll_lock_select	:	string	:=	"not_active_lcff_pll_lock";
		rstctrl_tx_lcff_pll_rstb_select	:	string	:=	"not_active_lcff_pll_rstb";
		rstctrl_tx_pcs_rst_n_inv	:	string	:=	"false";
		rstctrl_tx_pcs_rst_n_select	:	string	:=	"not_active_tx_pcs_rst";
		rstctrl_tx_pma_rstb_inv	:	string	:=	"false";
		rstctrl_tx_pma_syncp_inv	:	string	:=	"false";
		rstctrl_tx_pma_syncp_select	:	string	:=	"not_active_tx_pma_syncp";
		rx_ast_parity	:	string	:=	"disable";
		rx_buffer_credit_alloc	:	string	:=	"balance";
		rx_buffer_fc_protect	:	integer	:=	68;
		rx_buffer_protect	:	integer	:=	68;
		rx_cdc_almost_empty	:	integer	:=	3;
		rx_cdc_almost_full	:	integer	:=	12;
		rx_cred_ctl_param	:	string	:=	"disable";
		rx_ei_l0s	:	string	:=	"disable";
		rx_l0s_count_idl	:	integer	:=	0;
		rx_ptr0_nonposted_dpram_max	:	integer	:=	0;
		rx_ptr0_nonposted_dpram_min	:	integer	:=	0;
		rx_ptr0_posted_dpram_max	:	integer	:=	0;
		rx_ptr0_posted_dpram_min	:	integer	:=	0;
		rx_runt_patch_dis	:	string	:=	"enable";
		rx_sop_ctrl	:	string	:=	"rx_sop_boundary_64";
		rx_trunc_patch_dis	:	string	:=	"enable";
		rx_use_prst	:	string	:=	"false";
		rx_use_prst_ep	:	string	:=	"true";
		rxbuf_ecc_corr_mask_dis	:	string	:=	"enable";
		rxdl_bad_sop_eop_filter_dis	:	string	:=	"rxdlbug1_enable_both";
		rxdl_bad_tlp_patch_dis	:	string	:=	"rxdlbug2_enable_both";
		rxdl_lcrc_patch_dis	:	string	:=	"rxdlbug3_enable_both";
		sameclock_nfts_count	:	integer	:=	0;
		sel_enable_pcs_rx_fifo_err	:	string	:=	"disable_sel";
		silicon_rev	:	string	:=	"20nm5es";
		sim_mode	:	string	:=	"disable";
		simple_ro_fifo_control_en	:	string	:=	"disable";
		single_rx_detect	:	string	:=	"detect_all_lanes";
		skp_os_gen3_count	:	integer	:=	0;
		skp_os_schedule_count	:	integer	:=	0;
		slot_number	:	integer	:=	0;
		slot_power_limit	:	integer	:=	0;
		slot_power_scale	:	integer	:=	0;
		slotclk_cfg	:	string	:=	"static_slotclkcfgon";
		ssid	:	integer	:=	0;
		ssvid	:	integer	:=	0;
		subsystem_device_id	:	integer	:=	57345;
		subsystem_vendor_id	:	integer	:=	4466;
		sup_mode	:	string	:=	"user_mode";
		surprise_down_error_support	:	string	:=	"false";
		tl_cfg_div	:	string	:=	"cfg_clk_div_7";
		tl_tx_check_parity_msg	:	string	:=	"disable";
		tph_completer	:	string	:=	"false";
		tx_ast_parity	:	string	:=	"disable";
		tx_cdc_almost_empty	:	integer	:=	5;
		tx_cdc_almost_full	:	integer	:=	12;
		tx_sop_ctrl	:	string	:=	"boundary_64";
		tx_swing	:	integer	:=	0;
		txdl_fair_arbiter_counter	:	integer	:=	0;
		txdl_fair_arbiter_en	:	string	:=	"enable";
		txrate_adv	:	string	:=	"capability";
		uc_calibration_en	:	string	:=	"uc_calibration_dis";
		use_aer	:	string	:=	"false";
		use_crc_forwarding	:	string	:=	"false";
		user_id	:	integer	:=	0;
		vc0_clk_enable	:	string	:=	"true";
		vc0_rx_buffer_memory_settings	:	string	:=	"000000000000000000000000000000000000";
		vc0_rx_flow_ctrl_compl_data	:	integer	:=	448;
		vc0_rx_flow_ctrl_compl_header	:	integer	:=	112;
		vc0_rx_flow_ctrl_nonposted_data	:	integer	:=	0;
		vc0_rx_flow_ctrl_nonposted_header	:	integer	:=	54;
		vc0_rx_flow_ctrl_posted_data	:	integer	:=	360;
		vc0_rx_flow_ctrl_posted_header	:	integer	:=	50;
		vc1_clk_enable	:	string	:=	"false";
		vc_arbitration	:	string	:=	"single_vc_arb";
		vc_enable	:	string	:=	"single_vc";
		vendor_id	:	integer	:=	4466;
		vsec_cap	:	integer	:=	0;
		vsec_id	:	integer	:=	4466;
		wrong_device_id	:	string	:=	"disable"
	);
	port (
		-- Architecture ports
		aer_msi_num	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		app_int_err	:	in	std_logic_vector(1 downto 0)	:=	"00";
		app_inta_sts	:	in	std_logic	:=	'0';
		app_msi_num	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		app_msi_req	:	in	std_logic	:=	'0';
		app_msi_tc	:	in	std_logic_vector(2 downto 0)	:=	"000";
		atpg_los_en_n	:	in	std_logic	:=	'0';
		avmm_address	:	in	std_logic_vector(9 downto 0)	:=	"0000000000";
		avmm_byte_en	:	in	std_logic_vector(1 downto 0)	:=	"00";
		avmm_clk	:	in	std_logic	:=	'0';
		avmm_read	:	in	std_logic	:=	'0';
		avmm_rst_n	:	in	std_logic	:=	'0';
		avmm_write	:	in	std_logic	:=	'0';
		avmm_writedata	:	in	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		bist_scanen	:	in	std_logic	:=	'0';
		bist_scanin	:	in	std_logic	:=	'0';
		bisten_rcv_n	:	in	std_logic	:=	'0';
		bisten_rpl_n	:	in	std_logic	:=	'0';
		bistmode_n	:	in	std_logic	:=	'0';
		cfg_link2csr_pld	:	in	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		cfg_prmbus_pld	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		chnl_cal_done0	:	in	std_logic	:=	'0';
		chnl_cal_done1	:	in	std_logic	:=	'0';
		chnl_cal_done2	:	in	std_logic	:=	'0';
		chnl_cal_done3	:	in	std_logic	:=	'0';
		chnl_cal_done4	:	in	std_logic	:=	'0';
		chnl_cal_done5	:	in	std_logic	:=	'0';
		chnl_cal_done6	:	in	std_logic	:=	'0';
		chnl_cal_done7	:	in	std_logic	:=	'0';
		core_clk_in	:	in	std_logic	:=	'0';
		core_crst	:	in	std_logic	:=	'0';
		core_por	:	in	std_logic	:=	'0';
		core_rst	:	in	std_logic	:=	'0';
		core_srst	:	in	std_logic	:=	'0';
		cpl_err	:	in	std_logic_vector(6 downto 0)	:=	"0000000";
		cpl_pending	:	in	std_logic	:=	'0';
		cseb_rddata	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		cseb_rddata_parity	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		cseb_rdresponse	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		cseb_waitrequest	:	in	std_logic	:=	'0';
		cseb_wrresp_valid	:	in	std_logic	:=	'0';
		cseb_wrresponse	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		csr_cbdin	:	in	std_logic	:=	'0';
		csr_clk	:	in	std_logic	:=	'0';
		csr_din	:	in	std_logic	:=	'0';
		csr_en	:	in	std_logic	:=	'0';
		csr_enscan	:	in	std_logic	:=	'0';
		csr_entest	:	in	std_logic	:=	'0';
		csr_in	:	in	std_logic	:=	'0';
		csr_load_csr	:	in	std_logic	:=	'0';
		csr_pipe_in	:	in	std_logic	:=	'0';
		csr_seg	:	in	std_logic	:=	'0';
		csr_tcsrin	:	in	std_logic	:=	'0';
		csr_tverify	:	in	std_logic	:=	'0';
		cvp_config_done	:	in	std_logic	:=	'0';
		cvp_config_error	:	in	std_logic	:=	'0';
		cvp_config_ready	:	in	std_logic	:=	'0';
		cvp_en	:	in	std_logic	:=	'0';
		egress_blk_err	:	in	std_logic	:=	'0';
		entest	:	in	std_logic	:=	'0';
		flr_reset	:	in	std_logic	:=	'0';
		force_tx_eidle	:	in	std_logic	:=	'0';
		fref_clk0	:	in	std_logic	:=	'0';
		fref_clk1	:	in	std_logic	:=	'0';
		fref_clk2	:	in	std_logic	:=	'0';
		fref_clk3	:	in	std_logic	:=	'0';
		fref_clk4	:	in	std_logic	:=	'0';
		fref_clk5	:	in	std_logic	:=	'0';
		fref_clk6	:	in	std_logic	:=	'0';
		fref_clk7	:	in	std_logic	:=	'0';
		frzlogic	:	in	std_logic	:=	'0';
		frzreg	:	in	std_logic	:=	'0';
		hold_ltssm_rec	:	in	std_logic	:=	'0';
		hpg_ctrler	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		iocsrrdy_dly	:	in	std_logic	:=	'0';
		lmi_addr	:	in	std_logic_vector(11 downto 0)	:=	"000000000000";
		lmi_din	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		lmi_rden	:	in	std_logic	:=	'0';
		lmi_wren	:	in	std_logic	:=	'0';
		m10k_select	:	in	std_logic_vector(2 downto 0)	:=	"000";
		mask_tx_pll_lock0	:	in	std_logic	:=	'0';
		mask_tx_pll_lock1	:	in	std_logic	:=	'0';
		mask_tx_pll_lock2	:	in	std_logic	:=	'0';
		mask_tx_pll_lock3	:	in	std_logic	:=	'0';
		mask_tx_pll_lock4	:	in	std_logic	:=	'0';
		mask_tx_pll_lock5	:	in	std_logic	:=	'0';
		mask_tx_pll_lock6	:	in	std_logic	:=	'0';
		mask_tx_pll_lock7	:	in	std_logic	:=	'0';
		mem_hip_test_enable	:	in	std_logic	:=	'0';
		mem_regscanen_n	:	in	std_logic	:=	'0';
		mem_rscin_rcv_bot	:	in	std_logic	:=	'0';
		mem_rscin_rcv_top	:	in	std_logic	:=	'0';
		mem_rscin_rtry	:	in	std_logic	:=	'0';
		nfrzdrv	:	in	std_logic	:=	'0';
		npor	:	in	std_logic	:=	'0';
		pclk_central	:	in	std_logic	:=	'0';
		pclk_ch0	:	in	std_logic	:=	'0';
		pclk_ch1	:	in	std_logic	:=	'0';
		pex_msi_num	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		phy_rst	:	in	std_logic	:=	'0';
		phy_srst	:	in	std_logic	:=	'0';
		phystatus0	:	in	std_logic	:=	'0';
		phystatus1	:	in	std_logic	:=	'0';
		phystatus2	:	in	std_logic	:=	'0';
		phystatus3	:	in	std_logic	:=	'0';
		phystatus4	:	in	std_logic	:=	'0';
		phystatus5	:	in	std_logic	:=	'0';
		phystatus6	:	in	std_logic	:=	'0';
		phystatus7	:	in	std_logic	:=	'0';
		pin_perst_n	:	in	std_logic	:=	'0';
		pld_clk	:	in	std_logic	:=	'0';
		pld_clrhip_n	:	in	std_logic	:=	'0';
		pld_clrpcship_n	:	in	std_logic	:=	'0';
		pld_clrpmapcship_n	:	in	std_logic	:=	'0';
		pld_core_ready	:	in	std_logic	:=	'0';
		pld_gp_status	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		pld_perst_n	:	in	std_logic	:=	'0';
		pll_cal_done0	:	in	std_logic	:=	'0';
		pll_cal_done1	:	in	std_logic	:=	'0';
		pll_cal_done2	:	in	std_logic	:=	'0';
		pll_cal_done3	:	in	std_logic	:=	'0';
		pll_cal_done4	:	in	std_logic	:=	'0';
		pll_cal_done5	:	in	std_logic	:=	'0';
		pll_cal_done6	:	in	std_logic	:=	'0';
		pll_cal_done7	:	in	std_logic	:=	'0';
		pll_fixed_clk_central	:	in	std_logic	:=	'0';
		pll_fixed_clk_ch0	:	in	std_logic	:=	'0';
		pll_fixed_clk_ch1	:	in	std_logic	:=	'0';
		plniotri	:	in	std_logic	:=	'0';
		pm_auxpwr	:	in	std_logic	:=	'0';
		pm_data	:	in	std_logic_vector(9 downto 0)	:=	"0000000000";
		pm_event	:	in	std_logic	:=	'0';
		pm_exit_d0_ack	:	in	std_logic	:=	'0';
		pme_to_cr	:	in	std_logic	:=	'0';
		reserved_clk_in	:	in	std_logic	:=	'0';
		reserved_in	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		rx_cred_ctl	:	in	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		rx_pll_freq_lock0	:	in	std_logic	:=	'0';
		rx_pll_freq_lock1	:	in	std_logic	:=	'0';
		rx_pll_freq_lock2	:	in	std_logic	:=	'0';
		rx_pll_freq_lock3	:	in	std_logic	:=	'0';
		rx_pll_freq_lock4	:	in	std_logic	:=	'0';
		rx_pll_freq_lock5	:	in	std_logic	:=	'0';
		rx_pll_freq_lock6	:	in	std_logic	:=	'0';
		rx_pll_freq_lock7	:	in	std_logic	:=	'0';
		rx_pll_phase_lock0	:	in	std_logic	:=	'0';
		rx_pll_phase_lock1	:	in	std_logic	:=	'0';
		rx_pll_phase_lock2	:	in	std_logic	:=	'0';
		rx_pll_phase_lock3	:	in	std_logic	:=	'0';
		rx_pll_phase_lock4	:	in	std_logic	:=	'0';
		rx_pll_phase_lock5	:	in	std_logic	:=	'0';
		rx_pll_phase_lock6	:	in	std_logic	:=	'0';
		rx_pll_phase_lock7	:	in	std_logic	:=	'0';
		rx_st_mask	:	in	std_logic	:=	'0';
		rx_st_ready	:	in	std_logic	:=	'0';
		rxblkst0	:	in	std_logic	:=	'0';
		rxblkst1	:	in	std_logic	:=	'0';
		rxblkst2	:	in	std_logic	:=	'0';
		rxblkst3	:	in	std_logic	:=	'0';
		rxblkst4	:	in	std_logic	:=	'0';
		rxblkst5	:	in	std_logic	:=	'0';
		rxblkst6	:	in	std_logic	:=	'0';
		rxblkst7	:	in	std_logic	:=	'0';
		rxdata0	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata1	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata2	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata3	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata4	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata5	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata6	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata7	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdatak0	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak1	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak2	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak3	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak4	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak5	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak6	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak7	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdataskip0	:	in	std_logic	:=	'0';
		rxdataskip1	:	in	std_logic	:=	'0';
		rxdataskip2	:	in	std_logic	:=	'0';
		rxdataskip3	:	in	std_logic	:=	'0';
		rxdataskip4	:	in	std_logic	:=	'0';
		rxdataskip5	:	in	std_logic	:=	'0';
		rxdataskip6	:	in	std_logic	:=	'0';
		rxdataskip7	:	in	std_logic	:=	'0';
		rxelecidle0	:	in	std_logic	:=	'0';
		rxelecidle1	:	in	std_logic	:=	'0';
		rxelecidle2	:	in	std_logic	:=	'0';
		rxelecidle3	:	in	std_logic	:=	'0';
		rxelecidle4	:	in	std_logic	:=	'0';
		rxelecidle5	:	in	std_logic	:=	'0';
		rxelecidle6	:	in	std_logic	:=	'0';
		rxelecidle7	:	in	std_logic	:=	'0';
		rxfreqlocked0	:	in	std_logic	:=	'0';
		rxfreqlocked1	:	in	std_logic	:=	'0';
		rxfreqlocked2	:	in	std_logic	:=	'0';
		rxfreqlocked3	:	in	std_logic	:=	'0';
		rxfreqlocked4	:	in	std_logic	:=	'0';
		rxfreqlocked5	:	in	std_logic	:=	'0';
		rxfreqlocked6	:	in	std_logic	:=	'0';
		rxfreqlocked7	:	in	std_logic	:=	'0';
		rxstatus0	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus1	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus2	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus3	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus4	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus5	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus6	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus7	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxsynchd0	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd1	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd2	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd3	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd4	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd5	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd6	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd7	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxvalid0	:	in	std_logic	:=	'0';
		rxvalid1	:	in	std_logic	:=	'0';
		rxvalid2	:	in	std_logic	:=	'0';
		rxvalid3	:	in	std_logic	:=	'0';
		rxvalid4	:	in	std_logic	:=	'0';
		rxvalid5	:	in	std_logic	:=	'0';
		rxvalid6	:	in	std_logic	:=	'0';
		rxvalid7	:	in	std_logic	:=	'0';
		scan_mode_n	:	in	std_logic	:=	'0';
		scan_shift_n	:	in	std_logic	:=	'0';
		sw_ctmod	:	in	std_logic_vector(1 downto 0)	:=	"00";
		swdn_in	:	in	std_logic_vector(2 downto 0)	:=	"000";
		swup_in	:	in	std_logic_vector(6 downto 0)	:=	"0000000";
		test_in_1_hip	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		test_in_hip	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		test_pl_dbg_eqin	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		tx_cred_cons_select	:	in	std_logic	:=	'0';
		tx_cred_fc_sel	:	in	std_logic_vector(1 downto 0)	:=	"00";
		tx_lcff_pll_lock0	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock1	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock2	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock3	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock4	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock5	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock6	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock7	:	in	std_logic	:=	'0';
		tx_st_data	:	in	std_logic_vector(255 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		tx_st_empty	:	in	std_logic_vector(1 downto 0)	:=	"00";
		tx_st_eop	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		tx_st_err	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		tx_st_parity	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		tx_st_sop	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		tx_st_valid	:	in	std_logic	:=	'0';
		user_mode	:	in	std_logic	:=	'0';
		sta_hd_altpe3_hip_core_top_hd_altpe3_hip_core_u_clkmux_core_clk_cnt_reg_0_0_Q	:	out	std_logic	:=	'0';
		sta_hd_altpe3_hip_core_top_hd_altpe3_hip_core_u_clkmux_core_clk_cnt_reg_1_0_Q	:	out	std_logic	:=	'0';
		sta_hd_altpe3_hip_core_top_hd_altpe3_hip_core_u_clkmux_core_clk_cnt_reg_2_0_Q	:	out	std_logic	:=	'0';
		app_inta_ack	:	out	std_logic	:=	'0';
		app_msi_ack	:	out	std_logic	:=	'0';
		avmm_readdata	:	out	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		cfg_par_err	:	out	std_logic	:=	'0';
		core_clk_out	:	out	std_logic	:=	'0';
		cseb_addr	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		cseb_addr_parity	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		cseb_be	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		cseb_is_shadow	:	out	std_logic	:=	'0';
		cseb_rden	:	out	std_logic	:=	'0';
		cseb_wrdata	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		cseb_wrdata_parity	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		cseb_wren	:	out	std_logic	:=	'0';
		cseb_wrresp_req	:	out	std_logic	:=	'0';
		csr_dout	:	out	std_logic	:=	'0';
		csr_out	:	out	std_logic	:=	'0';
		csr_pipe_out	:	out	std_logic	:=	'0';
		current_coeff0	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff1	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff2	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff3	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff4	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff5	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff6	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff7	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_rxpreset0	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset1	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset2	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset3	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset4	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset5	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset6	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset7	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_speed	:	out	std_logic_vector(1 downto 0)	:=	"00";
		cvp_clk	:	out	std_logic	:=	'0';
		cvp_config	:	out	std_logic	:=	'0';
		cvp_data	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		cvp_full_config	:	out	std_logic	:=	'0';
		cvp_start_xfer	:	out	std_logic	:=	'0';
		dl_up	:	out	std_logic	:=	'0';
		dlup_exit	:	out	std_logic	:=	'0';
		eidle_infer_sel0	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel1	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel2	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel3	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel4	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel5	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel6	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel7	:	out	std_logic_vector(2 downto 0)	:=	"000";
		ev_128ns	:	out	std_logic	:=	'0';
		ev_1us	:	out	std_logic	:=	'0';
		flr_sts	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n0	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n1	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n2	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n3	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n4	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n5	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n6	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n7	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n0	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n1	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n2	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n3	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n4	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n5	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n6	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n7	:	out	std_logic	:=	'0';
		hotrst_exit	:	out	std_logic	:=	'0';
		int_status	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		k_hip_pcs_chnl_en	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		k_hrc_chnl_en	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		k_hrc_chnl_txpll_master_cgb_rst_en	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		k_hrc_chnl_txpll_rst_en	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		l2_exit	:	out	std_logic	:=	'0';
		lane_act	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		lmi_ack	:	out	std_logic	:=	'0';
		lmi_dout	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		ltssm_state	:	out	std_logic_vector(4 downto 0)	:=	"00000";
		mem_rscout_rcv_bot	:	out	std_logic	:=	'0';
		mem_rscout_rcv_top	:	out	std_logic	:=	'0';
		mem_rscout_rtry	:	out	std_logic	:=	'0';
		pld_clk_in_use	:	out	std_logic	:=	'0';
		pld_gp_ctrl	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		pm_exit_d0_req	:	out	std_logic	:=	'0';
		pme_to_sr	:	out	std_logic	:=	'0';
		powerdown0	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown1	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown2	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown3	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown4	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown5	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown6	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown7	:	out	std_logic_vector(1 downto 0)	:=	"00";
		r2c_unc_ecc	:	out	std_logic	:=	'0';
		rate0	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate1	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate2	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate3	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate4	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate5	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate6	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate7	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate_ctrl	:	out	std_logic_vector(1 downto 0)	:=	"00";
		reserved_clk_out	:	out	std_logic	:=	'0';
		reserved_out	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		reset_status	:	out	std_logic	:=	'0';
		retry_corr_ecc	:	out	std_logic	:=	'0';
		retry_unc_ecc	:	out	std_logic	:=	'0';
		rx_corr_ecc	:	out	std_logic	:=	'0';
		rx_cred_status	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		rx_par_err	:	out	std_logic	:=	'0';
		rx_pcs_rst_n0	:	out	std_logic	:=	'0';
		rx_pcs_rst_n1	:	out	std_logic	:=	'0';
		rx_pcs_rst_n2	:	out	std_logic	:=	'0';
		rx_pcs_rst_n3	:	out	std_logic	:=	'0';
		rx_pcs_rst_n4	:	out	std_logic	:=	'0';
		rx_pcs_rst_n5	:	out	std_logic	:=	'0';
		rx_pcs_rst_n6	:	out	std_logic	:=	'0';
		rx_pcs_rst_n7	:	out	std_logic	:=	'0';
		rx_pma_rstb0	:	out	std_logic	:=	'0';
		rx_pma_rstb1	:	out	std_logic	:=	'0';
		rx_pma_rstb2	:	out	std_logic	:=	'0';
		rx_pma_rstb3	:	out	std_logic	:=	'0';
		rx_pma_rstb4	:	out	std_logic	:=	'0';
		rx_pma_rstb5	:	out	std_logic	:=	'0';
		rx_pma_rstb6	:	out	std_logic	:=	'0';
		rx_pma_rstb7	:	out	std_logic	:=	'0';
		rx_st_bardec1	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		rx_st_bardec2	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		rx_st_be	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rx_st_data	:	out	std_logic_vector(255 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		rx_st_empty	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rx_st_eop	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		rx_st_err	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		rx_st_parity	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rx_st_sop	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		rx_st_valid	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		rxfc_cplbuf_ovf	:	out	std_logic	:=	'0';
		rxfc_cplovf_tag	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		rxpolarity0	:	out	std_logic	:=	'0';
		rxpolarity1	:	out	std_logic	:=	'0';
		rxpolarity2	:	out	std_logic	:=	'0';
		rxpolarity3	:	out	std_logic	:=	'0';
		rxpolarity4	:	out	std_logic	:=	'0';
		rxpolarity5	:	out	std_logic	:=	'0';
		rxpolarity6	:	out	std_logic	:=	'0';
		rxpolarity7	:	out	std_logic	:=	'0';
		serr_out	:	out	std_logic	:=	'0';
		swdn_out	:	out	std_logic_vector(6 downto 0)	:=	"0000000";
		swup_out	:	out	std_logic_vector(2 downto 0)	:=	"000";
		test_fref_clk	:	out	std_logic	:=	'0';
		test_out_1_hip	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		test_out_hip	:	out	std_logic_vector(255 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		tl_cfg_add	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		tl_cfg_ctl	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		tl_cfg_sts	:	out	std_logic_vector(52 downto 0)	:=	"00000000000000000000000000000000000000000000000000000";
		tl_cfg_sts_wr	:	out	std_logic	:=	'0';
		tx_cred_data_fc	:	out	std_logic_vector(11 downto 0)	:=	"000000000000";
		tx_cred_fc_hip_cons	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		tx_cred_fc_infinite	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		tx_cred_hdr_fc	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		tx_deemph0	:	out	std_logic	:=	'0';
		tx_deemph1	:	out	std_logic	:=	'0';
		tx_deemph2	:	out	std_logic	:=	'0';
		tx_deemph3	:	out	std_logic	:=	'0';
		tx_deemph4	:	out	std_logic	:=	'0';
		tx_deemph5	:	out	std_logic	:=	'0';
		tx_deemph6	:	out	std_logic	:=	'0';
		tx_deemph7	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb0	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb1	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb2	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb3	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb4	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb5	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb6	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb7	:	out	std_logic	:=	'0';
		tx_margin0	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin1	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin2	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin3	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin4	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin5	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin6	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin7	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_par_err	:	out	std_logic_vector(1 downto 0)	:=	"00";
		tx_pcs_rst_n0	:	out	std_logic	:=	'0';
		tx_pcs_rst_n1	:	out	std_logic	:=	'0';
		tx_pcs_rst_n2	:	out	std_logic	:=	'0';
		tx_pcs_rst_n3	:	out	std_logic	:=	'0';
		tx_pcs_rst_n4	:	out	std_logic	:=	'0';
		tx_pcs_rst_n5	:	out	std_logic	:=	'0';
		tx_pcs_rst_n6	:	out	std_logic	:=	'0';
		tx_pcs_rst_n7	:	out	std_logic	:=	'0';
		tx_pma_syncp0	:	out	std_logic	:=	'0';
		tx_pma_syncp1	:	out	std_logic	:=	'0';
		tx_pma_syncp2	:	out	std_logic	:=	'0';
		tx_pma_syncp3	:	out	std_logic	:=	'0';
		tx_pma_syncp4	:	out	std_logic	:=	'0';
		tx_pma_syncp5	:	out	std_logic	:=	'0';
		tx_pma_syncp6	:	out	std_logic	:=	'0';
		tx_pma_syncp7	:	out	std_logic	:=	'0';
		tx_st_ready	:	out	std_logic	:=	'0';
		txblkst0	:	out	std_logic	:=	'0';
		txblkst1	:	out	std_logic	:=	'0';
		txblkst2	:	out	std_logic	:=	'0';
		txblkst3	:	out	std_logic	:=	'0';
		txblkst4	:	out	std_logic	:=	'0';
		txblkst5	:	out	std_logic	:=	'0';
		txblkst6	:	out	std_logic	:=	'0';
		txblkst7	:	out	std_logic	:=	'0';
		txcompl0	:	out	std_logic	:=	'0';
		txcompl1	:	out	std_logic	:=	'0';
		txcompl2	:	out	std_logic	:=	'0';
		txcompl3	:	out	std_logic	:=	'0';
		txcompl4	:	out	std_logic	:=	'0';
		txcompl5	:	out	std_logic	:=	'0';
		txcompl6	:	out	std_logic	:=	'0';
		txcompl7	:	out	std_logic	:=	'0';
		txdata0	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata1	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata2	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata3	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata4	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata5	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata6	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata7	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdatak0	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak1	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak2	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak3	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak4	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak5	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak6	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak7	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdataskip0	:	out	std_logic	:=	'0';
		txdataskip1	:	out	std_logic	:=	'0';
		txdataskip2	:	out	std_logic	:=	'0';
		txdataskip3	:	out	std_logic	:=	'0';
		txdataskip4	:	out	std_logic	:=	'0';
		txdataskip5	:	out	std_logic	:=	'0';
		txdataskip6	:	out	std_logic	:=	'0';
		txdataskip7	:	out	std_logic	:=	'0';
		txdetectrx0	:	out	std_logic	:=	'0';
		txdetectrx1	:	out	std_logic	:=	'0';
		txdetectrx2	:	out	std_logic	:=	'0';
		txdetectrx3	:	out	std_logic	:=	'0';
		txdetectrx4	:	out	std_logic	:=	'0';
		txdetectrx5	:	out	std_logic	:=	'0';
		txdetectrx6	:	out	std_logic	:=	'0';
		txdetectrx7	:	out	std_logic	:=	'0';
		txelecidle0	:	out	std_logic	:=	'0';
		txelecidle1	:	out	std_logic	:=	'0';
		txelecidle2	:	out	std_logic	:=	'0';
		txelecidle3	:	out	std_logic	:=	'0';
		txelecidle4	:	out	std_logic	:=	'0';
		txelecidle5	:	out	std_logic	:=	'0';
		txelecidle6	:	out	std_logic	:=	'0';
		txelecidle7	:	out	std_logic	:=	'0';
		txst_prot_err	:	out	std_logic	:=	'0';
		txswing0	:	out	std_logic	:=	'0';
		txswing1	:	out	std_logic	:=	'0';
		txswing2	:	out	std_logic	:=	'0';
		txswing3	:	out	std_logic	:=	'0';
		txswing4	:	out	std_logic	:=	'0';
		txswing5	:	out	std_logic	:=	'0';
		txswing6	:	out	std_logic	:=	'0';
		txswing7	:	out	std_logic	:=	'0';
		txsynchd0	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd1	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd2	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd3	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd4	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd5	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd6	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd7	:	out	std_logic_vector(1 downto 0)	:=	"00";
		wake_oen	:	out	std_logic	:=	'0'
	);
end component;

begin



inst : twentynm_hssi_gen3_x8_pcie_hip_encrypted
	generic map (
		-- Instance parameters
		acknack_base	=>	acknack_base_int,
		acknack_set	=>	acknack_set,
		advance_error_reporting	=>	advance_error_reporting,
		app_interface_width	=>	app_interface_width,
		arb_upfc_30us_counter	=>	arb_upfc_30us_counter_int,
		arb_upfc_30us_en	=>	arb_upfc_30us_en,
		aspm_config_management	=>	aspm_config_management,
		aspm_patch_disable	=>	aspm_patch_disable,
		ast_width_rx	=>	ast_width_rx,
		ast_width_tx	=>	ast_width_tx,
		atomic_malformed	=>	atomic_malformed,
		atomic_op_completer_32bit	=>	atomic_op_completer_32bit,
		atomic_op_completer_64bit	=>	atomic_op_completer_64bit,
		atomic_op_routing	=>	atomic_op_routing,
		auto_msg_drop_enable	=>	auto_msg_drop_enable,
		avmm_cvp_inter_sel_csr_ctrl	=>	avmm_cvp_inter_sel_csr_ctrl,
		avmm_dprio_broadcast_en_csr_ctrl	=>	avmm_dprio_broadcast_en_csr_ctrl,
		avmm_force_inter_sel_csr_ctrl	=>	avmm_force_inter_sel_csr_ctrl,
		avmm_power_iso_en_csr_ctrl	=>	avmm_power_iso_en_csr_ctrl,
		bar0_size_mask	=>	bar0_size_mask_int,
		bar0_type	=>	bar0_type,
		bar1_size_mask	=>	bar1_size_mask_int,
		bar1_type	=>	bar1_type,
		bar2_size_mask	=>	bar2_size_mask_int,
		bar2_type	=>	bar2_type,
		bar3_size_mask	=>	bar3_size_mask_int,
		bar3_type	=>	bar3_type,
		bar4_size_mask	=>	bar4_size_mask_int,
		bar4_type	=>	bar4_type,
		bar5_size_mask	=>	bar5_size_mask_int,
		bar5_type	=>	bar5_type,
		base_counter_sel	=>	base_counter_sel,
		bist_memory_settings	=>	bist_memory_settings,
		bridge_port_ssid_support	=>	bridge_port_ssid_support,
		bridge_port_vga_enable	=>	bridge_port_vga_enable,
		bypass_cdc	=>	bypass_cdc,
		bypass_clk_switch	=>	bypass_clk_switch,
		bypass_tl	=>	bypass_tl,
		capab_rate_rxcfg_en	=>	capab_rate_rxcfg_en,
		cas_completer_128bit	=>	cas_completer_128bit,
		cdc_clk_relation	=>	cdc_clk_relation,
		cdc_dummy_insert_limit	=>	cdc_dummy_insert_limit_int,
		cfg_parchk_ena	=>	cfg_parchk_ena,
		cfgbp_req_recov_disable	=>	cfgbp_req_recov_disable,
		class_code	=>	class_code_int,
		clock_pwr_management	=>	clock_pwr_management,
		completion_timeout	=>	completion_timeout,
		core_clk_divider	=>	core_clk_divider,
		core_clk_freq_mhz	=>	core_clk_freq_mhz,
		core_clk_out_sel	=>	core_clk_out_sel,
		core_clk_sel	=>	core_clk_sel,
		core_clk_source	=>	core_clk_source,
		cseb_bar_match_checking	=>	cseb_bar_match_checking,
		cseb_config_bypass	=>	cseb_config_bypass,
		cseb_cpl_status_during_cvp	=>	cseb_cpl_status_during_cvp,
		cseb_cpl_tag_checking	=>	cseb_cpl_tag_checking,
		cseb_disable_auto_crs	=>	cseb_disable_auto_crs,
		cseb_extend_pci	=>	cseb_extend_pci,
		cseb_extend_pcie	=>	cseb_extend_pcie,
		cseb_min_error_checking	=>	cseb_min_error_checking,
		cseb_route_to_avl_rx_st	=>	cseb_route_to_avl_rx_st,
		cseb_temp_busy_crs	=>	cseb_temp_busy_crs,
		cvp_clk_reset	=>	cvp_clk_reset,
		cvp_data_compressed	=>	cvp_data_compressed,
		cvp_data_encrypted	=>	cvp_data_encrypted,
		cvp_enable	=>	cvp_enable,
		cvp_mode_reset	=>	cvp_mode_reset,
		cvp_rate_sel	=>	cvp_rate_sel,
		d0_pme	=>	d0_pme,
		d1_pme	=>	d1_pme,
		d1_support	=>	d1_support,
		d2_pme	=>	d2_pme,
		d2_support	=>	d2_support,
		d3_cold_pme	=>	d3_cold_pme,
		d3_hot_pme	=>	d3_hot_pme,
		data_pack_rx	=>	data_pack_rx,
		deemphasis_enable	=>	deemphasis_enable,
		deskew_comma	=>	deskew_comma,
		device_id	=>	device_id_int,
		device_number	=>	device_number_int,
		device_specific_init	=>	device_specific_init,
		dft_clock_obsrv_en	=>	dft_clock_obsrv_en,
		dft_clock_obsrv_sel	=>	dft_clock_obsrv_sel,
		diffclock_nfts_count	=>	diffclock_nfts_count_int,
		dis_cplovf	=>	dis_cplovf,
		dis_paritychk	=>	dis_paritychk,
		disable_link_x2_support	=>	disable_link_x2_support,
		disable_snoop_packet	=>	disable_snoop_packet,
		dl_tx_check_parity_edb	=>	dl_tx_check_parity_edb,
		dll_active_report_support	=>	dll_active_report_support,
		early_dl_up	=>	early_dl_up,
		eco_fb332688_dis	=>	eco_fb332688_dis,
		ecrc_check_capable	=>	ecrc_check_capable,
		ecrc_gen_capable	=>	ecrc_gen_capable,
		egress_block_err_report_ena	=>	egress_block_err_report_ena,
		ei_delay_powerdown_count	=>	ei_delay_powerdown_count_int,
		eie_before_nfts_count	=>	eie_before_nfts_count_int,
		electromech_interlock	=>	electromech_interlock,
		en_ieiupdatefc	=>	en_ieiupdatefc,
		en_lane_errchk	=>	en_lane_errchk,
		en_phystatus_dly	=>	en_phystatus_dly,
		ena_ido_cpl	=>	ena_ido_cpl,
		ena_ido_req	=>	ena_ido_req,
		enable_adapter_half_rate_mode	=>	enable_adapter_half_rate_mode,
		enable_ch01_pclk_out	=>	enable_ch01_pclk_out,
		enable_ch0_pclk_out	=>	enable_ch0_pclk_out,
		enable_completion_timeout_disable	=>	enable_completion_timeout_disable,
		enable_directed_spd_chng	=>	enable_directed_spd_chng,
		enable_function_msix_support	=>	enable_function_msix_support,
		enable_l0s_aspm	=>	enable_l0s_aspm,
		enable_l1_aspm	=>	enable_l1_aspm,
		enable_rx_buffer_checking	=>	enable_rx_buffer_checking,
		enable_rx_reordering	=>	enable_rx_reordering,
		enable_slot_register	=>	enable_slot_register,
		endpoint_l0_latency	=>	endpoint_l0_latency_int,
		endpoint_l1_latency	=>	endpoint_l1_latency_int,
		eql_rq_int_en_number	=>	eql_rq_int_en_number_int,
		errmgt_fcpe_patch_dis	=>	errmgt_fcpe_patch_dis,
		errmgt_fep_patch_dis	=>	errmgt_fep_patch_dis,
		expansion_base_address_register	=>	expansion_base_address_register,
		extend_tag_field	=>	extend_tag_field,
		extended_format_field	=>	extended_format_field,
		extended_tag_reset	=>	extended_tag_reset,
		fc_init_timer	=>	fc_init_timer_int,
		flow_control_timeout_count	=>	flow_control_timeout_count_int,
		flow_control_update_count	=>	flow_control_update_count_int,
		flr_capability	=>	flr_capability,
		force_dis_to_det	=>	force_dis_to_det,
		force_gen1_dis	=>	force_gen1_dis,
		force_tx_coeff_preset_lpbk	=>	force_tx_coeff_preset_lpbk,
		frame_err_patch_dis	=>	frame_err_patch_dis,
		func_mode	=>	func_mode,
		g3_bypass_equlz	=>	g3_bypass_equlz,
		g3_coeff_done_tmout	=>	g3_coeff_done_tmout,
		g3_deskew_char	=>	g3_deskew_char,
		g3_dis_be_frm_err	=>	g3_dis_be_frm_err,
		g3_dn_rx_hint_eqlz_0	=>	g3_dn_rx_hint_eqlz_0_int,
		g3_dn_rx_hint_eqlz_1	=>	g3_dn_rx_hint_eqlz_1_int,
		g3_dn_rx_hint_eqlz_2	=>	g3_dn_rx_hint_eqlz_2_int,
		g3_dn_rx_hint_eqlz_3	=>	g3_dn_rx_hint_eqlz_3_int,
		g3_dn_rx_hint_eqlz_4	=>	g3_dn_rx_hint_eqlz_4_int,
		g3_dn_rx_hint_eqlz_5	=>	g3_dn_rx_hint_eqlz_5_int,
		g3_dn_rx_hint_eqlz_6	=>	g3_dn_rx_hint_eqlz_6_int,
		g3_dn_rx_hint_eqlz_7	=>	g3_dn_rx_hint_eqlz_7_int,
		g3_dn_tx_preset_eqlz_0	=>	g3_dn_tx_preset_eqlz_0_int,
		g3_dn_tx_preset_eqlz_1	=>	g3_dn_tx_preset_eqlz_1_int,
		g3_dn_tx_preset_eqlz_2	=>	g3_dn_tx_preset_eqlz_2_int,
		g3_dn_tx_preset_eqlz_3	=>	g3_dn_tx_preset_eqlz_3_int,
		g3_dn_tx_preset_eqlz_4	=>	g3_dn_tx_preset_eqlz_4_int,
		g3_dn_tx_preset_eqlz_5	=>	g3_dn_tx_preset_eqlz_5_int,
		g3_dn_tx_preset_eqlz_6	=>	g3_dn_tx_preset_eqlz_6_int,
		g3_dn_tx_preset_eqlz_7	=>	g3_dn_tx_preset_eqlz_7_int,
		g3_force_ber_max	=>	g3_force_ber_max,
		g3_force_ber_min	=>	g3_force_ber_min,
		g3_lnk_trn_rx_ts	=>	g3_lnk_trn_rx_ts,
		g3_ltssm_eq_dbg	=>	g3_ltssm_eq_dbg,
		g3_ltssm_rec_dbg	=>	g3_ltssm_rec_dbg,
		g3_pause_ltssm_rec_en	=>	g3_pause_ltssm_rec_en,
		g3_quiesce_guarant	=>	g3_quiesce_guarant,
		g3_redo_equlz_dis	=>	g3_redo_equlz_dis,
		g3_redo_equlz_en	=>	g3_redo_equlz_en,
		g3_up_rx_hint_eqlz_0	=>	g3_up_rx_hint_eqlz_0_int,
		g3_up_rx_hint_eqlz_1	=>	g3_up_rx_hint_eqlz_1_int,
		g3_up_rx_hint_eqlz_2	=>	g3_up_rx_hint_eqlz_2_int,
		g3_up_rx_hint_eqlz_3	=>	g3_up_rx_hint_eqlz_3_int,
		g3_up_rx_hint_eqlz_4	=>	g3_up_rx_hint_eqlz_4_int,
		g3_up_rx_hint_eqlz_5	=>	g3_up_rx_hint_eqlz_5_int,
		g3_up_rx_hint_eqlz_6	=>	g3_up_rx_hint_eqlz_6_int,
		g3_up_rx_hint_eqlz_7	=>	g3_up_rx_hint_eqlz_7_int,
		g3_up_tx_preset_eqlz_0	=>	g3_up_tx_preset_eqlz_0_int,
		g3_up_tx_preset_eqlz_1	=>	g3_up_tx_preset_eqlz_1_int,
		g3_up_tx_preset_eqlz_2	=>	g3_up_tx_preset_eqlz_2_int,
		g3_up_tx_preset_eqlz_3	=>	g3_up_tx_preset_eqlz_3_int,
		g3_up_tx_preset_eqlz_4	=>	g3_up_tx_preset_eqlz_4_int,
		g3_up_tx_preset_eqlz_5	=>	g3_up_tx_preset_eqlz_5_int,
		g3_up_tx_preset_eqlz_6	=>	g3_up_tx_preset_eqlz_6_int,
		g3_up_tx_preset_eqlz_7	=>	g3_up_tx_preset_eqlz_7_int,
		gen123_lane_rate_mode	=>	gen123_lane_rate_mode,
		gen2_diffclock_nfts_count	=>	gen2_diffclock_nfts_count_int,
		gen2_pma_pll_usage	=>	gen2_pma_pll_usage,
		gen2_sameclock_nfts_count	=>	gen2_sameclock_nfts_count_int,
		gen3_coeff_1	=>	gen3_coeff_1_int,
		gen3_coeff_10	=>	gen3_coeff_10_int,
		gen3_coeff_10_ber_meas	=>	gen3_coeff_10_ber_meas_int,
		gen3_coeff_10_nxtber_less	=>	gen3_coeff_10_nxtber_less_int,
		gen3_coeff_10_nxtber_more	=>	gen3_coeff_10_nxtber_more_int,
		gen3_coeff_10_preset_hint	=>	gen3_coeff_10_preset_hint_int,
		gen3_coeff_10_reqber	=>	gen3_coeff_10_reqber_int,
		gen3_coeff_10_sel	=>	gen3_coeff_10_sel,
		gen3_coeff_11	=>	gen3_coeff_11_int,
		gen3_coeff_11_ber_meas	=>	gen3_coeff_11_ber_meas_int,
		gen3_coeff_11_nxtber_less	=>	gen3_coeff_11_nxtber_less_int,
		gen3_coeff_11_nxtber_more	=>	gen3_coeff_11_nxtber_more_int,
		gen3_coeff_11_preset_hint	=>	gen3_coeff_11_preset_hint_int,
		gen3_coeff_11_reqber	=>	gen3_coeff_11_reqber_int,
		gen3_coeff_11_sel	=>	gen3_coeff_11_sel,
		gen3_coeff_12	=>	gen3_coeff_12_int,
		gen3_coeff_12_ber_meas	=>	gen3_coeff_12_ber_meas_int,
		gen3_coeff_12_nxtber_less	=>	gen3_coeff_12_nxtber_less_int,
		gen3_coeff_12_nxtber_more	=>	gen3_coeff_12_nxtber_more_int,
		gen3_coeff_12_preset_hint	=>	gen3_coeff_12_preset_hint_int,
		gen3_coeff_12_reqber	=>	gen3_coeff_12_reqber_int,
		gen3_coeff_12_sel	=>	gen3_coeff_12_sel,
		gen3_coeff_13	=>	gen3_coeff_13_int,
		gen3_coeff_13_ber_meas	=>	gen3_coeff_13_ber_meas_int,
		gen3_coeff_13_nxtber_less	=>	gen3_coeff_13_nxtber_less_int,
		gen3_coeff_13_nxtber_more	=>	gen3_coeff_13_nxtber_more_int,
		gen3_coeff_13_preset_hint	=>	gen3_coeff_13_preset_hint_int,
		gen3_coeff_13_reqber	=>	gen3_coeff_13_reqber_int,
		gen3_coeff_13_sel	=>	gen3_coeff_13_sel,
		gen3_coeff_14	=>	gen3_coeff_14_int,
		gen3_coeff_14_ber_meas	=>	gen3_coeff_14_ber_meas_int,
		gen3_coeff_14_nxtber_less	=>	gen3_coeff_14_nxtber_less_int,
		gen3_coeff_14_nxtber_more	=>	gen3_coeff_14_nxtber_more_int,
		gen3_coeff_14_preset_hint	=>	gen3_coeff_14_preset_hint_int,
		gen3_coeff_14_reqber	=>	gen3_coeff_14_reqber_int,
		gen3_coeff_14_sel	=>	gen3_coeff_14_sel,
		gen3_coeff_15	=>	gen3_coeff_15_int,
		gen3_coeff_15_ber_meas	=>	gen3_coeff_15_ber_meas_int,
		gen3_coeff_15_nxtber_less	=>	gen3_coeff_15_nxtber_less_int,
		gen3_coeff_15_nxtber_more	=>	gen3_coeff_15_nxtber_more_int,
		gen3_coeff_15_preset_hint	=>	gen3_coeff_15_preset_hint_int,
		gen3_coeff_15_reqber	=>	gen3_coeff_15_reqber_int,
		gen3_coeff_15_sel	=>	gen3_coeff_15_sel,
		gen3_coeff_16	=>	gen3_coeff_16_int,
		gen3_coeff_16_ber_meas	=>	gen3_coeff_16_ber_meas_int,
		gen3_coeff_16_nxtber_less	=>	gen3_coeff_16_nxtber_less_int,
		gen3_coeff_16_nxtber_more	=>	gen3_coeff_16_nxtber_more_int,
		gen3_coeff_16_preset_hint	=>	gen3_coeff_16_preset_hint_int,
		gen3_coeff_16_reqber	=>	gen3_coeff_16_reqber_int,
		gen3_coeff_16_sel	=>	gen3_coeff_16_sel,
		gen3_coeff_17	=>	gen3_coeff_17_int,
		gen3_coeff_17_ber_meas	=>	gen3_coeff_17_ber_meas_int,
		gen3_coeff_17_nxtber_less	=>	gen3_coeff_17_nxtber_less_int,
		gen3_coeff_17_nxtber_more	=>	gen3_coeff_17_nxtber_more_int,
		gen3_coeff_17_preset_hint	=>	gen3_coeff_17_preset_hint_int,
		gen3_coeff_17_reqber	=>	gen3_coeff_17_reqber_int,
		gen3_coeff_17_sel	=>	gen3_coeff_17_sel,
		gen3_coeff_18	=>	gen3_coeff_18_int,
		gen3_coeff_18_ber_meas	=>	gen3_coeff_18_ber_meas_int,
		gen3_coeff_18_nxtber_less	=>	gen3_coeff_18_nxtber_less_int,
		gen3_coeff_18_nxtber_more	=>	gen3_coeff_18_nxtber_more_int,
		gen3_coeff_18_preset_hint	=>	gen3_coeff_18_preset_hint_int,
		gen3_coeff_18_reqber	=>	gen3_coeff_18_reqber_int,
		gen3_coeff_18_sel	=>	gen3_coeff_18_sel,
		gen3_coeff_19	=>	gen3_coeff_19_int,
		gen3_coeff_19_ber_meas	=>	gen3_coeff_19_ber_meas_int,
		gen3_coeff_19_nxtber_less	=>	gen3_coeff_19_nxtber_less_int,
		gen3_coeff_19_nxtber_more	=>	gen3_coeff_19_nxtber_more_int,
		gen3_coeff_19_preset_hint	=>	gen3_coeff_19_preset_hint_int,
		gen3_coeff_19_reqber	=>	gen3_coeff_19_reqber_int,
		gen3_coeff_19_sel	=>	gen3_coeff_19_sel,
		gen3_coeff_1_ber_meas	=>	gen3_coeff_1_ber_meas_int,
		gen3_coeff_1_nxtber_less	=>	gen3_coeff_1_nxtber_less_int,
		gen3_coeff_1_nxtber_more	=>	gen3_coeff_1_nxtber_more_int,
		gen3_coeff_1_preset_hint	=>	gen3_coeff_1_preset_hint_int,
		gen3_coeff_1_reqber	=>	gen3_coeff_1_reqber_int,
		gen3_coeff_1_sel	=>	gen3_coeff_1_sel,
		gen3_coeff_2	=>	gen3_coeff_2_int,
		gen3_coeff_20	=>	gen3_coeff_20_int,
		gen3_coeff_20_ber_meas	=>	gen3_coeff_20_ber_meas_int,
		gen3_coeff_20_nxtber_less	=>	gen3_coeff_20_nxtber_less_int,
		gen3_coeff_20_nxtber_more	=>	gen3_coeff_20_nxtber_more_int,
		gen3_coeff_20_preset_hint	=>	gen3_coeff_20_preset_hint_int,
		gen3_coeff_20_reqber	=>	gen3_coeff_20_reqber_int,
		gen3_coeff_20_sel	=>	gen3_coeff_20_sel,
		gen3_coeff_21	=>	gen3_coeff_21_int,
		gen3_coeff_21_ber_meas	=>	gen3_coeff_21_ber_meas_int,
		gen3_coeff_21_nxtber_less	=>	gen3_coeff_21_nxtber_less_int,
		gen3_coeff_21_nxtber_more	=>	gen3_coeff_21_nxtber_more_int,
		gen3_coeff_21_preset_hint	=>	gen3_coeff_21_preset_hint_int,
		gen3_coeff_21_reqber	=>	gen3_coeff_21_reqber_int,
		gen3_coeff_21_sel	=>	gen3_coeff_21_sel,
		gen3_coeff_22	=>	gen3_coeff_22_int,
		gen3_coeff_22_ber_meas	=>	gen3_coeff_22_ber_meas_int,
		gen3_coeff_22_nxtber_less	=>	gen3_coeff_22_nxtber_less_int,
		gen3_coeff_22_nxtber_more	=>	gen3_coeff_22_nxtber_more_int,
		gen3_coeff_22_preset_hint	=>	gen3_coeff_22_preset_hint_int,
		gen3_coeff_22_reqber	=>	gen3_coeff_22_reqber_int,
		gen3_coeff_22_sel	=>	gen3_coeff_22_sel,
		gen3_coeff_23	=>	gen3_coeff_23_int,
		gen3_coeff_23_ber_meas	=>	gen3_coeff_23_ber_meas_int,
		gen3_coeff_23_nxtber_less	=>	gen3_coeff_23_nxtber_less_int,
		gen3_coeff_23_nxtber_more	=>	gen3_coeff_23_nxtber_more_int,
		gen3_coeff_23_preset_hint	=>	gen3_coeff_23_preset_hint_int,
		gen3_coeff_23_reqber	=>	gen3_coeff_23_reqber_int,
		gen3_coeff_23_sel	=>	gen3_coeff_23_sel,
		gen3_coeff_24	=>	gen3_coeff_24_int,
		gen3_coeff_24_ber_meas	=>	gen3_coeff_24_ber_meas_int,
		gen3_coeff_24_nxtber_less	=>	gen3_coeff_24_nxtber_less_int,
		gen3_coeff_24_nxtber_more	=>	gen3_coeff_24_nxtber_more_int,
		gen3_coeff_24_preset_hint	=>	gen3_coeff_24_preset_hint_int,
		gen3_coeff_24_reqber	=>	gen3_coeff_24_reqber_int,
		gen3_coeff_24_sel	=>	gen3_coeff_24_sel,
		gen3_coeff_2_ber_meas	=>	gen3_coeff_2_ber_meas_int,
		gen3_coeff_2_nxtber_less	=>	gen3_coeff_2_nxtber_less_int,
		gen3_coeff_2_nxtber_more	=>	gen3_coeff_2_nxtber_more_int,
		gen3_coeff_2_preset_hint	=>	gen3_coeff_2_preset_hint_int,
		gen3_coeff_2_reqber	=>	gen3_coeff_2_reqber_int,
		gen3_coeff_2_sel	=>	gen3_coeff_2_sel,
		gen3_coeff_3	=>	gen3_coeff_3_int,
		gen3_coeff_3_ber_meas	=>	gen3_coeff_3_ber_meas_int,
		gen3_coeff_3_nxtber_less	=>	gen3_coeff_3_nxtber_less_int,
		gen3_coeff_3_nxtber_more	=>	gen3_coeff_3_nxtber_more_int,
		gen3_coeff_3_preset_hint	=>	gen3_coeff_3_preset_hint_int,
		gen3_coeff_3_reqber	=>	gen3_coeff_3_reqber_int,
		gen3_coeff_3_sel	=>	gen3_coeff_3_sel,
		gen3_coeff_4	=>	gen3_coeff_4_int,
		gen3_coeff_4_ber_meas	=>	gen3_coeff_4_ber_meas_int,
		gen3_coeff_4_nxtber_less	=>	gen3_coeff_4_nxtber_less_int,
		gen3_coeff_4_nxtber_more	=>	gen3_coeff_4_nxtber_more_int,
		gen3_coeff_4_preset_hint	=>	gen3_coeff_4_preset_hint_int,
		gen3_coeff_4_reqber	=>	gen3_coeff_4_reqber_int,
		gen3_coeff_4_sel	=>	gen3_coeff_4_sel,
		gen3_coeff_5	=>	gen3_coeff_5_int,
		gen3_coeff_5_ber_meas	=>	gen3_coeff_5_ber_meas_int,
		gen3_coeff_5_nxtber_less	=>	gen3_coeff_5_nxtber_less_int,
		gen3_coeff_5_nxtber_more	=>	gen3_coeff_5_nxtber_more_int,
		gen3_coeff_5_preset_hint	=>	gen3_coeff_5_preset_hint_int,
		gen3_coeff_5_reqber	=>	gen3_coeff_5_reqber_int,
		gen3_coeff_5_sel	=>	gen3_coeff_5_sel,
		gen3_coeff_6	=>	gen3_coeff_6_int,
		gen3_coeff_6_ber_meas	=>	gen3_coeff_6_ber_meas_int,
		gen3_coeff_6_nxtber_less	=>	gen3_coeff_6_nxtber_less_int,
		gen3_coeff_6_nxtber_more	=>	gen3_coeff_6_nxtber_more_int,
		gen3_coeff_6_preset_hint	=>	gen3_coeff_6_preset_hint_int,
		gen3_coeff_6_reqber	=>	gen3_coeff_6_reqber_int,
		gen3_coeff_6_sel	=>	gen3_coeff_6_sel,
		gen3_coeff_7	=>	gen3_coeff_7_int,
		gen3_coeff_7_ber_meas	=>	gen3_coeff_7_ber_meas_int,
		gen3_coeff_7_nxtber_less	=>	gen3_coeff_7_nxtber_less_int,
		gen3_coeff_7_nxtber_more	=>	gen3_coeff_7_nxtber_more_int,
		gen3_coeff_7_preset_hint	=>	gen3_coeff_7_preset_hint_int,
		gen3_coeff_7_reqber	=>	gen3_coeff_7_reqber_int,
		gen3_coeff_7_sel	=>	gen3_coeff_7_sel,
		gen3_coeff_8	=>	gen3_coeff_8_int,
		gen3_coeff_8_ber_meas	=>	gen3_coeff_8_ber_meas_int,
		gen3_coeff_8_nxtber_less	=>	gen3_coeff_8_nxtber_less_int,
		gen3_coeff_8_nxtber_more	=>	gen3_coeff_8_nxtber_more_int,
		gen3_coeff_8_preset_hint	=>	gen3_coeff_8_preset_hint_int,
		gen3_coeff_8_reqber	=>	gen3_coeff_8_reqber_int,
		gen3_coeff_8_sel	=>	gen3_coeff_8_sel,
		gen3_coeff_9	=>	gen3_coeff_9_int,
		gen3_coeff_9_ber_meas	=>	gen3_coeff_9_ber_meas_int,
		gen3_coeff_9_nxtber_less	=>	gen3_coeff_9_nxtber_less_int,
		gen3_coeff_9_nxtber_more	=>	gen3_coeff_9_nxtber_more_int,
		gen3_coeff_9_preset_hint	=>	gen3_coeff_9_preset_hint_int,
		gen3_coeff_9_reqber	=>	gen3_coeff_9_reqber_int,
		gen3_coeff_9_sel	=>	gen3_coeff_9_sel,
		gen3_coeff_delay_count	=>	gen3_coeff_delay_count_int,
		gen3_coeff_errchk	=>	gen3_coeff_errchk,
		gen3_dcbal_en	=>	gen3_dcbal_en,
		gen3_diffclock_nfts_count	=>	gen3_diffclock_nfts_count_int,
		gen3_force_local_coeff	=>	gen3_force_local_coeff,
		gen3_full_swing	=>	gen3_full_swing_int,
		gen3_half_swing	=>	gen3_half_swing,
		gen3_low_freq	=>	gen3_low_freq_int,
		gen3_paritychk	=>	gen3_paritychk,
		gen3_pl_framing_err_dis	=>	gen3_pl_framing_err_dis,
		gen3_preset_coeff_1	=>	gen3_preset_coeff_1_int,
		gen3_preset_coeff_10	=>	gen3_preset_coeff_10_int,
		gen3_preset_coeff_11	=>	gen3_preset_coeff_11_int,
		gen3_preset_coeff_2	=>	gen3_preset_coeff_2_int,
		gen3_preset_coeff_3	=>	gen3_preset_coeff_3_int,
		gen3_preset_coeff_4	=>	gen3_preset_coeff_4_int,
		gen3_preset_coeff_5	=>	gen3_preset_coeff_5_int,
		gen3_preset_coeff_6	=>	gen3_preset_coeff_6_int,
		gen3_preset_coeff_7	=>	gen3_preset_coeff_7_int,
		gen3_preset_coeff_8	=>	gen3_preset_coeff_8_int,
		gen3_preset_coeff_9	=>	gen3_preset_coeff_9_int,
		gen3_reset_eieos_cnt_bit	=>	gen3_reset_eieos_cnt_bit,
		gen3_rxfreqlock_counter	=>	gen3_rxfreqlock_counter_int,
		gen3_sameclock_nfts_count	=>	gen3_sameclock_nfts_count_int,
		gen3_scrdscr_bypass	=>	gen3_scrdscr_bypass,
		gen3_skip_ph2_ph3	=>	gen3_skip_ph2_ph3,
		hard_reset_bypass	=>	hard_reset_bypass,
		hard_rst_sig_chnl_en	=>	hard_rst_sig_chnl_en,
		hard_rst_tx_pll_rst_chnl_en	=>	hard_rst_tx_pll_rst_chnl_en,
		hip_ac_pwr_clk_freq_in_hz	=>	hip_ac_pwr_clk_freq_in_hz_int,
		hip_ac_pwr_uw_per_mhz	=>	hip_ac_pwr_uw_per_mhz_int,
		hip_base_address	=>	hip_base_address_int,
		hip_clock_dis	=>	hip_clock_dis,
		hip_hard_reset	=>	hip_hard_reset,
		hip_pcs_sig_chnl_en	=>	hip_pcs_sig_chnl_en,
		hot_plug_support	=>	hot_plug_support_int,
		hrc_chnl_txpll_master_cgb_rst_select	=>	hrc_chnl_txpll_master_cgb_rst_select,
		hrdrstctrl_en	=>	hrdrstctrl_en,
		iei_enable_settings	=>	iei_enable_settings,
		indicator	=>	indicator_int,
		intel_id_access	=>	intel_id_access,
		interrupt_pin	=>	interrupt_pin,
		io_window_addr_width	=>	io_window_addr_width,
		jtag_id	=>	jtag_id,
		ko_compl_data	=>	ko_compl_data_int,
		ko_compl_header	=>	ko_compl_header_int,
		l01_entry_latency	=>	l01_entry_latency_int,
		l0_exit_latency_diffclock	=>	l0_exit_latency_diffclock_int,
		l0_exit_latency_sameclock	=>	l0_exit_latency_sameclock_int,
		l0s_adj_rply_timer_dis	=>	l0s_adj_rply_timer_dis,
		l1_exit_latency_diffclock	=>	l1_exit_latency_diffclock_int,
		l1_exit_latency_sameclock	=>	l1_exit_latency_sameclock_int,
		l2_async_logic	=>	l2_async_logic,
		lane_mask	=>	lane_mask,
		lane_rate	=>	lane_rate,
		link_width	=>	link_width,
		lmi_hold_off_cfg_timer_en	=>	lmi_hold_off_cfg_timer_en,
		low_priority_vc	=>	low_priority_vc,
		ltr_mechanism	=>	ltr_mechanism,
		ltssm_1ms_timeout	=>	ltssm_1ms_timeout,
		ltssm_freqlocked_check	=>	ltssm_freqlocked_check,
		malformed_tlp_truncate_en	=>	malformed_tlp_truncate_en,
		max_link_width	=>	max_link_width,
		max_payload_size	=>	max_payload_size,
		maximum_current	=>	maximum_current_int,
		millisecond_cycle_count	=>	millisecond_cycle_count_int,
		msi_64bit_addressing_capable	=>	msi_64bit_addressing_capable,
		msi_masking_capable	=>	msi_masking_capable,
		msi_multi_message_capable	=>	msi_multi_message_capable,
		msi_support	=>	msi_support,
		msix_pba_bir	=>	msix_pba_bir_int,
		msix_pba_offset	=>	msix_pba_offset_int,
		msix_table_bir	=>	msix_table_bir_int,
		msix_table_offset	=>	msix_table_offset_int,
		msix_table_size	=>	msix_table_size_int,
		national_inst_thru_enhance	=>	national_inst_thru_enhance,
		no_command_completed	=>	no_command_completed,
		no_soft_reset	=>	no_soft_reset,
		not_use_k_gbl_bits	=>	not_use_k_gbl_bits,
		operating_voltage	=>	operating_voltage,
		pcie_base_spec	=>	pcie_base_spec,
		pcie_mode	=>	pcie_mode,
		pcie_spec_1p0_compliance	=>	pcie_spec_1p0_compliance,
		pcie_spec_version	=>	pcie_spec_version,
		pclk_out_sel	=>	pclk_out_sel,
		pld_in_use_reg	=>	pld_in_use_reg,
		pm_latency_patch_dis	=>	pm_latency_patch_dis,
		pm_txdl_patch_dis	=>	pm_txdl_patch_dis,
		pme_clock	=>	pme_clock,
		port_link_number	=>	port_link_number_int,
		port_type	=>	port_type,
		powerdown_mode	=>	powerdown_mode,
		prefetchable_mem_window_addr_width	=>	prefetchable_mem_window_addr_width,
		r2c_mask_easy	=>	r2c_mask_easy,
		r2c_mask_enable	=>	r2c_mask_enable,
		rec_frqlk_mon_en	=>	rec_frqlk_mon_en,
		register_pipe_signals	=>	register_pipe_signals,
		retry_buffer_last_active_address	=>	retry_buffer_last_active_address_int,
		retry_buffer_memory_settings	=>	retry_buffer_memory_settings,
		retry_ecc_corr_mask_dis	=>	retry_ecc_corr_mask_dis,
		revision_id	=>	revision_id_int,
		role_based_error_reporting	=>	role_based_error_reporting,
		rp_bug_fix_pri_sec_stat_reg	=>	rp_bug_fix_pri_sec_stat_reg_int,
		rpltim_base	=>	rpltim_base_int,
		rpltim_set	=>	rpltim_set,
		rstctl_ltssm_dis	=>	rstctl_ltssm_dis,
		rstctrl_1ms_count_fref_clk	=>	rstctrl_1ms_count_fref_clk_int,
		rstctrl_1us_count_fref_clk	=>	rstctrl_1us_count_fref_clk_int,
		rstctrl_altpe3_crst_n_inv	=>	rstctrl_altpe3_crst_n_inv,
		rstctrl_altpe3_rst_n_inv	=>	rstctrl_altpe3_rst_n_inv,
		rstctrl_altpe3_srst_n_inv	=>	rstctrl_altpe3_srst_n_inv,
		rstctrl_chnl_cal_done_select	=>	rstctrl_chnl_cal_done_select,
		rstctrl_debug_en	=>	rstctrl_debug_en,
		rstctrl_force_inactive_rst	=>	rstctrl_force_inactive_rst,
		rstctrl_fref_clk_select	=>	rstctrl_fref_clk_select,
		rstctrl_hard_block_enable	=>	rstctrl_hard_block_enable,
		rstctrl_hip_ep	=>	rstctrl_hip_ep,
		rstctrl_mask_tx_pll_lock_select	=>	rstctrl_mask_tx_pll_lock_select,
		rstctrl_perst_enable	=>	rstctrl_perst_enable,
		rstctrl_perstn_select	=>	rstctrl_perstn_select,
		rstctrl_pld_clr	=>	rstctrl_pld_clr,
		rstctrl_pll_cal_done_select	=>	rstctrl_pll_cal_done_select,
		rstctrl_rx_pcs_rst_n_inv	=>	rstctrl_rx_pcs_rst_n_inv,
		rstctrl_rx_pcs_rst_n_select	=>	rstctrl_rx_pcs_rst_n_select,
		rstctrl_rx_pll_freq_lock_select	=>	rstctrl_rx_pll_freq_lock_select,
		rstctrl_rx_pll_lock_select	=>	rstctrl_rx_pll_lock_select,
		rstctrl_rx_pma_rstb_inv	=>	rstctrl_rx_pma_rstb_inv,
		rstctrl_rx_pma_rstb_select	=>	rstctrl_rx_pma_rstb_select,
		rstctrl_timer_a	=>	rstctrl_timer_a_int,
		rstctrl_timer_a_type	=>	rstctrl_timer_a_type,
		rstctrl_timer_b	=>	rstctrl_timer_b_int,
		rstctrl_timer_b_type	=>	rstctrl_timer_b_type,
		rstctrl_timer_c	=>	rstctrl_timer_c_int,
		rstctrl_timer_c_type	=>	rstctrl_timer_c_type,
		rstctrl_timer_d	=>	rstctrl_timer_d_int,
		rstctrl_timer_d_type	=>	rstctrl_timer_d_type,
		rstctrl_timer_e	=>	rstctrl_timer_e_int,
		rstctrl_timer_e_type	=>	rstctrl_timer_e_type,
		rstctrl_timer_f	=>	rstctrl_timer_f_int,
		rstctrl_timer_f_type	=>	rstctrl_timer_f_type,
		rstctrl_timer_g	=>	rstctrl_timer_g_int,
		rstctrl_timer_g_type	=>	rstctrl_timer_g_type,
		rstctrl_timer_h	=>	rstctrl_timer_h_int,
		rstctrl_timer_h_type	=>	rstctrl_timer_h_type,
		rstctrl_timer_i	=>	rstctrl_timer_i_int,
		rstctrl_timer_i_type	=>	rstctrl_timer_i_type,
		rstctrl_timer_j	=>	rstctrl_timer_j_int,
		rstctrl_timer_j_type	=>	rstctrl_timer_j_type,
		rstctrl_tx_lcff_pll_lock_select	=>	rstctrl_tx_lcff_pll_lock_select,
		rstctrl_tx_lcff_pll_rstb_select	=>	rstctrl_tx_lcff_pll_rstb_select,
		rstctrl_tx_pcs_rst_n_inv	=>	rstctrl_tx_pcs_rst_n_inv,
		rstctrl_tx_pcs_rst_n_select	=>	rstctrl_tx_pcs_rst_n_select,
		rstctrl_tx_pma_rstb_inv	=>	rstctrl_tx_pma_rstb_inv,
		rstctrl_tx_pma_syncp_inv	=>	rstctrl_tx_pma_syncp_inv,
		rstctrl_tx_pma_syncp_select	=>	rstctrl_tx_pma_syncp_select,
		rx_ast_parity	=>	rx_ast_parity,
		rx_buffer_credit_alloc	=>	rx_buffer_credit_alloc,
		rx_buffer_fc_protect	=>	rx_buffer_fc_protect_int,
		rx_buffer_protect	=>	rx_buffer_protect_int,
		rx_cdc_almost_empty	=>	rx_cdc_almost_empty_int,
		rx_cdc_almost_full	=>	rx_cdc_almost_full_int,
		rx_cred_ctl_param	=>	rx_cred_ctl_param,
		rx_ei_l0s	=>	rx_ei_l0s,
		rx_l0s_count_idl	=>	rx_l0s_count_idl_int,
		rx_ptr0_nonposted_dpram_max	=>	rx_ptr0_nonposted_dpram_max_int,
		rx_ptr0_nonposted_dpram_min	=>	rx_ptr0_nonposted_dpram_min_int,
		rx_ptr0_posted_dpram_max	=>	rx_ptr0_posted_dpram_max_int,
		rx_ptr0_posted_dpram_min	=>	rx_ptr0_posted_dpram_min_int,
		rx_runt_patch_dis	=>	rx_runt_patch_dis,
		rx_sop_ctrl	=>	rx_sop_ctrl,
		rx_trunc_patch_dis	=>	rx_trunc_patch_dis,
		rx_use_prst	=>	rx_use_prst,
		rx_use_prst_ep	=>	rx_use_prst_ep,
		rxbuf_ecc_corr_mask_dis	=>	rxbuf_ecc_corr_mask_dis,
		rxdl_bad_sop_eop_filter_dis	=>	rxdl_bad_sop_eop_filter_dis,
		rxdl_bad_tlp_patch_dis	=>	rxdl_bad_tlp_patch_dis,
		rxdl_lcrc_patch_dis	=>	rxdl_lcrc_patch_dis,
		sameclock_nfts_count	=>	sameclock_nfts_count_int,
		sel_enable_pcs_rx_fifo_err	=>	sel_enable_pcs_rx_fifo_err,
		silicon_rev	=>	silicon_rev,
		sim_mode	=>	sim_mode,
		simple_ro_fifo_control_en	=>	simple_ro_fifo_control_en,
		single_rx_detect	=>	single_rx_detect,
		skp_os_gen3_count	=>	skp_os_gen3_count_int,
		skp_os_schedule_count	=>	skp_os_schedule_count_int,
		slot_number	=>	slot_number_int,
		slot_power_limit	=>	slot_power_limit_int,
		slot_power_scale	=>	slot_power_scale_int,
		slotclk_cfg	=>	slotclk_cfg,
		ssid	=>	ssid_int,
		ssvid	=>	ssvid_int,
		subsystem_device_id	=>	subsystem_device_id_int,
		subsystem_vendor_id	=>	subsystem_vendor_id_int,
		sup_mode	=>	sup_mode,
		surprise_down_error_support	=>	surprise_down_error_support,
		tl_cfg_div	=>	tl_cfg_div,
		tl_tx_check_parity_msg	=>	tl_tx_check_parity_msg,
		tph_completer	=>	tph_completer,
		tx_ast_parity	=>	tx_ast_parity,
		tx_cdc_almost_empty	=>	tx_cdc_almost_empty_int,
		tx_cdc_almost_full	=>	tx_cdc_almost_full_int,
		tx_sop_ctrl	=>	tx_sop_ctrl,
		tx_swing	=>	tx_swing_int,
		txdl_fair_arbiter_counter	=>	txdl_fair_arbiter_counter_int,
		txdl_fair_arbiter_en	=>	txdl_fair_arbiter_en,
		txrate_adv	=>	txrate_adv,
		uc_calibration_en	=>	uc_calibration_en,
		use_aer	=>	use_aer,
		use_crc_forwarding	=>	use_crc_forwarding,
		user_id	=>	user_id_int,
		vc0_clk_enable	=>	vc0_clk_enable,
		vc0_rx_buffer_memory_settings	=>	vc0_rx_buffer_memory_settings,
		vc0_rx_flow_ctrl_compl_data	=>	vc0_rx_flow_ctrl_compl_data_int,
		vc0_rx_flow_ctrl_compl_header	=>	vc0_rx_flow_ctrl_compl_header_int,
		vc0_rx_flow_ctrl_nonposted_data	=>	vc0_rx_flow_ctrl_nonposted_data_int,
		vc0_rx_flow_ctrl_nonposted_header	=>	vc0_rx_flow_ctrl_nonposted_header_int,
		vc0_rx_flow_ctrl_posted_data	=>	vc0_rx_flow_ctrl_posted_data_int,
		vc0_rx_flow_ctrl_posted_header	=>	vc0_rx_flow_ctrl_posted_header_int,
		vc1_clk_enable	=>	vc1_clk_enable,
		vc_arbitration	=>	vc_arbitration,
		vc_enable	=>	vc_enable,
		vendor_id	=>	vendor_id_int,
		vsec_cap	=>	vsec_cap_int,
		vsec_id	=>	vsec_id_int,
		wrong_device_id	=>	wrong_device_id
	)
	port map (
		-- Instance ports
		aer_msi_num	=>	aer_msi_num,
		app_int_err	=>	app_int_err,
		app_inta_sts	=>	app_inta_sts,
		app_msi_num	=>	app_msi_num,
		app_msi_req	=>	app_msi_req,
		app_msi_tc	=>	app_msi_tc,
		atpg_los_en_n	=>	atpg_los_en_n,
		avmm_address	=>	avmm_address,
		avmm_byte_en	=>	avmm_byte_en,
		avmm_clk	=>	avmm_clk,
		avmm_read	=>	avmm_read,
		avmm_rst_n	=>	avmm_rst_n,
		avmm_write	=>	avmm_write,
		avmm_writedata	=>	avmm_writedata,
		bist_scanen	=>	bist_scanen,
		bist_scanin	=>	bist_scanin,
		bisten_rcv_n	=>	bisten_rcv_n,
		bisten_rpl_n	=>	bisten_rpl_n,
		bistmode_n	=>	bistmode_n,
		cfg_link2csr_pld	=>	cfg_link2csr_pld,
		cfg_prmbus_pld	=>	cfg_prmbus_pld,
		chnl_cal_done0	=>	chnl_cal_done0,
		chnl_cal_done1	=>	chnl_cal_done1,
		chnl_cal_done2	=>	chnl_cal_done2,
		chnl_cal_done3	=>	chnl_cal_done3,
		chnl_cal_done4	=>	chnl_cal_done4,
		chnl_cal_done5	=>	chnl_cal_done5,
		chnl_cal_done6	=>	chnl_cal_done6,
		chnl_cal_done7	=>	chnl_cal_done7,
		core_clk_in	=>	core_clk_in,
		core_crst	=>	core_crst,
		core_por	=>	core_por,
		core_rst	=>	core_rst,
		core_srst	=>	core_srst,
		cpl_err	=>	cpl_err,
		cpl_pending	=>	cpl_pending,
		cseb_rddata	=>	cseb_rddata,
		cseb_rddata_parity	=>	cseb_rddata_parity,
		cseb_rdresponse	=>	cseb_rdresponse,
		cseb_waitrequest	=>	cseb_waitrequest,
		cseb_wrresp_valid	=>	cseb_wrresp_valid,
		cseb_wrresponse	=>	cseb_wrresponse,
		csr_cbdin	=>	csr_cbdin,
		csr_clk	=>	csr_clk,
		csr_din	=>	csr_din,
		csr_en	=>	csr_en,
		csr_enscan	=>	csr_enscan,
		csr_entest	=>	csr_entest,
		csr_in	=>	csr_in,
		csr_load_csr	=>	csr_load_csr,
		csr_pipe_in	=>	csr_pipe_in,
		csr_seg	=>	csr_seg,
		csr_tcsrin	=>	csr_tcsrin,
		csr_tverify	=>	csr_tverify,
		cvp_config_done	=>	cvp_config_done,
		cvp_config_error	=>	cvp_config_error,
		cvp_config_ready	=>	cvp_config_ready,
		cvp_en	=>	cvp_en,
		egress_blk_err	=>	egress_blk_err,
		entest	=>	entest,
		flr_reset	=>	flr_reset,
		force_tx_eidle	=>	force_tx_eidle,
		fref_clk0	=>	fref_clk0,
		fref_clk1	=>	fref_clk1,
		fref_clk2	=>	fref_clk2,
		fref_clk3	=>	fref_clk3,
		fref_clk4	=>	fref_clk4,
		fref_clk5	=>	fref_clk5,
		fref_clk6	=>	fref_clk6,
		fref_clk7	=>	fref_clk7,
		frzlogic	=>	frzlogic,
		frzreg	=>	frzreg,
		hold_ltssm_rec	=>	hold_ltssm_rec,
		hpg_ctrler	=>	hpg_ctrler,
		iocsrrdy_dly	=>	iocsrrdy_dly,
		lmi_addr	=>	lmi_addr,
		lmi_din	=>	lmi_din,
		lmi_rden	=>	lmi_rden,
		lmi_wren	=>	lmi_wren,
		m10k_select	=>	m10k_select,
		mask_tx_pll_lock0	=>	mask_tx_pll_lock0,
		mask_tx_pll_lock1	=>	mask_tx_pll_lock1,
		mask_tx_pll_lock2	=>	mask_tx_pll_lock2,
		mask_tx_pll_lock3	=>	mask_tx_pll_lock3,
		mask_tx_pll_lock4	=>	mask_tx_pll_lock4,
		mask_tx_pll_lock5	=>	mask_tx_pll_lock5,
		mask_tx_pll_lock6	=>	mask_tx_pll_lock6,
		mask_tx_pll_lock7	=>	mask_tx_pll_lock7,
		mem_hip_test_enable	=>	mem_hip_test_enable,
		mem_regscanen_n	=>	mem_regscanen_n,
		mem_rscin_rcv_bot	=>	mem_rscin_rcv_bot,
		mem_rscin_rcv_top	=>	mem_rscin_rcv_top,
		mem_rscin_rtry	=>	mem_rscin_rtry,
		nfrzdrv	=>	nfrzdrv,
		npor	=>	npor,
		pclk_central	=>	pclk_central,
		pclk_ch0	=>	pclk_ch0,
		pclk_ch1	=>	pclk_ch1,
		pex_msi_num	=>	pex_msi_num,
		phy_rst	=>	phy_rst,
		phy_srst	=>	phy_srst,
		phystatus0	=>	phystatus0,
		phystatus1	=>	phystatus1,
		phystatus2	=>	phystatus2,
		phystatus3	=>	phystatus3,
		phystatus4	=>	phystatus4,
		phystatus5	=>	phystatus5,
		phystatus6	=>	phystatus6,
		phystatus7	=>	phystatus7,
		pin_perst_n	=>	pin_perst_n,
		pld_clk	=>	pld_clk,
		pld_clrhip_n	=>	pld_clrhip_n,
		pld_clrpcship_n	=>	pld_clrpcship_n,
		pld_clrpmapcship_n	=>	pld_clrpmapcship_n,
		pld_core_ready	=>	pld_core_ready,
		pld_gp_status	=>	pld_gp_status,
		pld_perst_n	=>	pld_perst_n,
		pll_cal_done0	=>	pll_cal_done0,
		pll_cal_done1	=>	pll_cal_done1,
		pll_cal_done2	=>	pll_cal_done2,
		pll_cal_done3	=>	pll_cal_done3,
		pll_cal_done4	=>	pll_cal_done4,
		pll_cal_done5	=>	pll_cal_done5,
		pll_cal_done6	=>	pll_cal_done6,
		pll_cal_done7	=>	pll_cal_done7,
		pll_fixed_clk_central	=>	pll_fixed_clk_central,
		pll_fixed_clk_ch0	=>	pll_fixed_clk_ch0,
		pll_fixed_clk_ch1	=>	pll_fixed_clk_ch1,
		plniotri	=>	plniotri,
		pm_auxpwr	=>	pm_auxpwr,
		pm_data	=>	pm_data,
		pm_event	=>	pm_event,
		pm_exit_d0_ack	=>	pm_exit_d0_ack,
		pme_to_cr	=>	pme_to_cr,
		reserved_clk_in	=>	reserved_clk_in,
		reserved_in	=>	reserved_in,
		rx_cred_ctl	=>	rx_cred_ctl,
		rx_pll_freq_lock0	=>	rx_pll_freq_lock0,
		rx_pll_freq_lock1	=>	rx_pll_freq_lock1,
		rx_pll_freq_lock2	=>	rx_pll_freq_lock2,
		rx_pll_freq_lock3	=>	rx_pll_freq_lock3,
		rx_pll_freq_lock4	=>	rx_pll_freq_lock4,
		rx_pll_freq_lock5	=>	rx_pll_freq_lock5,
		rx_pll_freq_lock6	=>	rx_pll_freq_lock6,
		rx_pll_freq_lock7	=>	rx_pll_freq_lock7,
		rx_pll_phase_lock0	=>	rx_pll_phase_lock0,
		rx_pll_phase_lock1	=>	rx_pll_phase_lock1,
		rx_pll_phase_lock2	=>	rx_pll_phase_lock2,
		rx_pll_phase_lock3	=>	rx_pll_phase_lock3,
		rx_pll_phase_lock4	=>	rx_pll_phase_lock4,
		rx_pll_phase_lock5	=>	rx_pll_phase_lock5,
		rx_pll_phase_lock6	=>	rx_pll_phase_lock6,
		rx_pll_phase_lock7	=>	rx_pll_phase_lock7,
		rx_st_mask	=>	rx_st_mask,
		rx_st_ready	=>	rx_st_ready,
		rxblkst0	=>	rxblkst0,
		rxblkst1	=>	rxblkst1,
		rxblkst2	=>	rxblkst2,
		rxblkst3	=>	rxblkst3,
		rxblkst4	=>	rxblkst4,
		rxblkst5	=>	rxblkst5,
		rxblkst6	=>	rxblkst6,
		rxblkst7	=>	rxblkst7,
		rxdata0	=>	rxdata0,
		rxdata1	=>	rxdata1,
		rxdata2	=>	rxdata2,
		rxdata3	=>	rxdata3,
		rxdata4	=>	rxdata4,
		rxdata5	=>	rxdata5,
		rxdata6	=>	rxdata6,
		rxdata7	=>	rxdata7,
		rxdatak0	=>	rxdatak0,
		rxdatak1	=>	rxdatak1,
		rxdatak2	=>	rxdatak2,
		rxdatak3	=>	rxdatak3,
		rxdatak4	=>	rxdatak4,
		rxdatak5	=>	rxdatak5,
		rxdatak6	=>	rxdatak6,
		rxdatak7	=>	rxdatak7,
		rxdataskip0	=>	rxdataskip0,
		rxdataskip1	=>	rxdataskip1,
		rxdataskip2	=>	rxdataskip2,
		rxdataskip3	=>	rxdataskip3,
		rxdataskip4	=>	rxdataskip4,
		rxdataskip5	=>	rxdataskip5,
		rxdataskip6	=>	rxdataskip6,
		rxdataskip7	=>	rxdataskip7,
		rxelecidle0	=>	rxelecidle0,
		rxelecidle1	=>	rxelecidle1,
		rxelecidle2	=>	rxelecidle2,
		rxelecidle3	=>	rxelecidle3,
		rxelecidle4	=>	rxelecidle4,
		rxelecidle5	=>	rxelecidle5,
		rxelecidle6	=>	rxelecidle6,
		rxelecidle7	=>	rxelecidle7,
		rxfreqlocked0	=>	rxfreqlocked0,
		rxfreqlocked1	=>	rxfreqlocked1,
		rxfreqlocked2	=>	rxfreqlocked2,
		rxfreqlocked3	=>	rxfreqlocked3,
		rxfreqlocked4	=>	rxfreqlocked4,
		rxfreqlocked5	=>	rxfreqlocked5,
		rxfreqlocked6	=>	rxfreqlocked6,
		rxfreqlocked7	=>	rxfreqlocked7,
		rxstatus0	=>	rxstatus0,
		rxstatus1	=>	rxstatus1,
		rxstatus2	=>	rxstatus2,
		rxstatus3	=>	rxstatus3,
		rxstatus4	=>	rxstatus4,
		rxstatus5	=>	rxstatus5,
		rxstatus6	=>	rxstatus6,
		rxstatus7	=>	rxstatus7,
		rxsynchd0	=>	rxsynchd0,
		rxsynchd1	=>	rxsynchd1,
		rxsynchd2	=>	rxsynchd2,
		rxsynchd3	=>	rxsynchd3,
		rxsynchd4	=>	rxsynchd4,
		rxsynchd5	=>	rxsynchd5,
		rxsynchd6	=>	rxsynchd6,
		rxsynchd7	=>	rxsynchd7,
		rxvalid0	=>	rxvalid0,
		rxvalid1	=>	rxvalid1,
		rxvalid2	=>	rxvalid2,
		rxvalid3	=>	rxvalid3,
		rxvalid4	=>	rxvalid4,
		rxvalid5	=>	rxvalid5,
		rxvalid6	=>	rxvalid6,
		rxvalid7	=>	rxvalid7,
		scan_mode_n	=>	scan_mode_n,
		scan_shift_n	=>	scan_shift_n,
		sw_ctmod	=>	sw_ctmod,
		swdn_in	=>	swdn_in,
		swup_in	=>	swup_in,
		test_in_1_hip	=>	test_in_1_hip,
		test_in_hip	=>	test_in_hip,
		test_pl_dbg_eqin	=>	test_pl_dbg_eqin,
		tx_cred_cons_select	=>	tx_cred_cons_select,
		tx_cred_fc_sel	=>	tx_cred_fc_sel,
		tx_lcff_pll_lock0	=>	tx_lcff_pll_lock0,
		tx_lcff_pll_lock1	=>	tx_lcff_pll_lock1,
		tx_lcff_pll_lock2	=>	tx_lcff_pll_lock2,
		tx_lcff_pll_lock3	=>	tx_lcff_pll_lock3,
		tx_lcff_pll_lock4	=>	tx_lcff_pll_lock4,
		tx_lcff_pll_lock5	=>	tx_lcff_pll_lock5,
		tx_lcff_pll_lock6	=>	tx_lcff_pll_lock6,
		tx_lcff_pll_lock7	=>	tx_lcff_pll_lock7,
		tx_st_data	=>	tx_st_data,
		tx_st_empty	=>	tx_st_empty,
		tx_st_eop	=>	tx_st_eop,
		tx_st_err	=>	tx_st_err,
		tx_st_parity	=>	tx_st_parity,
		tx_st_sop	=>	tx_st_sop,
		tx_st_valid	=>	tx_st_valid,
		user_mode	=>	user_mode,
		sta_hd_altpe3_hip_core_top_hd_altpe3_hip_core_u_clkmux_core_clk_cnt_reg_0_0_Q	=>	sta_hd_altpe3_hip_core_top_hd_altpe3_hip_core_u_clkmux_core_clk_cnt_reg_0_0_Q,
		sta_hd_altpe3_hip_core_top_hd_altpe3_hip_core_u_clkmux_core_clk_cnt_reg_1_0_Q	=>	sta_hd_altpe3_hip_core_top_hd_altpe3_hip_core_u_clkmux_core_clk_cnt_reg_1_0_Q,
		sta_hd_altpe3_hip_core_top_hd_altpe3_hip_core_u_clkmux_core_clk_cnt_reg_2_0_Q	=>	sta_hd_altpe3_hip_core_top_hd_altpe3_hip_core_u_clkmux_core_clk_cnt_reg_2_0_Q,
		app_inta_ack	=>	app_inta_ack,
		app_msi_ack	=>	app_msi_ack,
		avmm_readdata	=>	avmm_readdata,
		cfg_par_err	=>	cfg_par_err,
		core_clk_out	=>	core_clk_out,
		cseb_addr	=>	cseb_addr,
		cseb_addr_parity	=>	cseb_addr_parity,
		cseb_be	=>	cseb_be,
		cseb_is_shadow	=>	cseb_is_shadow,
		cseb_rden	=>	cseb_rden,
		cseb_wrdata	=>	cseb_wrdata,
		cseb_wrdata_parity	=>	cseb_wrdata_parity,
		cseb_wren	=>	cseb_wren,
		cseb_wrresp_req	=>	cseb_wrresp_req,
		csr_dout	=>	csr_dout,
		csr_out	=>	csr_out,
		csr_pipe_out	=>	csr_pipe_out,
		current_coeff0	=>	current_coeff0,
		current_coeff1	=>	current_coeff1,
		current_coeff2	=>	current_coeff2,
		current_coeff3	=>	current_coeff3,
		current_coeff4	=>	current_coeff4,
		current_coeff5	=>	current_coeff5,
		current_coeff6	=>	current_coeff6,
		current_coeff7	=>	current_coeff7,
		current_rxpreset0	=>	current_rxpreset0,
		current_rxpreset1	=>	current_rxpreset1,
		current_rxpreset2	=>	current_rxpreset2,
		current_rxpreset3	=>	current_rxpreset3,
		current_rxpreset4	=>	current_rxpreset4,
		current_rxpreset5	=>	current_rxpreset5,
		current_rxpreset6	=>	current_rxpreset6,
		current_rxpreset7	=>	current_rxpreset7,
		current_speed	=>	current_speed,
		cvp_clk	=>	cvp_clk,
		cvp_config	=>	cvp_config,
		cvp_data	=>	cvp_data,
		cvp_full_config	=>	cvp_full_config,
		cvp_start_xfer	=>	cvp_start_xfer,
		dl_up	=>	dl_up,
		dlup_exit	=>	dlup_exit,
		eidle_infer_sel0	=>	eidle_infer_sel0,
		eidle_infer_sel1	=>	eidle_infer_sel1,
		eidle_infer_sel2	=>	eidle_infer_sel2,
		eidle_infer_sel3	=>	eidle_infer_sel3,
		eidle_infer_sel4	=>	eidle_infer_sel4,
		eidle_infer_sel5	=>	eidle_infer_sel5,
		eidle_infer_sel6	=>	eidle_infer_sel6,
		eidle_infer_sel7	=>	eidle_infer_sel7,
		ev_128ns	=>	ev_128ns,
		ev_1us	=>	ev_1us,
		flr_sts	=>	flr_sts,
		g3_rx_pcs_rst_n0	=>	g3_rx_pcs_rst_n0,
		g3_rx_pcs_rst_n1	=>	g3_rx_pcs_rst_n1,
		g3_rx_pcs_rst_n2	=>	g3_rx_pcs_rst_n2,
		g3_rx_pcs_rst_n3	=>	g3_rx_pcs_rst_n3,
		g3_rx_pcs_rst_n4	=>	g3_rx_pcs_rst_n4,
		g3_rx_pcs_rst_n5	=>	g3_rx_pcs_rst_n5,
		g3_rx_pcs_rst_n6	=>	g3_rx_pcs_rst_n6,
		g3_rx_pcs_rst_n7	=>	g3_rx_pcs_rst_n7,
		g3_tx_pcs_rst_n0	=>	g3_tx_pcs_rst_n0,
		g3_tx_pcs_rst_n1	=>	g3_tx_pcs_rst_n1,
		g3_tx_pcs_rst_n2	=>	g3_tx_pcs_rst_n2,
		g3_tx_pcs_rst_n3	=>	g3_tx_pcs_rst_n3,
		g3_tx_pcs_rst_n4	=>	g3_tx_pcs_rst_n4,
		g3_tx_pcs_rst_n5	=>	g3_tx_pcs_rst_n5,
		g3_tx_pcs_rst_n6	=>	g3_tx_pcs_rst_n6,
		g3_tx_pcs_rst_n7	=>	g3_tx_pcs_rst_n7,
		hotrst_exit	=>	hotrst_exit,
		int_status	=>	int_status,
		k_hip_pcs_chnl_en	=>	k_hip_pcs_chnl_en,
		k_hrc_chnl_en	=>	k_hrc_chnl_en,
		k_hrc_chnl_txpll_master_cgb_rst_en	=>	k_hrc_chnl_txpll_master_cgb_rst_en,
		k_hrc_chnl_txpll_rst_en	=>	k_hrc_chnl_txpll_rst_en,
		l2_exit	=>	l2_exit,
		lane_act	=>	lane_act,
		lmi_ack	=>	lmi_ack,
		lmi_dout	=>	lmi_dout,
		ltssm_state	=>	ltssm_state,
		mem_rscout_rcv_bot	=>	mem_rscout_rcv_bot,
		mem_rscout_rcv_top	=>	mem_rscout_rcv_top,
		mem_rscout_rtry	=>	mem_rscout_rtry,
		pld_clk_in_use	=>	pld_clk_in_use,
		pld_gp_ctrl	=>	pld_gp_ctrl,
		pm_exit_d0_req	=>	pm_exit_d0_req,
		pme_to_sr	=>	pme_to_sr,
		powerdown0	=>	powerdown0,
		powerdown1	=>	powerdown1,
		powerdown2	=>	powerdown2,
		powerdown3	=>	powerdown3,
		powerdown4	=>	powerdown4,
		powerdown5	=>	powerdown5,
		powerdown6	=>	powerdown6,
		powerdown7	=>	powerdown7,
		r2c_unc_ecc	=>	r2c_unc_ecc,
		rate0	=>	rate0,
		rate1	=>	rate1,
		rate2	=>	rate2,
		rate3	=>	rate3,
		rate4	=>	rate4,
		rate5	=>	rate5,
		rate6	=>	rate6,
		rate7	=>	rate7,
		rate_ctrl	=>	rate_ctrl,
		reserved_clk_out	=>	reserved_clk_out,
		reserved_out	=>	reserved_out,
		reset_status	=>	reset_status,
		retry_corr_ecc	=>	retry_corr_ecc,
		retry_unc_ecc	=>	retry_unc_ecc,
		rx_corr_ecc	=>	rx_corr_ecc,
		rx_cred_status	=>	rx_cred_status,
		rx_par_err	=>	rx_par_err,
		rx_pcs_rst_n0	=>	rx_pcs_rst_n0,
		rx_pcs_rst_n1	=>	rx_pcs_rst_n1,
		rx_pcs_rst_n2	=>	rx_pcs_rst_n2,
		rx_pcs_rst_n3	=>	rx_pcs_rst_n3,
		rx_pcs_rst_n4	=>	rx_pcs_rst_n4,
		rx_pcs_rst_n5	=>	rx_pcs_rst_n5,
		rx_pcs_rst_n6	=>	rx_pcs_rst_n6,
		rx_pcs_rst_n7	=>	rx_pcs_rst_n7,
		rx_pma_rstb0	=>	rx_pma_rstb0,
		rx_pma_rstb1	=>	rx_pma_rstb1,
		rx_pma_rstb2	=>	rx_pma_rstb2,
		rx_pma_rstb3	=>	rx_pma_rstb3,
		rx_pma_rstb4	=>	rx_pma_rstb4,
		rx_pma_rstb5	=>	rx_pma_rstb5,
		rx_pma_rstb6	=>	rx_pma_rstb6,
		rx_pma_rstb7	=>	rx_pma_rstb7,
		rx_st_bardec1	=>	rx_st_bardec1,
		rx_st_bardec2	=>	rx_st_bardec2,
		rx_st_be	=>	rx_st_be,
		rx_st_data	=>	rx_st_data,
		rx_st_empty	=>	rx_st_empty,
		rx_st_eop	=>	rx_st_eop,
		rx_st_err	=>	rx_st_err,
		rx_st_parity	=>	rx_st_parity,
		rx_st_sop	=>	rx_st_sop,
		rx_st_valid	=>	rx_st_valid,
		rxfc_cplbuf_ovf	=>	rxfc_cplbuf_ovf,
		rxfc_cplovf_tag	=>	rxfc_cplovf_tag,
		rxpolarity0	=>	rxpolarity0,
		rxpolarity1	=>	rxpolarity1,
		rxpolarity2	=>	rxpolarity2,
		rxpolarity3	=>	rxpolarity3,
		rxpolarity4	=>	rxpolarity4,
		rxpolarity5	=>	rxpolarity5,
		rxpolarity6	=>	rxpolarity6,
		rxpolarity7	=>	rxpolarity7,
		serr_out	=>	serr_out,
		swdn_out	=>	swdn_out,
		swup_out	=>	swup_out,
		test_fref_clk	=>	test_fref_clk,
		test_out_1_hip	=>	test_out_1_hip,
		test_out_hip	=>	test_out_hip,
		tl_cfg_add	=>	tl_cfg_add,
		tl_cfg_ctl	=>	tl_cfg_ctl,
		tl_cfg_sts	=>	tl_cfg_sts,
		tl_cfg_sts_wr	=>	tl_cfg_sts_wr,
		tx_cred_data_fc	=>	tx_cred_data_fc,
		tx_cred_fc_hip_cons	=>	tx_cred_fc_hip_cons,
		tx_cred_fc_infinite	=>	tx_cred_fc_infinite,
		tx_cred_hdr_fc	=>	tx_cred_hdr_fc,
		tx_deemph0	=>	tx_deemph0,
		tx_deemph1	=>	tx_deemph1,
		tx_deemph2	=>	tx_deemph2,
		tx_deemph3	=>	tx_deemph3,
		tx_deemph4	=>	tx_deemph4,
		tx_deemph5	=>	tx_deemph5,
		tx_deemph6	=>	tx_deemph6,
		tx_deemph7	=>	tx_deemph7,
		tx_lcff_pll_rstb0	=>	tx_lcff_pll_rstb0,
		tx_lcff_pll_rstb1	=>	tx_lcff_pll_rstb1,
		tx_lcff_pll_rstb2	=>	tx_lcff_pll_rstb2,
		tx_lcff_pll_rstb3	=>	tx_lcff_pll_rstb3,
		tx_lcff_pll_rstb4	=>	tx_lcff_pll_rstb4,
		tx_lcff_pll_rstb5	=>	tx_lcff_pll_rstb5,
		tx_lcff_pll_rstb6	=>	tx_lcff_pll_rstb6,
		tx_lcff_pll_rstb7	=>	tx_lcff_pll_rstb7,
		tx_margin0	=>	tx_margin0,
		tx_margin1	=>	tx_margin1,
		tx_margin2	=>	tx_margin2,
		tx_margin3	=>	tx_margin3,
		tx_margin4	=>	tx_margin4,
		tx_margin5	=>	tx_margin5,
		tx_margin6	=>	tx_margin6,
		tx_margin7	=>	tx_margin7,
		tx_par_err	=>	tx_par_err,
		tx_pcs_rst_n0	=>	tx_pcs_rst_n0,
		tx_pcs_rst_n1	=>	tx_pcs_rst_n1,
		tx_pcs_rst_n2	=>	tx_pcs_rst_n2,
		tx_pcs_rst_n3	=>	tx_pcs_rst_n3,
		tx_pcs_rst_n4	=>	tx_pcs_rst_n4,
		tx_pcs_rst_n5	=>	tx_pcs_rst_n5,
		tx_pcs_rst_n6	=>	tx_pcs_rst_n6,
		tx_pcs_rst_n7	=>	tx_pcs_rst_n7,
		tx_pma_syncp0	=>	tx_pma_syncp0,
		tx_pma_syncp1	=>	tx_pma_syncp1,
		tx_pma_syncp2	=>	tx_pma_syncp2,
		tx_pma_syncp3	=>	tx_pma_syncp3,
		tx_pma_syncp4	=>	tx_pma_syncp4,
		tx_pma_syncp5	=>	tx_pma_syncp5,
		tx_pma_syncp6	=>	tx_pma_syncp6,
		tx_pma_syncp7	=>	tx_pma_syncp7,
		tx_st_ready	=>	tx_st_ready,
		txblkst0	=>	txblkst0,
		txblkst1	=>	txblkst1,
		txblkst2	=>	txblkst2,
		txblkst3	=>	txblkst3,
		txblkst4	=>	txblkst4,
		txblkst5	=>	txblkst5,
		txblkst6	=>	txblkst6,
		txblkst7	=>	txblkst7,
		txcompl0	=>	txcompl0,
		txcompl1	=>	txcompl1,
		txcompl2	=>	txcompl2,
		txcompl3	=>	txcompl3,
		txcompl4	=>	txcompl4,
		txcompl5	=>	txcompl5,
		txcompl6	=>	txcompl6,
		txcompl7	=>	txcompl7,
		txdata0	=>	txdata0,
		txdata1	=>	txdata1,
		txdata2	=>	txdata2,
		txdata3	=>	txdata3,
		txdata4	=>	txdata4,
		txdata5	=>	txdata5,
		txdata6	=>	txdata6,
		txdata7	=>	txdata7,
		txdatak0	=>	txdatak0,
		txdatak1	=>	txdatak1,
		txdatak2	=>	txdatak2,
		txdatak3	=>	txdatak3,
		txdatak4	=>	txdatak4,
		txdatak5	=>	txdatak5,
		txdatak6	=>	txdatak6,
		txdatak7	=>	txdatak7,
		txdataskip0	=>	txdataskip0,
		txdataskip1	=>	txdataskip1,
		txdataskip2	=>	txdataskip2,
		txdataskip3	=>	txdataskip3,
		txdataskip4	=>	txdataskip4,
		txdataskip5	=>	txdataskip5,
		txdataskip6	=>	txdataskip6,
		txdataskip7	=>	txdataskip7,
		txdetectrx0	=>	txdetectrx0,
		txdetectrx1	=>	txdetectrx1,
		txdetectrx2	=>	txdetectrx2,
		txdetectrx3	=>	txdetectrx3,
		txdetectrx4	=>	txdetectrx4,
		txdetectrx5	=>	txdetectrx5,
		txdetectrx6	=>	txdetectrx6,
		txdetectrx7	=>	txdetectrx7,
		txelecidle0	=>	txelecidle0,
		txelecidle1	=>	txelecidle1,
		txelecidle2	=>	txelecidle2,
		txelecidle3	=>	txelecidle3,
		txelecidle4	=>	txelecidle4,
		txelecidle5	=>	txelecidle5,
		txelecidle6	=>	txelecidle6,
		txelecidle7	=>	txelecidle7,
		txst_prot_err	=>	txst_prot_err,
		txswing0	=>	txswing0,
		txswing1	=>	txswing1,
		txswing2	=>	txswing2,
		txswing3	=>	txswing3,
		txswing4	=>	txswing4,
		txswing5	=>	txswing5,
		txswing6	=>	txswing6,
		txswing7	=>	txswing7,
		txsynchd0	=>	txsynchd0,
		txsynchd1	=>	txsynchd1,
		txsynchd2	=>	txsynchd2,
		txsynchd3	=>	txsynchd3,
		txsynchd4	=>	txsynchd4,
		txsynchd5	=>	txsynchd5,
		txsynchd6	=>	txsynchd6,
		txsynchd7	=>	txsynchd7,
		wake_oen	=>	wake_oen
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_krfec_rx_pcs	is
	generic (
		-- Entity parameters
		blksync_cor_en	:	string	:=	"detect";
		bypass_gb	:	string	:=	"bypass_dis";
		clr_ctrl	:	string	:=	"both_enabled";
		ctrl_bit_reverse	:	string	:=	"ctrl_bit_reverse_dis";
		data_bit_reverse	:	string	:=	"data_bit_reverse_dis";
		dv_start	:	string	:=	"with_blklock";
		err_mark_type	:	string	:=	"err_mark_10g";
		error_marking_en	:	string	:=	"err_mark_dis";
		low_latency_en	:	string	:=	"disable";
		lpbk_mode	:	string	:=	"lpbk_dis";
		parity_invalid_enum	:	bit_vector	:=	B"00001000";
		parity_valid_num	:	bit_vector	:=	B"0100";
		pipeln_blksync	:	string	:=	"enable";
		pipeln_descrm	:	string	:=	"enable";
		pipeln_errcorrect	:	string	:=	"enable";
		pipeln_errtrap_ind	:	string	:=	"enable";
		pipeln_errtrap_lfsr	:	string	:=	"enable";
		pipeln_errtrap_loc	:	string	:=	"enable";
		pipeln_errtrap_pat	:	string	:=	"enable";
		pipeln_gearbox	:	string	:=	"enable";
		pipeln_syndrm	:	string	:=	"enable";
		pipeln_trans_dec	:	string	:=	"enable";
		prot_mode	:	string	:=	"disable_mode";
		receive_order	:	string	:=	"receive_lsb";
		reconfig_settings	:	string	:=	"{}";
		rx_testbus_sel	:	string	:=	"overall";
		signal_ok_en	:	string	:=	"sig_ok_dis";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		rx_clr_counters	:	in	std_logic	:=	'0';
		rx_data_in	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		rx_krfec_clk	:	in	std_logic	:=	'0';
		rx_master_clk	:	in	std_logic	:=	'0';
		rx_master_clk_rst_n	:	in	std_logic	:=	'0';
		rx_signal_ok_in	:	in	std_logic	:=	'0';
		scan_mode_n	:	in	std_logic	:=	'0';
		scan_rst_n	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_blk_lock_krfec_reg	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_blk_lock_krfec_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_diag_data_status_krfec_reg	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_diag_data_status_krfec_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_frame_krfec_reg	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_frame_krfec_txclk_reg	:	out	std_logic	:=	'0';
		rx_block_lock	:	out	std_logic	:=	'0';
		rx_control_out	:	out	std_logic_vector(9 downto 0)	:=	"0000000000";
		rx_data_out	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		rx_data_status	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rx_data_valid_out	:	out	std_logic	:=	'0';
		rx_frame	:	out	std_logic	:=	'0';
		rx_signal_ok_out	:	out	std_logic	:=	'0';
		rx_test_data	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000"
	);
end twentynm_hssi_krfec_rx_pcs;

architecture behavior of twentynm_hssi_krfec_rx_pcs	is

constant parity_invalid_enum_int	:	integer	:=	bin2int(parity_invalid_enum);
constant parity_valid_num_int	:	integer	:=	bin2int(parity_valid_num);



component	twentynm_hssi_krfec_rx_pcs_encrypted
	generic (
		-- Architecture parameters
		blksync_cor_en	:	string	:=	"detect";
		bypass_gb	:	string	:=	"bypass_dis";
		clr_ctrl	:	string	:=	"both_enabled";
		ctrl_bit_reverse	:	string	:=	"ctrl_bit_reverse_dis";
		data_bit_reverse	:	string	:=	"data_bit_reverse_dis";
		dv_start	:	string	:=	"with_blklock";
		err_mark_type	:	string	:=	"err_mark_10g";
		error_marking_en	:	string	:=	"err_mark_dis";
		low_latency_en	:	string	:=	"disable";
		lpbk_mode	:	string	:=	"lpbk_dis";
		parity_invalid_enum	:	integer	:=	8;
		parity_valid_num	:	integer	:=	4;
		pipeln_blksync	:	string	:=	"enable";
		pipeln_descrm	:	string	:=	"enable";
		pipeln_errcorrect	:	string	:=	"enable";
		pipeln_errtrap_ind	:	string	:=	"enable";
		pipeln_errtrap_lfsr	:	string	:=	"enable";
		pipeln_errtrap_loc	:	string	:=	"enable";
		pipeln_errtrap_pat	:	string	:=	"enable";
		pipeln_gearbox	:	string	:=	"enable";
		pipeln_syndrm	:	string	:=	"enable";
		pipeln_trans_dec	:	string	:=	"enable";
		prot_mode	:	string	:=	"disable_mode";
		receive_order	:	string	:=	"receive_lsb";
		reconfig_settings	:	string	:=	"{}";
		rx_testbus_sel	:	string	:=	"overall";
		signal_ok_en	:	string	:=	"sig_ok_dis";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode"
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		rx_clr_counters	:	in	std_logic	:=	'0';
		rx_data_in	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		rx_krfec_clk	:	in	std_logic	:=	'0';
		rx_master_clk	:	in	std_logic	:=	'0';
		rx_master_clk_rst_n	:	in	std_logic	:=	'0';
		rx_signal_ok_in	:	in	std_logic	:=	'0';
		scan_mode_n	:	in	std_logic	:=	'0';
		scan_rst_n	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_blk_lock_krfec_reg	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_blk_lock_krfec_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_diag_data_status_krfec_reg	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_diag_data_status_krfec_txclk_reg	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_frame_krfec_reg	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_frame_krfec_txclk_reg	:	out	std_logic	:=	'0';
		rx_block_lock	:	out	std_logic	:=	'0';
		rx_control_out	:	out	std_logic_vector(9 downto 0)	:=	"0000000000";
		rx_data_out	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		rx_data_status	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rx_data_valid_out	:	out	std_logic	:=	'0';
		rx_frame	:	out	std_logic	:=	'0';
		rx_signal_ok_out	:	out	std_logic	:=	'0';
		rx_test_data	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000"
	);
end component;

begin



inst : twentynm_hssi_krfec_rx_pcs_encrypted
	generic map (
		-- Instance parameters
		blksync_cor_en	=>	blksync_cor_en,
		bypass_gb	=>	bypass_gb,
		clr_ctrl	=>	clr_ctrl,
		ctrl_bit_reverse	=>	ctrl_bit_reverse,
		data_bit_reverse	=>	data_bit_reverse,
		dv_start	=>	dv_start,
		err_mark_type	=>	err_mark_type,
		error_marking_en	=>	error_marking_en,
		low_latency_en	=>	low_latency_en,
		lpbk_mode	=>	lpbk_mode,
		parity_invalid_enum	=>	parity_invalid_enum_int,
		parity_valid_num	=>	parity_valid_num_int,
		pipeln_blksync	=>	pipeln_blksync,
		pipeln_descrm	=>	pipeln_descrm,
		pipeln_errcorrect	=>	pipeln_errcorrect,
		pipeln_errtrap_ind	=>	pipeln_errtrap_ind,
		pipeln_errtrap_lfsr	=>	pipeln_errtrap_lfsr,
		pipeln_errtrap_loc	=>	pipeln_errtrap_loc,
		pipeln_errtrap_pat	=>	pipeln_errtrap_pat,
		pipeln_gearbox	=>	pipeln_gearbox,
		pipeln_syndrm	=>	pipeln_syndrm,
		pipeln_trans_dec	=>	pipeln_trans_dec,
		prot_mode	=>	prot_mode,
		receive_order	=>	receive_order,
		reconfig_settings	=>	reconfig_settings,
		rx_testbus_sel	=>	rx_testbus_sel,
		signal_ok_en	=>	signal_ok_en,
		silicon_rev	=>	silicon_rev,
		sup_mode	=>	sup_mode
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		rx_clr_counters	=>	rx_clr_counters,
		rx_data_in	=>	rx_data_in,
		rx_krfec_clk	=>	rx_krfec_clk,
		rx_master_clk	=>	rx_master_clk,
		rx_master_clk_rst_n	=>	rx_master_clk_rst_n,
		rx_signal_ok_in	=>	rx_signal_ok_in,
		scan_mode_n	=>	scan_mode_n,
		scan_rst_n	=>	scan_rst_n,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		pld_10g_krfec_rx_blk_lock_krfec_reg	=>	pld_10g_krfec_rx_blk_lock_krfec_reg,
		pld_10g_krfec_rx_blk_lock_krfec_txclk_reg	=>	pld_10g_krfec_rx_blk_lock_krfec_txclk_reg,
		pld_10g_krfec_rx_diag_data_status_krfec_reg	=>	pld_10g_krfec_rx_diag_data_status_krfec_reg,
		pld_10g_krfec_rx_diag_data_status_krfec_txclk_reg	=>	pld_10g_krfec_rx_diag_data_status_krfec_txclk_reg,
		pld_10g_krfec_rx_frame_krfec_reg	=>	pld_10g_krfec_rx_frame_krfec_reg,
		pld_10g_krfec_rx_frame_krfec_txclk_reg	=>	pld_10g_krfec_rx_frame_krfec_txclk_reg,
		rx_block_lock	=>	rx_block_lock,
		rx_control_out	=>	rx_control_out,
		rx_data_out	=>	rx_data_out,
		rx_data_status	=>	rx_data_status,
		rx_data_valid_out	=>	rx_data_valid_out,
		rx_frame	=>	rx_frame,
		rx_signal_ok_out	=>	rx_signal_ok_out,
		rx_test_data	=>	rx_test_data
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_krfec_tx_pcs	is
	generic (
		-- Entity parameters
		burst_err	:	string	:=	"burst_err_dis";
		burst_err_len	:	string	:=	"burst_err_len1";
		ctrl_bit_reverse	:	string	:=	"ctrl_bit_reverse_dis";
		data_bit_reverse	:	string	:=	"data_bit_reverse_dis";
		enc_frame_query	:	string	:=	"enc_query_dis";
		low_latency_en	:	string	:=	"disable";
		pipeln_encoder	:	string	:=	"enable";
		pipeln_scrambler	:	string	:=	"enable";
		prot_mode	:	string	:=	"disable_mode";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode";
		transcode_err	:	string	:=	"trans_err_dis";
		transmit_order	:	string	:=	"transmit_lsb";
		tx_testbus_sel	:	string	:=	"overall"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		tx_control_in	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		tx_data_in	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		tx_data_valid_in	:	in	std_logic	:=	'0';
		tx_krfec_clk	:	in	std_logic	:=	'0';
		tx_master_clk	:	in	std_logic	:=	'0';
		tx_master_clk_rst_n	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		pld_10g_krfec_tx_frame_krfec_reg	:	out	std_logic	:=	'0';
		pld_krfec_tx_alignment_plddirect_reg	:	out	std_logic	:=	'0';
		pld_krfec_tx_alignment_reg	:	out	std_logic	:=	'0';
		tx_alignment	:	out	std_logic	:=	'0';
		tx_data_out	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		tx_frame	:	out	std_logic	:=	'0';
		tx_test_data	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000"
	);
end twentynm_hssi_krfec_tx_pcs;

architecture behavior of twentynm_hssi_krfec_tx_pcs	is




component	twentynm_hssi_krfec_tx_pcs_encrypted
	generic (
		-- Architecture parameters
		burst_err	:	string	:=	"burst_err_dis";
		burst_err_len	:	string	:=	"burst_err_len1";
		ctrl_bit_reverse	:	string	:=	"ctrl_bit_reverse_dis";
		data_bit_reverse	:	string	:=	"data_bit_reverse_dis";
		enc_frame_query	:	string	:=	"enc_query_dis";
		low_latency_en	:	string	:=	"disable";
		pipeln_encoder	:	string	:=	"enable";
		pipeln_scrambler	:	string	:=	"enable";
		prot_mode	:	string	:=	"disable_mode";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode";
		transcode_err	:	string	:=	"trans_err_dis";
		transmit_order	:	string	:=	"transmit_lsb";
		tx_testbus_sel	:	string	:=	"overall"
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		tx_control_in	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		tx_data_in	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		tx_data_valid_in	:	in	std_logic	:=	'0';
		tx_krfec_clk	:	in	std_logic	:=	'0';
		tx_master_clk	:	in	std_logic	:=	'0';
		tx_master_clk_rst_n	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		pld_10g_krfec_tx_frame_krfec_reg	:	out	std_logic	:=	'0';
		pld_krfec_tx_alignment_plddirect_reg	:	out	std_logic	:=	'0';
		pld_krfec_tx_alignment_reg	:	out	std_logic	:=	'0';
		tx_alignment	:	out	std_logic	:=	'0';
		tx_data_out	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		tx_frame	:	out	std_logic	:=	'0';
		tx_test_data	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000"
	);
end component;

begin



inst : twentynm_hssi_krfec_tx_pcs_encrypted
	generic map (
		-- Instance parameters
		burst_err	=>	burst_err,
		burst_err_len	=>	burst_err_len,
		ctrl_bit_reverse	=>	ctrl_bit_reverse,
		data_bit_reverse	=>	data_bit_reverse,
		enc_frame_query	=>	enc_frame_query,
		low_latency_en	=>	low_latency_en,
		pipeln_encoder	=>	pipeln_encoder,
		pipeln_scrambler	=>	pipeln_scrambler,
		prot_mode	=>	prot_mode,
		silicon_rev	=>	silicon_rev,
		sup_mode	=>	sup_mode,
		transcode_err	=>	transcode_err,
		transmit_order	=>	transmit_order,
		tx_testbus_sel	=>	tx_testbus_sel
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		tx_control_in	=>	tx_control_in,
		tx_data_in	=>	tx_data_in,
		tx_data_valid_in	=>	tx_data_valid_in,
		tx_krfec_clk	=>	tx_krfec_clk,
		tx_master_clk	=>	tx_master_clk,
		tx_master_clk_rst_n	=>	tx_master_clk_rst_n,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		pld_10g_krfec_tx_frame_krfec_reg	=>	pld_10g_krfec_tx_frame_krfec_reg,
		pld_krfec_tx_alignment_plddirect_reg	=>	pld_krfec_tx_alignment_plddirect_reg,
		pld_krfec_tx_alignment_reg	=>	pld_krfec_tx_alignment_reg,
		tx_alignment	=>	tx_alignment,
		tx_data_out	=>	tx_data_out,
		tx_frame	=>	tx_frame,
		tx_test_data	=>	tx_test_data
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_pipe_gen1_2	is
	generic (
		-- Entity parameters
		elec_idle_delay_val	:	bit_vector	:=	B"000";
		error_replace_pad	:	string	:=	"replace_edb";
		hip_mode	:	string	:=	"dis_hip";
		ind_error_reporting	:	string	:=	"dis_ind_error_reporting";
		phystatus_delay_val	:	bit_vector	:=	B"000";
		phystatus_rst_toggle	:	string	:=	"dis_phystatus_rst_toggle";
		pipe_byte_de_serializer_en	:	string	:=	"dont_care_bds";
		prot_mode	:	string	:=	"pipe_g1";
		reconfig_settings	:	string	:=	"{}";
		rpre_emph_a_val	:	bit_vector	:=	B"000000";
		rpre_emph_b_val	:	bit_vector	:=	B"000000";
		rpre_emph_c_val	:	bit_vector	:=	B"000000";
		rpre_emph_d_val	:	bit_vector	:=	B"000000";
		rpre_emph_e_val	:	bit_vector	:=	B"000000";
		rvod_sel_a_val	:	bit_vector	:=	B"000000";
		rvod_sel_b_val	:	bit_vector	:=	B"000000";
		rvod_sel_c_val	:	bit_vector	:=	B"000000";
		rvod_sel_d_val	:	bit_vector	:=	B"000000";
		rvod_sel_e_val	:	bit_vector	:=	B"000000";
		rx_pipe_enable	:	string	:=	"dis_pipe_rx";
		rxdetect_bypass	:	string	:=	"dis_rxdetect_bypass";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode";
		tx_pipe_enable	:	string	:=	"dis_pipe_tx";
		txswing	:	string	:=	"dis_txswing"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		pcie_switch	:	in	std_logic	:=	'0';
		pipe_rx_clk	:	in	std_logic	:=	'0';
		pipe_tx_clk	:	in	std_logic	:=	'0';
		power_state_transition_done	:	in	std_logic	:=	'0';
		power_state_transition_done_ena	:	in	std_logic	:=	'0';
		powerdown	:	in	std_logic_vector(1 downto 0)	:=	"00";
		refclk_b	:	in	std_logic	:=	'0';
		refclk_b_reset	:	in	std_logic	:=	'0';
		rev_loopbk_pcs_gen3	:	in	std_logic	:=	'0';
		revloopback	:	in	std_logic	:=	'0';
		rx_detect_valid	:	in	std_logic	:=	'0';
		rx_found	:	in	std_logic	:=	'0';
		rx_pipe_reset	:	in	std_logic	:=	'0';
		rxd	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		rxelectricalidle	:	in	std_logic	:=	'0';
		rxelectricalidle_pcs_gen3	:	in	std_logic	:=	'0';
		rxpolarity	:	in	std_logic	:=	'0';
		rxpolarity_pcs_gen3	:	in	std_logic	:=	'0';
		sigdetni	:	in	std_logic	:=	'0';
		speed_change	:	in	std_logic	:=	'0';
		tx_elec_idle_comp	:	in	std_logic	:=	'0';
		tx_pipe_reset	:	in	std_logic	:=	'0';
		txd_ch	:	in	std_logic_vector(43 downto 0)	:=	"00000000000000000000000000000000000000000000";
		txdeemph	:	in	std_logic	:=	'0';
		txdetectrxloopback	:	in	std_logic	:=	'0';
		txelecidle	:	in	std_logic	:=	'0';
		txmargin	:	in	std_logic_vector(2 downto 0)	:=	"000";
		txswingport	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		pld_8g_rxpolarity_pipe3_reg	:	out	std_logic	:=	'0';
		current_coeff	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		phystatus	:	out	std_logic	:=	'0';
		polarity_inversion_rx	:	out	std_logic	:=	'0';
		rev_loopbk	:	out	std_logic	:=	'0';
		rxd_ch	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		rxelecidle	:	out	std_logic	:=	'0';
		rxelectricalidle_out	:	out	std_logic	:=	'0';
		rxstatus	:	out	std_logic_vector(2 downto 0)	:=	"000";
		rxvalid	:	out	std_logic	:=	'0';
		tx_elec_idle_out	:	out	std_logic	:=	'0';
		txd	:	out	std_logic_vector(43 downto 0)	:=	"00000000000000000000000000000000000000000000";
		txdetectrx	:	out	std_logic	:=	'0'
	);
end twentynm_hssi_pipe_gen1_2;

architecture behavior of twentynm_hssi_pipe_gen1_2	is

constant elec_idle_delay_val_int	:	integer	:=	bin2int(elec_idle_delay_val);
constant phystatus_delay_val_int	:	integer	:=	bin2int(phystatus_delay_val);
constant rpre_emph_a_val_int	:	integer	:=	bin2int(rpre_emph_a_val);
constant rpre_emph_b_val_int	:	integer	:=	bin2int(rpre_emph_b_val);
constant rpre_emph_c_val_int	:	integer	:=	bin2int(rpre_emph_c_val);
constant rpre_emph_d_val_int	:	integer	:=	bin2int(rpre_emph_d_val);
constant rpre_emph_e_val_int	:	integer	:=	bin2int(rpre_emph_e_val);
constant rvod_sel_a_val_int	:	integer	:=	bin2int(rvod_sel_a_val);
constant rvod_sel_b_val_int	:	integer	:=	bin2int(rvod_sel_b_val);
constant rvod_sel_c_val_int	:	integer	:=	bin2int(rvod_sel_c_val);
constant rvod_sel_d_val_int	:	integer	:=	bin2int(rvod_sel_d_val);
constant rvod_sel_e_val_int	:	integer	:=	bin2int(rvod_sel_e_val);



component	twentynm_hssi_pipe_gen1_2_encrypted
	generic (
		-- Architecture parameters
		elec_idle_delay_val	:	integer	:=	0;
		error_replace_pad	:	string	:=	"replace_edb";
		hip_mode	:	string	:=	"dis_hip";
		ind_error_reporting	:	string	:=	"dis_ind_error_reporting";
		phystatus_delay_val	:	integer	:=	0;
		phystatus_rst_toggle	:	string	:=	"dis_phystatus_rst_toggle";
		pipe_byte_de_serializer_en	:	string	:=	"dont_care_bds";
		prot_mode	:	string	:=	"pipe_g1";
		reconfig_settings	:	string	:=	"{}";
		rpre_emph_a_val	:	integer	:=	0;
		rpre_emph_b_val	:	integer	:=	0;
		rpre_emph_c_val	:	integer	:=	0;
		rpre_emph_d_val	:	integer	:=	0;
		rpre_emph_e_val	:	integer	:=	0;
		rvod_sel_a_val	:	integer	:=	0;
		rvod_sel_b_val	:	integer	:=	0;
		rvod_sel_c_val	:	integer	:=	0;
		rvod_sel_d_val	:	integer	:=	0;
		rvod_sel_e_val	:	integer	:=	0;
		rx_pipe_enable	:	string	:=	"dis_pipe_rx";
		rxdetect_bypass	:	string	:=	"dis_rxdetect_bypass";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode";
		tx_pipe_enable	:	string	:=	"dis_pipe_tx";
		txswing	:	string	:=	"dis_txswing"
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		pcie_switch	:	in	std_logic	:=	'0';
		pipe_rx_clk	:	in	std_logic	:=	'0';
		pipe_tx_clk	:	in	std_logic	:=	'0';
		power_state_transition_done	:	in	std_logic	:=	'0';
		power_state_transition_done_ena	:	in	std_logic	:=	'0';
		powerdown	:	in	std_logic_vector(1 downto 0)	:=	"00";
		refclk_b	:	in	std_logic	:=	'0';
		refclk_b_reset	:	in	std_logic	:=	'0';
		rev_loopbk_pcs_gen3	:	in	std_logic	:=	'0';
		revloopback	:	in	std_logic	:=	'0';
		rx_detect_valid	:	in	std_logic	:=	'0';
		rx_found	:	in	std_logic	:=	'0';
		rx_pipe_reset	:	in	std_logic	:=	'0';
		rxd	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		rxelectricalidle	:	in	std_logic	:=	'0';
		rxelectricalidle_pcs_gen3	:	in	std_logic	:=	'0';
		rxpolarity	:	in	std_logic	:=	'0';
		rxpolarity_pcs_gen3	:	in	std_logic	:=	'0';
		sigdetni	:	in	std_logic	:=	'0';
		speed_change	:	in	std_logic	:=	'0';
		tx_elec_idle_comp	:	in	std_logic	:=	'0';
		tx_pipe_reset	:	in	std_logic	:=	'0';
		txd_ch	:	in	std_logic_vector(43 downto 0)	:=	"00000000000000000000000000000000000000000000";
		txdeemph	:	in	std_logic	:=	'0';
		txdetectrxloopback	:	in	std_logic	:=	'0';
		txelecidle	:	in	std_logic	:=	'0';
		txmargin	:	in	std_logic_vector(2 downto 0)	:=	"000";
		txswingport	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		pld_8g_rxpolarity_pipe3_reg	:	out	std_logic	:=	'0';
		current_coeff	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		phystatus	:	out	std_logic	:=	'0';
		polarity_inversion_rx	:	out	std_logic	:=	'0';
		rev_loopbk	:	out	std_logic	:=	'0';
		rxd_ch	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		rxelecidle	:	out	std_logic	:=	'0';
		rxelectricalidle_out	:	out	std_logic	:=	'0';
		rxstatus	:	out	std_logic_vector(2 downto 0)	:=	"000";
		rxvalid	:	out	std_logic	:=	'0';
		tx_elec_idle_out	:	out	std_logic	:=	'0';
		txd	:	out	std_logic_vector(43 downto 0)	:=	"00000000000000000000000000000000000000000000";
		txdetectrx	:	out	std_logic	:=	'0'
	);
end component;

begin



inst : twentynm_hssi_pipe_gen1_2_encrypted
	generic map (
		-- Instance parameters
		elec_idle_delay_val	=>	elec_idle_delay_val_int,
		error_replace_pad	=>	error_replace_pad,
		hip_mode	=>	hip_mode,
		ind_error_reporting	=>	ind_error_reporting,
		phystatus_delay_val	=>	phystatus_delay_val_int,
		phystatus_rst_toggle	=>	phystatus_rst_toggle,
		pipe_byte_de_serializer_en	=>	pipe_byte_de_serializer_en,
		prot_mode	=>	prot_mode,
		reconfig_settings	=>	reconfig_settings,
		rpre_emph_a_val	=>	rpre_emph_a_val_int,
		rpre_emph_b_val	=>	rpre_emph_b_val_int,
		rpre_emph_c_val	=>	rpre_emph_c_val_int,
		rpre_emph_d_val	=>	rpre_emph_d_val_int,
		rpre_emph_e_val	=>	rpre_emph_e_val_int,
		rvod_sel_a_val	=>	rvod_sel_a_val_int,
		rvod_sel_b_val	=>	rvod_sel_b_val_int,
		rvod_sel_c_val	=>	rvod_sel_c_val_int,
		rvod_sel_d_val	=>	rvod_sel_d_val_int,
		rvod_sel_e_val	=>	rvod_sel_e_val_int,
		rx_pipe_enable	=>	rx_pipe_enable,
		rxdetect_bypass	=>	rxdetect_bypass,
		silicon_rev	=>	silicon_rev,
		sup_mode	=>	sup_mode,
		tx_pipe_enable	=>	tx_pipe_enable,
		txswing	=>	txswing
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		pcie_switch	=>	pcie_switch,
		pipe_rx_clk	=>	pipe_rx_clk,
		pipe_tx_clk	=>	pipe_tx_clk,
		power_state_transition_done	=>	power_state_transition_done,
		power_state_transition_done_ena	=>	power_state_transition_done_ena,
		powerdown	=>	powerdown,
		refclk_b	=>	refclk_b,
		refclk_b_reset	=>	refclk_b_reset,
		rev_loopbk_pcs_gen3	=>	rev_loopbk_pcs_gen3,
		revloopback	=>	revloopback,
		rx_detect_valid	=>	rx_detect_valid,
		rx_found	=>	rx_found,
		rx_pipe_reset	=>	rx_pipe_reset,
		rxd	=>	rxd,
		rxelectricalidle	=>	rxelectricalidle,
		rxelectricalidle_pcs_gen3	=>	rxelectricalidle_pcs_gen3,
		rxpolarity	=>	rxpolarity,
		rxpolarity_pcs_gen3	=>	rxpolarity_pcs_gen3,
		sigdetni	=>	sigdetni,
		speed_change	=>	speed_change,
		tx_elec_idle_comp	=>	tx_elec_idle_comp,
		tx_pipe_reset	=>	tx_pipe_reset,
		txd_ch	=>	txd_ch,
		txdeemph	=>	txdeemph,
		txdetectrxloopback	=>	txdetectrxloopback,
		txelecidle	=>	txelecidle,
		txmargin	=>	txmargin,
		txswingport	=>	txswingport,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		pld_8g_rxpolarity_pipe3_reg	=>	pld_8g_rxpolarity_pipe3_reg,
		current_coeff	=>	current_coeff,
		phystatus	=>	phystatus,
		polarity_inversion_rx	=>	polarity_inversion_rx,
		rev_loopbk	=>	rev_loopbk,
		rxd_ch	=>	rxd_ch,
		rxelecidle	=>	rxelecidle,
		rxelectricalidle_out	=>	rxelectricalidle_out,
		rxstatus	=>	rxstatus,
		rxvalid	=>	rxvalid,
		tx_elec_idle_out	=>	tx_elec_idle_out,
		txd	=>	txd,
		txdetectrx	=>	txdetectrx
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_pipe_gen3	is
	generic (
		-- Entity parameters
		bypass_rx_detection_enable	:	string	:=	"false";
		bypass_rx_preset	:	bit_vector	:=	B"000";
		bypass_rx_preset_enable	:	string	:=	"false";
		bypass_tx_coefficent	:	bit_vector	:=	B"000000000000000000";
		bypass_tx_coefficent_enable	:	string	:=	"false";
		elecidle_delay_g3	:	bit_vector	:=	B"110";
		ind_error_reporting	:	string	:=	"dis_ind_error_reporting";
		mode	:	string	:=	"pipe_g1";
		phy_status_delay_g12	:	bit_vector	:=	B"101";
		phy_status_delay_g3	:	bit_vector	:=	B"101";
		phystatus_rst_toggle_g12	:	string	:=	"dis_phystatus_rst_toggle";
		phystatus_rst_toggle_g3	:	string	:=	"dis_phystatus_rst_toggle_g3";
		rate_match_pad_insertion	:	string	:=	"dis_rm_fifo_pad_ins";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode";
		test_out_sel	:	string	:=	"disable_test_out"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		blk_algnd_int	:	in	std_logic	:=	'0';
		clkcomp_delete_int	:	in	std_logic	:=	'0';
		clkcomp_insert_int	:	in	std_logic	:=	'0';
		clkcomp_overfl_int	:	in	std_logic	:=	'0';
		clkcomp_undfl_int	:	in	std_logic	:=	'0';
		current_coeff	:	in	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_rxpreset	:	in	std_logic_vector(2 downto 0)	:=	"000";
		err_decode_int	:	in	std_logic	:=	'0';
		pcs_asn_bundling_in	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		pipe_tx_clk	:	in	std_logic	:=	'0';
		pipe_tx_rstn	:	in	std_logic	:=	'0';
		pma_rx_detect_valid	:	in	std_logic	:=	'0';
		pma_rx_found	:	in	std_logic	:=	'0';
		pma_signal_det	:	in	std_logic	:=	'0';
		powerdown	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rcv_lfsr_chk_int	:	in	std_logic	:=	'0';
		rx_blk_start_int	:	in	std_logic	:=	'0';
		rx_sync_hdr_int	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rx_test_out	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		rxd_8gpcs_in	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		rxdata_int	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdatak_int	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdataskip_int	:	in	std_logic	:=	'0';
		rxelecidle_8gpcs_in	:	in	std_logic	:=	'0';
		rxpolarity	:	in	std_logic	:=	'0';
		tx_blk_start	:	in	std_logic	:=	'0';
		tx_sync_hdr	:	in	std_logic_vector(1 downto 0)	:=	"00";
		tx_test_out	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		txcompliance	:	in	std_logic	:=	'0';
		txdata	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdatak	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		txdataskip	:	in	std_logic	:=	'0';
		txdeemph	:	in	std_logic	:=	'0';
		txdetectrxloopback	:	in	std_logic	:=	'0';
		txelecidle	:	in	std_logic	:=	'0';
		txmargin	:	in	std_logic_vector(2 downto 0)	:=	"000";
		txswing	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		dis_pc_byte	:	out	std_logic	:=	'0';
		gen3_clk_sel	:	out	std_logic	:=	'0';
		pcs_rst	:	out	std_logic	:=	'0';
		phystatus	:	out	std_logic	:=	'0';
		pma_current_coeff	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		pma_current_rxpreset	:	out	std_logic_vector(2 downto 0)	:=	"000";
		pma_rx_det_pd	:	out	std_logic	:=	'0';
		pma_tx_elec_idle	:	out	std_logic	:=	'0';
		pma_txdeemph	:	out	std_logic	:=	'0';
		pma_txdetectrx	:	out	std_logic	:=	'0';
		pma_txmargin	:	out	std_logic_vector(2 downto 0)	:=	"000";
		pma_txswing	:	out	std_logic	:=	'0';
		reset_pc_prts	:	out	std_logic	:=	'0';
		rev_lpbk_8gpcs_out	:	out	std_logic	:=	'0';
		rev_lpbk_int	:	out	std_logic	:=	'0';
		rx_blk_start	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		rx_sync_hdr	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rxd_8gpcs_out	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		rxdataskip	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		rxelecidle	:	out	std_logic	:=	'0';
		rxpolarity_8gpcs_out	:	out	std_logic	:=	'0';
		rxpolarity_int	:	out	std_logic	:=	'0';
		rxstatus	:	out	std_logic_vector(2 downto 0)	:=	"000";
		rxvalid	:	out	std_logic	:=	'0';
		shutdown_clk	:	out	std_logic	:=	'0';
		test_out	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		tx_blk_start_int	:	out	std_logic	:=	'0';
		tx_sync_hdr_int	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txdata_int	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdatak_int	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdataskip_int	:	out	std_logic	:=	'0'
	);
end twentynm_hssi_pipe_gen3;

architecture behavior of twentynm_hssi_pipe_gen3	is

constant bypass_rx_preset_int	:	integer	:=	bin2int(bypass_rx_preset);
constant bypass_tx_coefficent_int	:	integer	:=	bin2int(bypass_tx_coefficent);
constant elecidle_delay_g3_int	:	integer	:=	bin2int(elecidle_delay_g3);
constant phy_status_delay_g12_int	:	integer	:=	bin2int(phy_status_delay_g12);
constant phy_status_delay_g3_int	:	integer	:=	bin2int(phy_status_delay_g3);



component	twentynm_hssi_pipe_gen3_encrypted
	generic (
		-- Architecture parameters
		bypass_rx_detection_enable	:	string	:=	"false";
		bypass_rx_preset	:	integer	:=	0;
		bypass_rx_preset_enable	:	string	:=	"false";
		bypass_tx_coefficent	:	integer	:=	0;
		bypass_tx_coefficent_enable	:	string	:=	"false";
		elecidle_delay_g3	:	integer	:=	6;
		ind_error_reporting	:	string	:=	"dis_ind_error_reporting";
		mode	:	string	:=	"pipe_g1";
		phy_status_delay_g12	:	integer	:=	5;
		phy_status_delay_g3	:	integer	:=	5;
		phystatus_rst_toggle_g12	:	string	:=	"dis_phystatus_rst_toggle";
		phystatus_rst_toggle_g3	:	string	:=	"dis_phystatus_rst_toggle_g3";
		rate_match_pad_insertion	:	string	:=	"dis_rm_fifo_pad_ins";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode";
		test_out_sel	:	string	:=	"disable_test_out"
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		blk_algnd_int	:	in	std_logic	:=	'0';
		clkcomp_delete_int	:	in	std_logic	:=	'0';
		clkcomp_insert_int	:	in	std_logic	:=	'0';
		clkcomp_overfl_int	:	in	std_logic	:=	'0';
		clkcomp_undfl_int	:	in	std_logic	:=	'0';
		current_coeff	:	in	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_rxpreset	:	in	std_logic_vector(2 downto 0)	:=	"000";
		err_decode_int	:	in	std_logic	:=	'0';
		pcs_asn_bundling_in	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		pipe_tx_clk	:	in	std_logic	:=	'0';
		pipe_tx_rstn	:	in	std_logic	:=	'0';
		pma_rx_detect_valid	:	in	std_logic	:=	'0';
		pma_rx_found	:	in	std_logic	:=	'0';
		pma_signal_det	:	in	std_logic	:=	'0';
		powerdown	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rcv_lfsr_chk_int	:	in	std_logic	:=	'0';
		rx_blk_start_int	:	in	std_logic	:=	'0';
		rx_sync_hdr_int	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rx_test_out	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		rxd_8gpcs_in	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		rxdata_int	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdatak_int	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdataskip_int	:	in	std_logic	:=	'0';
		rxelecidle_8gpcs_in	:	in	std_logic	:=	'0';
		rxpolarity	:	in	std_logic	:=	'0';
		tx_blk_start	:	in	std_logic	:=	'0';
		tx_sync_hdr	:	in	std_logic_vector(1 downto 0)	:=	"00";
		tx_test_out	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		txcompliance	:	in	std_logic	:=	'0';
		txdata	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdatak	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		txdataskip	:	in	std_logic	:=	'0';
		txdeemph	:	in	std_logic	:=	'0';
		txdetectrxloopback	:	in	std_logic	:=	'0';
		txelecidle	:	in	std_logic	:=	'0';
		txmargin	:	in	std_logic_vector(2 downto 0)	:=	"000";
		txswing	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		dis_pc_byte	:	out	std_logic	:=	'0';
		gen3_clk_sel	:	out	std_logic	:=	'0';
		pcs_rst	:	out	std_logic	:=	'0';
		phystatus	:	out	std_logic	:=	'0';
		pma_current_coeff	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		pma_current_rxpreset	:	out	std_logic_vector(2 downto 0)	:=	"000";
		pma_rx_det_pd	:	out	std_logic	:=	'0';
		pma_tx_elec_idle	:	out	std_logic	:=	'0';
		pma_txdeemph	:	out	std_logic	:=	'0';
		pma_txdetectrx	:	out	std_logic	:=	'0';
		pma_txmargin	:	out	std_logic_vector(2 downto 0)	:=	"000";
		pma_txswing	:	out	std_logic	:=	'0';
		reset_pc_prts	:	out	std_logic	:=	'0';
		rev_lpbk_8gpcs_out	:	out	std_logic	:=	'0';
		rev_lpbk_int	:	out	std_logic	:=	'0';
		rx_blk_start	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		rx_sync_hdr	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rxd_8gpcs_out	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		rxdataskip	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		rxelecidle	:	out	std_logic	:=	'0';
		rxpolarity_8gpcs_out	:	out	std_logic	:=	'0';
		rxpolarity_int	:	out	std_logic	:=	'0';
		rxstatus	:	out	std_logic_vector(2 downto 0)	:=	"000";
		rxvalid	:	out	std_logic	:=	'0';
		shutdown_clk	:	out	std_logic	:=	'0';
		test_out	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		tx_blk_start_int	:	out	std_logic	:=	'0';
		tx_sync_hdr_int	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txdata_int	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdatak_int	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdataskip_int	:	out	std_logic	:=	'0'
	);
end component;

begin



inst : twentynm_hssi_pipe_gen3_encrypted
	generic map (
		-- Instance parameters
		bypass_rx_detection_enable	=>	bypass_rx_detection_enable,
		bypass_rx_preset	=>	bypass_rx_preset_int,
		bypass_rx_preset_enable	=>	bypass_rx_preset_enable,
		bypass_tx_coefficent	=>	bypass_tx_coefficent_int,
		bypass_tx_coefficent_enable	=>	bypass_tx_coefficent_enable,
		elecidle_delay_g3	=>	elecidle_delay_g3_int,
		ind_error_reporting	=>	ind_error_reporting,
		mode	=>	mode,
		phy_status_delay_g12	=>	phy_status_delay_g12_int,
		phy_status_delay_g3	=>	phy_status_delay_g3_int,
		phystatus_rst_toggle_g12	=>	phystatus_rst_toggle_g12,
		phystatus_rst_toggle_g3	=>	phystatus_rst_toggle_g3,
		rate_match_pad_insertion	=>	rate_match_pad_insertion,
		silicon_rev	=>	silicon_rev,
		sup_mode	=>	sup_mode,
		test_out_sel	=>	test_out_sel
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		blk_algnd_int	=>	blk_algnd_int,
		clkcomp_delete_int	=>	clkcomp_delete_int,
		clkcomp_insert_int	=>	clkcomp_insert_int,
		clkcomp_overfl_int	=>	clkcomp_overfl_int,
		clkcomp_undfl_int	=>	clkcomp_undfl_int,
		current_coeff	=>	current_coeff,
		current_rxpreset	=>	current_rxpreset,
		err_decode_int	=>	err_decode_int,
		pcs_asn_bundling_in	=>	pcs_asn_bundling_in,
		pipe_tx_clk	=>	pipe_tx_clk,
		pipe_tx_rstn	=>	pipe_tx_rstn,
		pma_rx_detect_valid	=>	pma_rx_detect_valid,
		pma_rx_found	=>	pma_rx_found,
		pma_signal_det	=>	pma_signal_det,
		powerdown	=>	powerdown,
		rcv_lfsr_chk_int	=>	rcv_lfsr_chk_int,
		rx_blk_start_int	=>	rx_blk_start_int,
		rx_sync_hdr_int	=>	rx_sync_hdr_int,
		rx_test_out	=>	rx_test_out,
		rxd_8gpcs_in	=>	rxd_8gpcs_in,
		rxdata_int	=>	rxdata_int,
		rxdatak_int	=>	rxdatak_int,
		rxdataskip_int	=>	rxdataskip_int,
		rxelecidle_8gpcs_in	=>	rxelecidle_8gpcs_in,
		rxpolarity	=>	rxpolarity,
		tx_blk_start	=>	tx_blk_start,
		tx_sync_hdr	=>	tx_sync_hdr,
		tx_test_out	=>	tx_test_out,
		txcompliance	=>	txcompliance,
		txdata	=>	txdata,
		txdatak	=>	txdatak,
		txdataskip	=>	txdataskip,
		txdeemph	=>	txdeemph,
		txdetectrxloopback	=>	txdetectrxloopback,
		txelecidle	=>	txelecidle,
		txmargin	=>	txmargin,
		txswing	=>	txswing,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		dis_pc_byte	=>	dis_pc_byte,
		gen3_clk_sel	=>	gen3_clk_sel,
		pcs_rst	=>	pcs_rst,
		phystatus	=>	phystatus,
		pma_current_coeff	=>	pma_current_coeff,
		pma_current_rxpreset	=>	pma_current_rxpreset,
		pma_rx_det_pd	=>	pma_rx_det_pd,
		pma_tx_elec_idle	=>	pma_tx_elec_idle,
		pma_txdeemph	=>	pma_txdeemph,
		pma_txdetectrx	=>	pma_txdetectrx,
		pma_txmargin	=>	pma_txmargin,
		pma_txswing	=>	pma_txswing,
		reset_pc_prts	=>	reset_pc_prts,
		rev_lpbk_8gpcs_out	=>	rev_lpbk_8gpcs_out,
		rev_lpbk_int	=>	rev_lpbk_int,
		rx_blk_start	=>	rx_blk_start,
		rx_sync_hdr	=>	rx_sync_hdr,
		rxd_8gpcs_out	=>	rxd_8gpcs_out,
		rxdataskip	=>	rxdataskip,
		rxelecidle	=>	rxelecidle,
		rxpolarity_8gpcs_out	=>	rxpolarity_8gpcs_out,
		rxpolarity_int	=>	rxpolarity_int,
		rxstatus	=>	rxstatus,
		rxvalid	=>	rxvalid,
		shutdown_clk	=>	shutdown_clk,
		test_out	=>	test_out,
		tx_blk_start_int	=>	tx_blk_start_int,
		tx_sync_hdr_int	=>	tx_sync_hdr_int,
		txdata_int	=>	txdata_int,
		txdatak_int	=>	txdatak_int,
		txdataskip_int	=>	txdataskip_int
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_pma_adaptation	is
	generic (
		-- Entity parameters
		adapt_dfe_control_sel	:	string	:=	"r_adapt_dfe_control_sel_0";
		adapt_dfe_sel	:	string	:=	"r_adapt_dfe_sel_0";
		adapt_mode	:	string	:=	"dfe_vga";
		adapt_vga_sel	:	string	:=	"r_adapt_vga_sel_0";
		adapt_vref_sel	:	string	:=	"r_adapt_vref_sel_0";
		adp_1s_ctle_bypass	:	string	:=	"radp_1s_ctle_bypass_0";
		adp_4s_ctle_bypass	:	string	:=	"radp_4s_ctle_bypass_0";
		adp_adapt_control_sel	:	string	:=	"radp_adapt_control_sel_0";
		adp_adapt_rstn	:	string	:=	"radp_adapt_rstn_1";
		adp_adapt_start	:	string	:=	"radp_adapt_start_0";
		adp_bist_auxpath_en	:	string	:=	"radp_bist_auxpath_disable";
		adp_bist_count_rstn	:	string	:=	"radp_bist_count_rstn_0";
		adp_bist_datapath_en	:	string	:=	"radp_bist_datapath_disable";
		adp_bist_mode	:	string	:=	"radp_bist_mode_0";
		adp_bist_odi_dfe_sel	:	string	:=	"radp_bist_odi_dfe_sel_0";
		adp_bist_spec_en	:	string	:=	"radp_bist_spec_en_0";
		adp_control_mux_bypass	:	string	:=	"radp_control_mux_bypass_0";
		adp_ctle_acgain_4s	:	string	:=	"radp_ctle_acgain_4s_0";
		adp_ctle_adapt_bw	:	string	:=	"radp_ctle_adapt_bw_3";
		adp_ctle_adapt_cycle_window	:	string	:=	"radp_ctle_adapt_cycle_window_6";
		adp_ctle_adapt_oneshot	:	string	:=	"radp_ctle_adapt_oneshot_1";
		adp_ctle_en	:	string	:=	"radp_ctle_disable";
		adp_ctle_eqz_1s_sel	:	string	:=	"radp_ctle_eqz_1s_sel_0";
		adp_ctle_force_spec_sign	:	string	:=	"radp_ctle_force_spec_sign_0";
		adp_ctle_hold_en	:	string	:=	"radp_ctle_not_held";
		adp_ctle_load	:	string	:=	"radp_ctle_load_0";
		adp_ctle_load_value	:	string	:=	"radp_ctle_load_value_0";
		adp_ctle_scale	:	string	:=	"radp_ctle_scale_0";
		adp_ctle_scale_en	:	string	:=	"radp_ctle_scale_en_0";
		adp_ctle_spec_sign	:	string	:=	"radp_ctle_spec_sign_0";
		adp_ctle_sweep_direction	:	string	:=	"radp_ctle_sweep_direction_1";
		adp_ctle_threshold	:	string	:=	"radp_ctle_threshold_0";
		adp_ctle_threshold_en	:	string	:=	"radp_ctle_threshold_en_0";
		adp_ctle_vref_polarity	:	string	:=	"radp_ctle_vref_polarity_0";
		adp_ctle_window	:	string	:=	"radp_ctle_window_0";
		adp_dfe_bw	:	string	:=	"radp_dfe_bw_3";
		adp_dfe_clkout_div_sel	:	string	:=	"radp_dfe_clkout_div_sel_0";
		adp_dfe_cycle	:	string	:=	"radp_dfe_cycle_6";
		adp_dfe_fltap_bypass	:	string	:=	"radp_dfe_fltap_bypass_0";
		adp_dfe_fltap_en	:	string	:=	"radp_dfe_fltap_disable";
		adp_dfe_fltap_hold_en	:	string	:=	"radp_dfe_fltap_not_held";
		adp_dfe_fltap_load	:	string	:=	"radp_dfe_fltap_load_0";
		adp_dfe_fltap_position	:	string	:=	"radp_dfe_fltap_position_0";
		adp_dfe_force_spec_sign	:	string	:=	"radp_dfe_force_spec_sign_0";
		adp_dfe_fxtap1	:	string	:=	"radp_dfe_fxtap1_0";
		adp_dfe_fxtap10	:	string	:=	"radp_dfe_fxtap10_0";
		adp_dfe_fxtap10_sgn	:	string	:=	"radp_dfe_fxtap10_sgn_0";
		adp_dfe_fxtap11	:	string	:=	"radp_dfe_fxtap11_0";
		adp_dfe_fxtap11_sgn	:	string	:=	"radp_dfe_fxtap11_sgn_0";
		adp_dfe_fxtap2	:	string	:=	"radp_dfe_fxtap2_0";
		adp_dfe_fxtap2_sgn	:	string	:=	"radp_dfe_fxtap2_sgn_0";
		adp_dfe_fxtap3	:	string	:=	"radp_dfe_fxtap3_0";
		adp_dfe_fxtap3_sgn	:	string	:=	"radp_dfe_fxtap3_sgn_0";
		adp_dfe_fxtap4	:	string	:=	"radp_dfe_fxtap4_0";
		adp_dfe_fxtap4_sgn	:	string	:=	"radp_dfe_fxtap4_sgn_0";
		adp_dfe_fxtap5	:	string	:=	"radp_dfe_fxtap5_0";
		adp_dfe_fxtap5_sgn	:	string	:=	"radp_dfe_fxtap5_sgn_0";
		adp_dfe_fxtap6	:	string	:=	"radp_dfe_fxtap6_0";
		adp_dfe_fxtap6_sgn	:	string	:=	"radp_dfe_fxtap6_sgn_0";
		adp_dfe_fxtap7	:	string	:=	"radp_dfe_fxtap7_0";
		adp_dfe_fxtap7_sgn	:	string	:=	"radp_dfe_fxtap7_sgn_0";
		adp_dfe_fxtap8	:	string	:=	"radp_dfe_fxtap8_0";
		adp_dfe_fxtap8_sgn	:	string	:=	"radp_dfe_fxtap8_sgn_0";
		adp_dfe_fxtap9	:	string	:=	"radp_dfe_fxtap9_0";
		adp_dfe_fxtap9_sgn	:	string	:=	"radp_dfe_fxtap9_sgn_0";
		adp_dfe_fxtap_bypass	:	string	:=	"radp_dfe_fxtap_bypass_0";
		adp_dfe_fxtap_en	:	string	:=	"radp_dfe_fxtap_disable";
		adp_dfe_fxtap_hold_en	:	string	:=	"radp_dfe_fxtap_not_held";
		adp_dfe_fxtap_load	:	string	:=	"radp_dfe_fxtap_load_0";
		adp_dfe_mode	:	string	:=	"radp_dfe_mode_0";
		adp_dfe_spec_sign	:	string	:=	"radp_dfe_spec_sign_0";
		adp_dfe_vref_polarity	:	string	:=	"radp_dfe_vref_polarity_0";
		adp_force_freqlock	:	string	:=	"radp_force_freqlock_off";
		adp_frame_capture	:	string	:=	"radp_frame_capture_0";
		adp_frame_en	:	string	:=	"radp_frame_en_0";
		adp_frame_odi_sel	:	string	:=	"radp_frame_odi_sel_0";
		adp_frame_out_sel	:	string	:=	"radp_frame_out_sel_0";
		adp_lfeq_fb_sel	:	string	:=	"radp_lfeq_fb_sel_0";
		adp_mode	:	string	:=	"radp_mode_0";
		adp_odi_control_sel	:	string	:=	"radp_odi_control_sel_0";
		adp_onetime_dfe	:	string	:=	"radp_onetime_dfe_0";
		adp_spec_avg_window	:	string	:=	"radp_spec_avg_window_4";
		adp_spec_trans_filter	:	string	:=	"radp_spec_trans_filter_2";
		adp_status_sel	:	string	:=	"radp_status_sel_0";
		adp_vga_bypass	:	string	:=	"radp_vga_bypass_0";
		adp_vga_en	:	string	:=	"radp_vga_disable";
		adp_vga_load	:	string	:=	"radp_vga_load_0";
		adp_vga_polarity	:	string	:=	"radp_vga_polarity_0";
		adp_vga_sel	:	string	:=	"radp_vga_sel_0";
		adp_vga_sweep_direction	:	string	:=	"radp_vga_sweep_direction_1";
		adp_vga_threshold	:	string	:=	"radp_vga_threshold_4";
		adp_vref_bw	:	string	:=	"radp_vref_bw_1";
		adp_vref_bypass	:	string	:=	"radp_vref_bypass_0";
		adp_vref_cycle	:	string	:=	"radp_vref_cycle_6";
		adp_vref_dfe_spec_en	:	string	:=	"radp_vref_dfe_spec_en_0";
		adp_vref_en	:	string	:=	"radp_vref_disable";
		adp_vref_hold_en	:	string	:=	"radp_vref_not_held";
		adp_vref_load	:	string	:=	"radp_vref_load_0";
		adp_vref_polarity	:	string	:=	"radp_vref_polarity_0";
		adp_vref_sel	:	string	:=	"radp_vref_sel_21";
		adp_vref_vga_level	:	string	:=	"radp_vref_vga_level_13";
		datarate	:	string	:=	"0 bps";
		initial_settings	:	string	:=	"true";
		odi_count_threshold	:	string	:=	"rodi_count_threshold_0";
		odi_dfe_spec_en	:	string	:=	"rodi_dfe_spec_en_0";
		odi_en	:	string	:=	"rodi_en_0";
		odi_mode	:	string	:=	"rodi_mode_0";
		odi_rstn	:	string	:=	"rodi_rstn_0";
		odi_spec_sel	:	string	:=	"rodi_spec_sel_0";
		odi_start	:	string	:=	"rodi_start_0";
		odi_vref_sel	:	string	:=	"rodi_vref_sel_0";
		optimal	:	string	:=	"false";
		prot_mode	:	string	:=	"basic_rx";
		rrx_pcie_eqz	:	string	:=	"rrx_pcie_eqz_0";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		adapt_reset	:	in	std_logic	:=	'0';
		adapt_start	:	in	std_logic	:=	'0';
		deser_clk	:	in	std_logic	:=	'0';
		deser_data	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		deser_error	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		deser_odi	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		deser_odi_clk	:	in	std_logic	:=	'0';
		global_pipe_se	:	in	std_logic	:=	'0';
		i_rxpreset	:	in	std_logic_vector(2 downto 0)	:=	"000";
		radp_ctle_hold_en	:	in	std_logic	:=	'0';
		radp_ctle_patt_en	:	in	std_logic	:=	'0';
		radp_ctle_preset_sel	:	in	std_logic	:=	'0';
		radp_enable_max_lfeq_scale	:	in	std_logic	:=	'0';
		radp_lfeq_hold_en	:	in	std_logic	:=	'0';
		radp_vga_polarity	:	in	std_logic	:=	'0';
		rx_pllfreqlock	:	in	std_logic	:=	'0';
		scan_clk	:	in	std_logic	:=	'0';
		scan_in	:	in	std_logic_vector(9 downto 0)	:=	"0000000000";
		test_mode	:	in	std_logic	:=	'0';
		test_se	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		ctle_acgain_4s	:	out	std_logic_vector(27 downto 0)	:=	"0000000000000000000000000000";
		ctle_eqz_1s_sel	:	out	std_logic_vector(14 downto 0)	:=	"000000000000000";
		ctle_lfeq_fb_sel	:	out	std_logic_vector(6 downto 0)	:=	"0000000";
		dfe_adapt_en	:	out	std_logic	:=	'0';
		dfe_adp_clk	:	out	std_logic	:=	'0';
		dfe_fltap1	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		dfe_fltap1_sgn	:	out	std_logic	:=	'0';
		dfe_fltap2	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		dfe_fltap2_sgn	:	out	std_logic	:=	'0';
		dfe_fltap3	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		dfe_fltap3_sgn	:	out	std_logic	:=	'0';
		dfe_fltap4	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		dfe_fltap4_sgn	:	out	std_logic	:=	'0';
		dfe_fltap_bypdeser	:	out	std_logic	:=	'0';
		dfe_fltap_position	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		dfe_fxtap1	:	out	std_logic_vector(6 downto 0)	:=	"0000000";
		dfe_fxtap2	:	out	std_logic_vector(6 downto 0)	:=	"0000000";
		dfe_fxtap2_sgn	:	out	std_logic	:=	'0';
		dfe_fxtap3	:	out	std_logic_vector(6 downto 0)	:=	"0000000";
		dfe_fxtap3_sgn	:	out	std_logic	:=	'0';
		dfe_fxtap4	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		dfe_fxtap4_sgn	:	out	std_logic	:=	'0';
		dfe_fxtap5	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		dfe_fxtap5_sgn	:	out	std_logic	:=	'0';
		dfe_fxtap6	:	out	std_logic_vector(4 downto 0)	:=	"00000";
		dfe_fxtap6_sgn	:	out	std_logic	:=	'0';
		dfe_fxtap7	:	out	std_logic_vector(4 downto 0)	:=	"00000";
		dfe_fxtap7_sgn	:	out	std_logic	:=	'0';
		dfe_spec_disable	:	out	std_logic	:=	'0';
		dfe_spec_sign_sel	:	out	std_logic	:=	'0';
		dfe_vref_sign_sel	:	out	std_logic	:=	'0';
		odi_vref	:	out	std_logic_vector(4 downto 0)	:=	"00000";
		scan_out	:	out	std_logic_vector(9 downto 0)	:=	"0000000000";
		status_bus	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		vga_sel	:	out	std_logic_vector(6 downto 0)	:=	"0000000";
		vref_sel	:	out	std_logic_vector(4 downto 0)	:=	"00000"
	);
end twentynm_hssi_pma_adaptation;

architecture behavior of twentynm_hssi_pma_adaptation	is




component	twentynm_hssi_pma_adaptation_encrypted
	generic (
		-- Architecture parameters
		adapt_dfe_control_sel	:	string	:=	"r_adapt_dfe_control_sel_0";
		adapt_dfe_sel	:	string	:=	"r_adapt_dfe_sel_0";
		adapt_mode	:	string	:=	"dfe_vga";
		adapt_vga_sel	:	string	:=	"r_adapt_vga_sel_0";
		adapt_vref_sel	:	string	:=	"r_adapt_vref_sel_0";
		adp_1s_ctle_bypass	:	string	:=	"radp_1s_ctle_bypass_0";
		adp_4s_ctle_bypass	:	string	:=	"radp_4s_ctle_bypass_0";
		adp_adapt_control_sel	:	string	:=	"radp_adapt_control_sel_0";
		adp_adapt_rstn	:	string	:=	"radp_adapt_rstn_1";
		adp_adapt_start	:	string	:=	"radp_adapt_start_0";
		adp_bist_auxpath_en	:	string	:=	"radp_bist_auxpath_disable";
		adp_bist_count_rstn	:	string	:=	"radp_bist_count_rstn_0";
		adp_bist_datapath_en	:	string	:=	"radp_bist_datapath_disable";
		adp_bist_mode	:	string	:=	"radp_bist_mode_0";
		adp_bist_odi_dfe_sel	:	string	:=	"radp_bist_odi_dfe_sel_0";
		adp_bist_spec_en	:	string	:=	"radp_bist_spec_en_0";
		adp_control_mux_bypass	:	string	:=	"radp_control_mux_bypass_0";
		adp_ctle_acgain_4s	:	string	:=	"radp_ctle_acgain_4s_0";
		adp_ctle_adapt_bw	:	string	:=	"radp_ctle_adapt_bw_3";
		adp_ctle_adapt_cycle_window	:	string	:=	"radp_ctle_adapt_cycle_window_6";
		adp_ctle_adapt_oneshot	:	string	:=	"radp_ctle_adapt_oneshot_1";
		adp_ctle_en	:	string	:=	"radp_ctle_disable";
		adp_ctle_eqz_1s_sel	:	string	:=	"radp_ctle_eqz_1s_sel_0";
		adp_ctle_force_spec_sign	:	string	:=	"radp_ctle_force_spec_sign_0";
		adp_ctle_hold_en	:	string	:=	"radp_ctle_not_held";
		adp_ctle_load	:	string	:=	"radp_ctle_load_0";
		adp_ctle_load_value	:	string	:=	"radp_ctle_load_value_0";
		adp_ctle_scale	:	string	:=	"radp_ctle_scale_0";
		adp_ctle_scale_en	:	string	:=	"radp_ctle_scale_en_0";
		adp_ctle_spec_sign	:	string	:=	"radp_ctle_spec_sign_0";
		adp_ctle_sweep_direction	:	string	:=	"radp_ctle_sweep_direction_1";
		adp_ctle_threshold	:	string	:=	"radp_ctle_threshold_0";
		adp_ctle_threshold_en	:	string	:=	"radp_ctle_threshold_en_0";
		adp_ctle_vref_polarity	:	string	:=	"radp_ctle_vref_polarity_0";
		adp_ctle_window	:	string	:=	"radp_ctle_window_0";
		adp_dfe_bw	:	string	:=	"radp_dfe_bw_3";
		adp_dfe_clkout_div_sel	:	string	:=	"radp_dfe_clkout_div_sel_0";
		adp_dfe_cycle	:	string	:=	"radp_dfe_cycle_6";
		adp_dfe_fltap_bypass	:	string	:=	"radp_dfe_fltap_bypass_0";
		adp_dfe_fltap_en	:	string	:=	"radp_dfe_fltap_disable";
		adp_dfe_fltap_hold_en	:	string	:=	"radp_dfe_fltap_not_held";
		adp_dfe_fltap_load	:	string	:=	"radp_dfe_fltap_load_0";
		adp_dfe_fltap_position	:	string	:=	"radp_dfe_fltap_position_0";
		adp_dfe_force_spec_sign	:	string	:=	"radp_dfe_force_spec_sign_0";
		adp_dfe_fxtap1	:	string	:=	"radp_dfe_fxtap1_0";
		adp_dfe_fxtap10	:	string	:=	"radp_dfe_fxtap10_0";
		adp_dfe_fxtap10_sgn	:	string	:=	"radp_dfe_fxtap10_sgn_0";
		adp_dfe_fxtap11	:	string	:=	"radp_dfe_fxtap11_0";
		adp_dfe_fxtap11_sgn	:	string	:=	"radp_dfe_fxtap11_sgn_0";
		adp_dfe_fxtap2	:	string	:=	"radp_dfe_fxtap2_0";
		adp_dfe_fxtap2_sgn	:	string	:=	"radp_dfe_fxtap2_sgn_0";
		adp_dfe_fxtap3	:	string	:=	"radp_dfe_fxtap3_0";
		adp_dfe_fxtap3_sgn	:	string	:=	"radp_dfe_fxtap3_sgn_0";
		adp_dfe_fxtap4	:	string	:=	"radp_dfe_fxtap4_0";
		adp_dfe_fxtap4_sgn	:	string	:=	"radp_dfe_fxtap4_sgn_0";
		adp_dfe_fxtap5	:	string	:=	"radp_dfe_fxtap5_0";
		adp_dfe_fxtap5_sgn	:	string	:=	"radp_dfe_fxtap5_sgn_0";
		adp_dfe_fxtap6	:	string	:=	"radp_dfe_fxtap6_0";
		adp_dfe_fxtap6_sgn	:	string	:=	"radp_dfe_fxtap6_sgn_0";
		adp_dfe_fxtap7	:	string	:=	"radp_dfe_fxtap7_0";
		adp_dfe_fxtap7_sgn	:	string	:=	"radp_dfe_fxtap7_sgn_0";
		adp_dfe_fxtap8	:	string	:=	"radp_dfe_fxtap8_0";
		adp_dfe_fxtap8_sgn	:	string	:=	"radp_dfe_fxtap8_sgn_0";
		adp_dfe_fxtap9	:	string	:=	"radp_dfe_fxtap9_0";
		adp_dfe_fxtap9_sgn	:	string	:=	"radp_dfe_fxtap9_sgn_0";
		adp_dfe_fxtap_bypass	:	string	:=	"radp_dfe_fxtap_bypass_0";
		adp_dfe_fxtap_en	:	string	:=	"radp_dfe_fxtap_disable";
		adp_dfe_fxtap_hold_en	:	string	:=	"radp_dfe_fxtap_not_held";
		adp_dfe_fxtap_load	:	string	:=	"radp_dfe_fxtap_load_0";
		adp_dfe_mode	:	string	:=	"radp_dfe_mode_0";
		adp_dfe_spec_sign	:	string	:=	"radp_dfe_spec_sign_0";
		adp_dfe_vref_polarity	:	string	:=	"radp_dfe_vref_polarity_0";
		adp_force_freqlock	:	string	:=	"radp_force_freqlock_off";
		adp_frame_capture	:	string	:=	"radp_frame_capture_0";
		adp_frame_en	:	string	:=	"radp_frame_en_0";
		adp_frame_odi_sel	:	string	:=	"radp_frame_odi_sel_0";
		adp_frame_out_sel	:	string	:=	"radp_frame_out_sel_0";
		adp_lfeq_fb_sel	:	string	:=	"radp_lfeq_fb_sel_0";
		adp_mode	:	string	:=	"radp_mode_0";
		adp_odi_control_sel	:	string	:=	"radp_odi_control_sel_0";
		adp_onetime_dfe	:	string	:=	"radp_onetime_dfe_0";
		adp_spec_avg_window	:	string	:=	"radp_spec_avg_window_4";
		adp_spec_trans_filter	:	string	:=	"radp_spec_trans_filter_2";
		adp_status_sel	:	string	:=	"radp_status_sel_0";
		adp_vga_bypass	:	string	:=	"radp_vga_bypass_0";
		adp_vga_en	:	string	:=	"radp_vga_disable";
		adp_vga_load	:	string	:=	"radp_vga_load_0";
		adp_vga_polarity	:	string	:=	"radp_vga_polarity_0";
		adp_vga_sel	:	string	:=	"radp_vga_sel_0";
		adp_vga_sweep_direction	:	string	:=	"radp_vga_sweep_direction_1";
		adp_vga_threshold	:	string	:=	"radp_vga_threshold_4";
		adp_vref_bw	:	string	:=	"radp_vref_bw_1";
		adp_vref_bypass	:	string	:=	"radp_vref_bypass_0";
		adp_vref_cycle	:	string	:=	"radp_vref_cycle_6";
		adp_vref_dfe_spec_en	:	string	:=	"radp_vref_dfe_spec_en_0";
		adp_vref_en	:	string	:=	"radp_vref_disable";
		adp_vref_hold_en	:	string	:=	"radp_vref_not_held";
		adp_vref_load	:	string	:=	"radp_vref_load_0";
		adp_vref_polarity	:	string	:=	"radp_vref_polarity_0";
		adp_vref_sel	:	string	:=	"radp_vref_sel_21";
		adp_vref_vga_level	:	string	:=	"radp_vref_vga_level_13";
		datarate	:	string	:=	"0 bps";
		initial_settings	:	string	:=	"true";
		odi_count_threshold	:	string	:=	"rodi_count_threshold_0";
		odi_dfe_spec_en	:	string	:=	"rodi_dfe_spec_en_0";
		odi_en	:	string	:=	"rodi_en_0";
		odi_mode	:	string	:=	"rodi_mode_0";
		odi_rstn	:	string	:=	"rodi_rstn_0";
		odi_spec_sel	:	string	:=	"rodi_spec_sel_0";
		odi_start	:	string	:=	"rodi_start_0";
		odi_vref_sel	:	string	:=	"rodi_vref_sel_0";
		optimal	:	string	:=	"false";
		prot_mode	:	string	:=	"basic_rx";
		rrx_pcie_eqz	:	string	:=	"rrx_pcie_eqz_0";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode"
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		adapt_reset	:	in	std_logic	:=	'0';
		adapt_start	:	in	std_logic	:=	'0';
		deser_clk	:	in	std_logic	:=	'0';
		deser_data	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		deser_error	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		deser_odi	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		deser_odi_clk	:	in	std_logic	:=	'0';
		global_pipe_se	:	in	std_logic	:=	'0';
		i_rxpreset	:	in	std_logic_vector(2 downto 0)	:=	"000";
		radp_ctle_hold_en	:	in	std_logic	:=	'0';
		radp_ctle_patt_en	:	in	std_logic	:=	'0';
		radp_ctle_preset_sel	:	in	std_logic	:=	'0';
		radp_enable_max_lfeq_scale	:	in	std_logic	:=	'0';
		radp_lfeq_hold_en	:	in	std_logic	:=	'0';
		radp_vga_polarity	:	in	std_logic	:=	'0';
		rx_pllfreqlock	:	in	std_logic	:=	'0';
		scan_clk	:	in	std_logic	:=	'0';
		scan_in	:	in	std_logic_vector(9 downto 0)	:=	"0000000000";
		test_mode	:	in	std_logic	:=	'0';
		test_se	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		ctle_acgain_4s	:	out	std_logic_vector(27 downto 0)	:=	"0000000000000000000000000000";
		ctle_eqz_1s_sel	:	out	std_logic_vector(14 downto 0)	:=	"000000000000000";
		ctle_lfeq_fb_sel	:	out	std_logic_vector(6 downto 0)	:=	"0000000";
		dfe_adapt_en	:	out	std_logic	:=	'0';
		dfe_adp_clk	:	out	std_logic	:=	'0';
		dfe_fltap1	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		dfe_fltap1_sgn	:	out	std_logic	:=	'0';
		dfe_fltap2	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		dfe_fltap2_sgn	:	out	std_logic	:=	'0';
		dfe_fltap3	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		dfe_fltap3_sgn	:	out	std_logic	:=	'0';
		dfe_fltap4	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		dfe_fltap4_sgn	:	out	std_logic	:=	'0';
		dfe_fltap_bypdeser	:	out	std_logic	:=	'0';
		dfe_fltap_position	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		dfe_fxtap1	:	out	std_logic_vector(6 downto 0)	:=	"0000000";
		dfe_fxtap2	:	out	std_logic_vector(6 downto 0)	:=	"0000000";
		dfe_fxtap2_sgn	:	out	std_logic	:=	'0';
		dfe_fxtap3	:	out	std_logic_vector(6 downto 0)	:=	"0000000";
		dfe_fxtap3_sgn	:	out	std_logic	:=	'0';
		dfe_fxtap4	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		dfe_fxtap4_sgn	:	out	std_logic	:=	'0';
		dfe_fxtap5	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		dfe_fxtap5_sgn	:	out	std_logic	:=	'0';
		dfe_fxtap6	:	out	std_logic_vector(4 downto 0)	:=	"00000";
		dfe_fxtap6_sgn	:	out	std_logic	:=	'0';
		dfe_fxtap7	:	out	std_logic_vector(4 downto 0)	:=	"00000";
		dfe_fxtap7_sgn	:	out	std_logic	:=	'0';
		dfe_spec_disable	:	out	std_logic	:=	'0';
		dfe_spec_sign_sel	:	out	std_logic	:=	'0';
		dfe_vref_sign_sel	:	out	std_logic	:=	'0';
		odi_vref	:	out	std_logic_vector(4 downto 0)	:=	"00000";
		scan_out	:	out	std_logic_vector(9 downto 0)	:=	"0000000000";
		status_bus	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		vga_sel	:	out	std_logic_vector(6 downto 0)	:=	"0000000";
		vref_sel	:	out	std_logic_vector(4 downto 0)	:=	"00000"
	);
end component;

begin



inst : twentynm_hssi_pma_adaptation_encrypted
	generic map (
		-- Instance parameters
		adapt_dfe_control_sel	=>	adapt_dfe_control_sel,
		adapt_dfe_sel	=>	adapt_dfe_sel,
		adapt_mode	=>	adapt_mode,
		adapt_vga_sel	=>	adapt_vga_sel,
		adapt_vref_sel	=>	adapt_vref_sel,
		adp_1s_ctle_bypass	=>	adp_1s_ctle_bypass,
		adp_4s_ctle_bypass	=>	adp_4s_ctle_bypass,
		adp_adapt_control_sel	=>	adp_adapt_control_sel,
		adp_adapt_rstn	=>	adp_adapt_rstn,
		adp_adapt_start	=>	adp_adapt_start,
		adp_bist_auxpath_en	=>	adp_bist_auxpath_en,
		adp_bist_count_rstn	=>	adp_bist_count_rstn,
		adp_bist_datapath_en	=>	adp_bist_datapath_en,
		adp_bist_mode	=>	adp_bist_mode,
		adp_bist_odi_dfe_sel	=>	adp_bist_odi_dfe_sel,
		adp_bist_spec_en	=>	adp_bist_spec_en,
		adp_control_mux_bypass	=>	adp_control_mux_bypass,
		adp_ctle_acgain_4s	=>	adp_ctle_acgain_4s,
		adp_ctle_adapt_bw	=>	adp_ctle_adapt_bw,
		adp_ctle_adapt_cycle_window	=>	adp_ctle_adapt_cycle_window,
		adp_ctle_adapt_oneshot	=>	adp_ctle_adapt_oneshot,
		adp_ctle_en	=>	adp_ctle_en,
		adp_ctle_eqz_1s_sel	=>	adp_ctle_eqz_1s_sel,
		adp_ctle_force_spec_sign	=>	adp_ctle_force_spec_sign,
		adp_ctle_hold_en	=>	adp_ctle_hold_en,
		adp_ctle_load	=>	adp_ctle_load,
		adp_ctle_load_value	=>	adp_ctle_load_value,
		adp_ctle_scale	=>	adp_ctle_scale,
		adp_ctle_scale_en	=>	adp_ctle_scale_en,
		adp_ctle_spec_sign	=>	adp_ctle_spec_sign,
		adp_ctle_sweep_direction	=>	adp_ctle_sweep_direction,
		adp_ctle_threshold	=>	adp_ctle_threshold,
		adp_ctle_threshold_en	=>	adp_ctle_threshold_en,
		adp_ctle_vref_polarity	=>	adp_ctle_vref_polarity,
		adp_ctle_window	=>	adp_ctle_window,
		adp_dfe_bw	=>	adp_dfe_bw,
		adp_dfe_clkout_div_sel	=>	adp_dfe_clkout_div_sel,
		adp_dfe_cycle	=>	adp_dfe_cycle,
		adp_dfe_fltap_bypass	=>	adp_dfe_fltap_bypass,
		adp_dfe_fltap_en	=>	adp_dfe_fltap_en,
		adp_dfe_fltap_hold_en	=>	adp_dfe_fltap_hold_en,
		adp_dfe_fltap_load	=>	adp_dfe_fltap_load,
		adp_dfe_fltap_position	=>	adp_dfe_fltap_position,
		adp_dfe_force_spec_sign	=>	adp_dfe_force_spec_sign,
		adp_dfe_fxtap1	=>	adp_dfe_fxtap1,
		adp_dfe_fxtap10	=>	adp_dfe_fxtap10,
		adp_dfe_fxtap10_sgn	=>	adp_dfe_fxtap10_sgn,
		adp_dfe_fxtap11	=>	adp_dfe_fxtap11,
		adp_dfe_fxtap11_sgn	=>	adp_dfe_fxtap11_sgn,
		adp_dfe_fxtap2	=>	adp_dfe_fxtap2,
		adp_dfe_fxtap2_sgn	=>	adp_dfe_fxtap2_sgn,
		adp_dfe_fxtap3	=>	adp_dfe_fxtap3,
		adp_dfe_fxtap3_sgn	=>	adp_dfe_fxtap3_sgn,
		adp_dfe_fxtap4	=>	adp_dfe_fxtap4,
		adp_dfe_fxtap4_sgn	=>	adp_dfe_fxtap4_sgn,
		adp_dfe_fxtap5	=>	adp_dfe_fxtap5,
		adp_dfe_fxtap5_sgn	=>	adp_dfe_fxtap5_sgn,
		adp_dfe_fxtap6	=>	adp_dfe_fxtap6,
		adp_dfe_fxtap6_sgn	=>	adp_dfe_fxtap6_sgn,
		adp_dfe_fxtap7	=>	adp_dfe_fxtap7,
		adp_dfe_fxtap7_sgn	=>	adp_dfe_fxtap7_sgn,
		adp_dfe_fxtap8	=>	adp_dfe_fxtap8,
		adp_dfe_fxtap8_sgn	=>	adp_dfe_fxtap8_sgn,
		adp_dfe_fxtap9	=>	adp_dfe_fxtap9,
		adp_dfe_fxtap9_sgn	=>	adp_dfe_fxtap9_sgn,
		adp_dfe_fxtap_bypass	=>	adp_dfe_fxtap_bypass,
		adp_dfe_fxtap_en	=>	adp_dfe_fxtap_en,
		adp_dfe_fxtap_hold_en	=>	adp_dfe_fxtap_hold_en,
		adp_dfe_fxtap_load	=>	adp_dfe_fxtap_load,
		adp_dfe_mode	=>	adp_dfe_mode,
		adp_dfe_spec_sign	=>	adp_dfe_spec_sign,
		adp_dfe_vref_polarity	=>	adp_dfe_vref_polarity,
		adp_force_freqlock	=>	adp_force_freqlock,
		adp_frame_capture	=>	adp_frame_capture,
		adp_frame_en	=>	adp_frame_en,
		adp_frame_odi_sel	=>	adp_frame_odi_sel,
		adp_frame_out_sel	=>	adp_frame_out_sel,
		adp_lfeq_fb_sel	=>	adp_lfeq_fb_sel,
		adp_mode	=>	adp_mode,
		adp_odi_control_sel	=>	adp_odi_control_sel,
		adp_onetime_dfe	=>	adp_onetime_dfe,
		adp_spec_avg_window	=>	adp_spec_avg_window,
		adp_spec_trans_filter	=>	adp_spec_trans_filter,
		adp_status_sel	=>	adp_status_sel,
		adp_vga_bypass	=>	adp_vga_bypass,
		adp_vga_en	=>	adp_vga_en,
		adp_vga_load	=>	adp_vga_load,
		adp_vga_polarity	=>	adp_vga_polarity,
		adp_vga_sel	=>	adp_vga_sel,
		adp_vga_sweep_direction	=>	adp_vga_sweep_direction,
		adp_vga_threshold	=>	adp_vga_threshold,
		adp_vref_bw	=>	adp_vref_bw,
		adp_vref_bypass	=>	adp_vref_bypass,
		adp_vref_cycle	=>	adp_vref_cycle,
		adp_vref_dfe_spec_en	=>	adp_vref_dfe_spec_en,
		adp_vref_en	=>	adp_vref_en,
		adp_vref_hold_en	=>	adp_vref_hold_en,
		adp_vref_load	=>	adp_vref_load,
		adp_vref_polarity	=>	adp_vref_polarity,
		adp_vref_sel	=>	adp_vref_sel,
		adp_vref_vga_level	=>	adp_vref_vga_level,
		datarate	=>	datarate,
		initial_settings	=>	initial_settings,
		odi_count_threshold	=>	odi_count_threshold,
		odi_dfe_spec_en	=>	odi_dfe_spec_en,
		odi_en	=>	odi_en,
		odi_mode	=>	odi_mode,
		odi_rstn	=>	odi_rstn,
		odi_spec_sel	=>	odi_spec_sel,
		odi_start	=>	odi_start,
		odi_vref_sel	=>	odi_vref_sel,
		optimal	=>	optimal,
		prot_mode	=>	prot_mode,
		rrx_pcie_eqz	=>	rrx_pcie_eqz,
		silicon_rev	=>	silicon_rev,
		sup_mode	=>	sup_mode
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		adapt_reset	=>	adapt_reset,
		adapt_start	=>	adapt_start,
		deser_clk	=>	deser_clk,
		deser_data	=>	deser_data,
		deser_error	=>	deser_error,
		deser_odi	=>	deser_odi,
		deser_odi_clk	=>	deser_odi_clk,
		global_pipe_se	=>	global_pipe_se,
		i_rxpreset	=>	i_rxpreset,
		radp_ctle_hold_en	=>	radp_ctle_hold_en,
		radp_ctle_patt_en	=>	radp_ctle_patt_en,
		radp_ctle_preset_sel	=>	radp_ctle_preset_sel,
		radp_enable_max_lfeq_scale	=>	radp_enable_max_lfeq_scale,
		radp_lfeq_hold_en	=>	radp_lfeq_hold_en,
		radp_vga_polarity	=>	radp_vga_polarity,
		rx_pllfreqlock	=>	rx_pllfreqlock,
		scan_clk	=>	scan_clk,
		scan_in	=>	scan_in,
		test_mode	=>	test_mode,
		test_se	=>	test_se,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		ctle_acgain_4s	=>	ctle_acgain_4s,
		ctle_eqz_1s_sel	=>	ctle_eqz_1s_sel,
		ctle_lfeq_fb_sel	=>	ctle_lfeq_fb_sel,
		dfe_adapt_en	=>	dfe_adapt_en,
		dfe_adp_clk	=>	dfe_adp_clk,
		dfe_fltap1	=>	dfe_fltap1,
		dfe_fltap1_sgn	=>	dfe_fltap1_sgn,
		dfe_fltap2	=>	dfe_fltap2,
		dfe_fltap2_sgn	=>	dfe_fltap2_sgn,
		dfe_fltap3	=>	dfe_fltap3,
		dfe_fltap3_sgn	=>	dfe_fltap3_sgn,
		dfe_fltap4	=>	dfe_fltap4,
		dfe_fltap4_sgn	=>	dfe_fltap4_sgn,
		dfe_fltap_bypdeser	=>	dfe_fltap_bypdeser,
		dfe_fltap_position	=>	dfe_fltap_position,
		dfe_fxtap1	=>	dfe_fxtap1,
		dfe_fxtap2	=>	dfe_fxtap2,
		dfe_fxtap2_sgn	=>	dfe_fxtap2_sgn,
		dfe_fxtap3	=>	dfe_fxtap3,
		dfe_fxtap3_sgn	=>	dfe_fxtap3_sgn,
		dfe_fxtap4	=>	dfe_fxtap4,
		dfe_fxtap4_sgn	=>	dfe_fxtap4_sgn,
		dfe_fxtap5	=>	dfe_fxtap5,
		dfe_fxtap5_sgn	=>	dfe_fxtap5_sgn,
		dfe_fxtap6	=>	dfe_fxtap6,
		dfe_fxtap6_sgn	=>	dfe_fxtap6_sgn,
		dfe_fxtap7	=>	dfe_fxtap7,
		dfe_fxtap7_sgn	=>	dfe_fxtap7_sgn,
		dfe_spec_disable	=>	dfe_spec_disable,
		dfe_spec_sign_sel	=>	dfe_spec_sign_sel,
		dfe_vref_sign_sel	=>	dfe_vref_sign_sel,
		odi_vref	=>	odi_vref,
		scan_out	=>	scan_out,
		status_bus	=>	status_bus,
		vga_sel	=>	vga_sel,
		vref_sel	=>	vref_sel
	);
end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_pma_aux	is
	generic (
		-- Entity parameters
		dprio_base_addr	:	bit_vector	:=	B"000000000";
		dprio_broadcast_en	:	string	:=	"dprio_broadcast_en_csr_ctrl_en";
		dprio_cvp_mdio_dis	:	string	:=	"dprio_cvp_mdio_dis_csr_ctrl_en";
		dprio_force_mdio_dis	:	string	:=	"dprio_force_mdio_dis_csr_ctrl_en";
		dprio_power_iso_en	:	string	:=	"dprio_power_iso_en_csr_ctrl_en";
		initial_settings	:	string	:=	"true";
		pm_aux_adc_vref_trim	:	string	:=	"adc_vref_trim_4";
		pm_aux_atb_bgbyp	:	string	:=	"atb_bg_ref";
		pm_aux_atb_en	:	string	:=	"atb_global_disable";
		pm_aux_atb_mode	:	string	:=	"atb_default";
		pm_aux_atbcmp_pdb	:	string	:=	"atb_comp_power_down";
		pm_aux_atben0	:	string	:=	"atben0_disable";
		pm_aux_atben0_hssi	:	string	:=	"atb0_hssi_precomp_open";
		pm_aux_atben0_io	:	string	:=	"atb0_io_precomp_open";
		pm_aux_atben0_swap	:	string	:=	"atben0_swap_disable";
		pm_aux_atben1	:	string	:=	"atben1_disable";
		pm_aux_atben1_hssi	:	string	:=	"atb1_hssi_precomp_open";
		pm_aux_atben1_io	:	string	:=	"atb1_io_precomp_open";
		pm_aux_atben1_swap	:	string	:=	"atben1_swap_disable";
		pm_aux_bg_powerdown	:	string	:=	"pm_aux_bg_power_up";
		pm_aux_bypass_bg_voltage_to_iconstant	:	string	:=	"pm_aux_normal_operation_for_iconstant";
		pm_aux_bypass_bg_voltage_to_itrack	:	string	:=	"pm_aux_normal_operation_for_itrack";
		pm_aux_comp_minus	:	string	:=	"atb_comp_minus_disconnect";
		pm_aux_comp_plus	:	string	:=	"atb_comp_plus_disconnect";
		pm_aux_dac_atb_outsel	:	string	:=	"dac_atb_out_off";
		pm_aux_dac_data	:	bit_vector	:=	B"000000000000";
		pm_aux_dac_data_sel	:	string	:=	"dac_data_dprio";
		pm_aux_dac_dmcn	:	bit_vector	:=	B"11111111111100";
		pm_aux_dac_dmcp	:	bit_vector	:=	B"11111111111100";
		pm_aux_dac_lst	:	string	:=	"dac_atb1_disable";
		pm_aux_dac_neg_trigger	:	string	:=	"dac_pos_edge_trigger";
		pm_aux_dac_pdb	:	string	:=	"dac_power_down";
		pm_aux_dac_resetb	:	string	:=	"dac_reset_off";
		pm_aux_dac_tstbus_sel	:	string	:=	"dac_tst_0";
		pm_aux_dac_vouten	:	string	:=	"dac_vout_dis";
		pm_aux_dac_vref_sel	:	string	:=	"dac_fs_full";
		pm_aux_dac_vref_trim	:	string	:=	"dac_vref_trim_4";
		pm_aux_dftcmp_pdb	:	string	:=	"dft_comp_power_down";
		pm_aux_iconstant_opt	:	string	:=	"iconstant_opt_50u";
		pm_aux_impctrl_tstbus	:	string	:=	"pm_aux_impctrl_tstbus_sel0";
		pm_aux_itracking_opt	:	string	:=	"itracking_opt_50u";
		pm_aux_lower_limit	:	bit_vector	:=	B"000000000000";
		pm_aux_refclk_div	:	string	:=	"refclk_div_bypass";
		pm_aux_rx_cal_override_value	:	string	:=	"pm_aux_rx_cal_override_value0";
		pm_aux_rx_cal_override_value_enable	:	string	:=	"pm_aux_rx_cal_override_value_disable";
		pm_aux_rx_imp	:	string	:=	"pm_aux_rx_imp_48";
		pm_aux_sar_atb_insel	:	string	:=	"sar_atb_in_off";
		pm_aux_sar_cal_b10	:	string	:=	"sar_b10_cap_off";
		pm_aux_sar_cal_b11	:	string	:=	"sar_b11_cap_off";
		pm_aux_sar_cal_b5	:	string	:=	"sar_b5_cap_off";
		pm_aux_sar_cal_b6	:	string	:=	"sar_b6_cap_off";
		pm_aux_sar_cal_b7	:	string	:=	"sar_b7_cap_off";
		pm_aux_sar_cal_b8	:	string	:=	"sar_b8_cap_off";
		pm_aux_sar_cal_b9	:	string	:=	"sar_b9_cap_off";
		pm_aux_sar_cal_ctrl	:	string	:=	"sar_rambit_cal";
		pm_aux_sar_cal_mode	:	string	:=	"sar_normal_mode";
		pm_aux_sar_cal_refn	:	string	:=	"sar_refn_sw_off";
		pm_aux_sar_cal_refp	:	string	:=	"sar_refp_sw_off";
		pm_aux_sar_cal_top	:	string	:=	"sar_top_sw_off";
		pm_aux_sar_ckskew	:	string	:=	"sar_skew1";
		pm_aux_sar_cmp_curr	:	string	:=	"sar_cmp_curr11";
		pm_aux_sar_dmcn	:	bit_vector	:=	B"11111111111100";
		pm_aux_sar_dmcp	:	bit_vector	:=	B"11111111111100";
		pm_aux_sar_inbuf_byp	:	string	:=	"sar_inbuf_en";
		pm_aux_sar_insel	:	string	:=	"sar_input_off";
		pm_aux_sar_lowrate	:	string	:=	"sar_normal_rate";
		pm_aux_sar_lst	:	string	:=	"sar_atb1_disable";
		pm_aux_sar_pdb	:	string	:=	"sar_power_down";
		pm_aux_sar_resetb	:	string	:=	"sar_reset_off";
		pm_aux_sar_tstbus_sel	:	string	:=	"sar_tst_0";
		pm_aux_sar_vcm_ctrl	:	string	:=	"sar_vcm_900mv";
		pm_aux_sar_vcm_en	:	string	:=	"sar_vcm_on";
		pm_aux_sel_fusetrim_cramtrim_adc_dac	:	string	:=	"sel_cramtrim_to_adc_dac";
		pm_aux_termination_cal_ctrl	:	string	:=	"pm_aux_termination_cal_ctrl_0";
		pm_aux_test_counter	:	string	:=	"pm_aux_test_counter_disable";
		pm_aux_tstmux_statreg	:	string	:=	"pm_aux_tstmux_statreg_0";
		pm_aux_tx_cal_override_value	:	string	:=	"pm_aux_tx_cal_override_value0";
		pm_aux_tx_cal_override_value_enable	:	string	:=	"pm_aux_tx_cal_override_value_disable";
		pm_aux_tx_imp	:	string	:=	"pm_aux_tx_imp_48";
		pm_aux_upper_limit	:	bit_vector	:=	B"000000000000";
		pm_aux_vgen_pdb	:	string	:=	"vref_power_down";
		pm_aux_vgen_sel	:	bit_vector	:=	B"100000";
		pm_aux_vrefen_minus	:	string	:=	"vref_comp_minus_disconnect";
		pm_aux_vrefen_plus	:	string	:=	"vref_comp_plus_disconnect";
		pma_aux_clock_select	:	string	:=	"pma_aux_clock_select_clkusr";
		powerdown_mode	:	string	:=	"powerdown";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode";
		xdprio_aux_wrap_xdprio_aux_cfg_dprio_sel_core	:	string	:=	"avalon_access_from_uc";
		xdprio_aux_wrap_xdprio_aux_uc_channel_base_addr	:	bit_vector	:=	B"00000000";
		ximpctrl_pm_aux_impctrl_sel_high_code	:	string	:=	"pm_aux_impctrl_tx_sel_high";
		ximpctrl_pm_aux_impctrl_tx_enable_eos_det	:	string	:=	"pm_aux_impctrl_tx_disable_eos_det";
		ximpctrl_pm_aux_impctrl_tx_ovwr_ncal	:	string	:=	"pm_aux_impctrl_tx_ovwr_pcal";
		ximpctrl_pm_aux_impctrl_tx_ovwr_state	:	string	:=	"pm_aux_impctrl_tx_ovwr_state_disable";
		ximpctrl_pm_aux_impctrl_tx_ovwr_state50	:	string	:=	"pm_aux_impctrl_tx_ovwr_state50";
		ximpctrl_pm_aux_impctrl_txcode_sel	:	string	:=	"pm_aux_impctrl_txcode_sel0"
	);
	port (
		-- Entity ports
		dprio_addr	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		dprio_clk	:	in	std_logic	:=	'0';
		dprio_read	:	in	std_logic	:=	'0';
		dprio_rst_n	:	in	std_logic	:=	'0';
		dprio_write	:	in	std_logic	:=	'0';
		dprio_writedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		pld_scan_mode_n	:	in	std_logic	:=	'0';
		pld_scan_shift_n	:	in	std_logic	:=	'0';
		scan_clk_in_impctrl	:	in	std_logic	:=	'0';
		scan_in_impctrl	:	in	std_logic	:=	'0';
		dft_flag_down	:	out	std_logic	:=	'0';
		dft_flag_up	:	out	std_logic	:=	'0';
		scan_out_impctrl	:	out	std_logic	:=	'0';
		tstmux_out	:	out	std_logic_vector(7 downto 0)	:=	"00000000"
	);
end twentynm_hssi_pma_aux;

architecture behavior of twentynm_hssi_pma_aux	is

constant dprio_base_addr_int	:	integer	:=	bin2int(dprio_base_addr);
constant pm_aux_dac_data_int	:	integer	:=	bin2int(pm_aux_dac_data);
constant pm_aux_dac_dmcn_int	:	integer	:=	bin2int(pm_aux_dac_dmcn);
constant pm_aux_dac_dmcp_int	:	integer	:=	bin2int(pm_aux_dac_dmcp);
constant pm_aux_lower_limit_int	:	integer	:=	bin2int(pm_aux_lower_limit);
constant pm_aux_sar_dmcn_int	:	integer	:=	bin2int(pm_aux_sar_dmcn);
constant pm_aux_sar_dmcp_int	:	integer	:=	bin2int(pm_aux_sar_dmcp);
constant pm_aux_upper_limit_int	:	integer	:=	bin2int(pm_aux_upper_limit);
constant pm_aux_vgen_sel_int	:	integer	:=	bin2int(pm_aux_vgen_sel);
constant xdprio_aux_wrap_xdprio_aux_uc_channel_base_addr_int	:	integer	:=	bin2int(xdprio_aux_wrap_xdprio_aux_uc_channel_base_addr);



component	twentynm_hssi_pma_aux_encrypted
	generic (
		-- Architecture parameters
		dprio_base_addr	:	integer	:=	0;
		dprio_broadcast_en	:	string	:=	"dprio_broadcast_en_csr_ctrl_en";
		dprio_cvp_mdio_dis	:	string	:=	"dprio_cvp_mdio_dis_csr_ctrl_en";
		dprio_force_mdio_dis	:	string	:=	"dprio_force_mdio_dis_csr_ctrl_en";
		dprio_power_iso_en	:	string	:=	"dprio_power_iso_en_csr_ctrl_en";
		initial_settings	:	string	:=	"true";
		pm_aux_adc_vref_trim	:	string	:=	"adc_vref_trim_4";
		pm_aux_atb_bgbyp	:	string	:=	"atb_bg_ref";
		pm_aux_atb_en	:	string	:=	"atb_global_disable";
		pm_aux_atb_mode	:	string	:=	"atb_default";
		pm_aux_atbcmp_pdb	:	string	:=	"atb_comp_power_down";
		pm_aux_atben0	:	string	:=	"atben0_disable";
		pm_aux_atben0_hssi	:	string	:=	"atb0_hssi_precomp_open";
		pm_aux_atben0_io	:	string	:=	"atb0_io_precomp_open";
		pm_aux_atben0_swap	:	string	:=	"atben0_swap_disable";
		pm_aux_atben1	:	string	:=	"atben1_disable";
		pm_aux_atben1_hssi	:	string	:=	"atb1_hssi_precomp_open";
		pm_aux_atben1_io	:	string	:=	"atb1_io_precomp_open";
		pm_aux_atben1_swap	:	string	:=	"atben1_swap_disable";
		pm_aux_bg_powerdown	:	string	:=	"pm_aux_bg_power_up";
		pm_aux_bypass_bg_voltage_to_iconstant	:	string	:=	"pm_aux_normal_operation_for_iconstant";
		pm_aux_bypass_bg_voltage_to_itrack	:	string	:=	"pm_aux_normal_operation_for_itrack";
		pm_aux_comp_minus	:	string	:=	"atb_comp_minus_disconnect";
		pm_aux_comp_plus	:	string	:=	"atb_comp_plus_disconnect";
		pm_aux_dac_atb_outsel	:	string	:=	"dac_atb_out_off";
		pm_aux_dac_data	:	integer	:=	0;
		pm_aux_dac_data_sel	:	string	:=	"dac_data_dprio";
		pm_aux_dac_dmcn	:	integer	:=	16380;
		pm_aux_dac_dmcp	:	integer	:=	16380;
		pm_aux_dac_lst	:	string	:=	"dac_atb1_disable";
		pm_aux_dac_neg_trigger	:	string	:=	"dac_pos_edge_trigger";
		pm_aux_dac_pdb	:	string	:=	"dac_power_down";
		pm_aux_dac_resetb	:	string	:=	"dac_reset_off";
		pm_aux_dac_tstbus_sel	:	string	:=	"dac_tst_0";
		pm_aux_dac_vouten	:	string	:=	"dac_vout_dis";
		pm_aux_dac_vref_sel	:	string	:=	"dac_fs_full";
		pm_aux_dac_vref_trim	:	string	:=	"dac_vref_trim_4";
		pm_aux_dftcmp_pdb	:	string	:=	"dft_comp_power_down";
		pm_aux_iconstant_opt	:	string	:=	"iconstant_opt_50u";
		pm_aux_impctrl_tstbus	:	string	:=	"pm_aux_impctrl_tstbus_sel0";
		pm_aux_itracking_opt	:	string	:=	"itracking_opt_50u";
		pm_aux_lower_limit	:	integer	:=	0;
		pm_aux_refclk_div	:	string	:=	"refclk_div_bypass";
		pm_aux_rx_cal_override_value	:	string	:=	"pm_aux_rx_cal_override_value0";
		pm_aux_rx_cal_override_value_enable	:	string	:=	"pm_aux_rx_cal_override_value_disable";
		pm_aux_rx_imp	:	string	:=	"pm_aux_rx_imp_48";
		pm_aux_sar_atb_insel	:	string	:=	"sar_atb_in_off";
		pm_aux_sar_cal_b10	:	string	:=	"sar_b10_cap_off";
		pm_aux_sar_cal_b11	:	string	:=	"sar_b11_cap_off";
		pm_aux_sar_cal_b5	:	string	:=	"sar_b5_cap_off";
		pm_aux_sar_cal_b6	:	string	:=	"sar_b6_cap_off";
		pm_aux_sar_cal_b7	:	string	:=	"sar_b7_cap_off";
		pm_aux_sar_cal_b8	:	string	:=	"sar_b8_cap_off";
		pm_aux_sar_cal_b9	:	string	:=	"sar_b9_cap_off";
		pm_aux_sar_cal_ctrl	:	string	:=	"sar_rambit_cal";
		pm_aux_sar_cal_mode	:	string	:=	"sar_normal_mode";
		pm_aux_sar_cal_refn	:	string	:=	"sar_refn_sw_off";
		pm_aux_sar_cal_refp	:	string	:=	"sar_refp_sw_off";
		pm_aux_sar_cal_top	:	string	:=	"sar_top_sw_off";
		pm_aux_sar_ckskew	:	string	:=	"sar_skew1";
		pm_aux_sar_cmp_curr	:	string	:=	"sar_cmp_curr11";
		pm_aux_sar_dmcn	:	integer	:=	16380;
		pm_aux_sar_dmcp	:	integer	:=	16380;
		pm_aux_sar_inbuf_byp	:	string	:=	"sar_inbuf_en";
		pm_aux_sar_insel	:	string	:=	"sar_input_off";
		pm_aux_sar_lowrate	:	string	:=	"sar_normal_rate";
		pm_aux_sar_lst	:	string	:=	"sar_atb1_disable";
		pm_aux_sar_pdb	:	string	:=	"sar_power_down";
		pm_aux_sar_resetb	:	string	:=	"sar_reset_off";
		pm_aux_sar_tstbus_sel	:	string	:=	"sar_tst_0";
		pm_aux_sar_vcm_ctrl	:	string	:=	"sar_vcm_900mv";
		pm_aux_sar_vcm_en	:	string	:=	"sar_vcm_on";
		pm_aux_sel_fusetrim_cramtrim_adc_dac	:	string	:=	"sel_cramtrim_to_adc_dac";
		pm_aux_termination_cal_ctrl	:	string	:=	"pm_aux_termination_cal_ctrl_0";
		pm_aux_test_counter	:	string	:=	"pm_aux_test_counter_disable";
		pm_aux_tstmux_statreg	:	string	:=	"pm_aux_tstmux_statreg_0";
		pm_aux_tx_cal_override_value	:	string	:=	"pm_aux_tx_cal_override_value0";
		pm_aux_tx_cal_override_value_enable	:	string	:=	"pm_aux_tx_cal_override_value_disable";
		pm_aux_tx_imp	:	string	:=	"pm_aux_tx_imp_48";
		pm_aux_upper_limit	:	integer	:=	0;
		pm_aux_vgen_pdb	:	string	:=	"vref_power_down";
		pm_aux_vgen_sel	:	integer	:=	32;
		pm_aux_vrefen_minus	:	string	:=	"vref_comp_minus_disconnect";
		pm_aux_vrefen_plus	:	string	:=	"vref_comp_plus_disconnect";
		pma_aux_clock_select	:	string	:=	"pma_aux_clock_select_clkusr";
		powerdown_mode	:	string	:=	"powerdown";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode";
		xdprio_aux_wrap_xdprio_aux_cfg_dprio_sel_core	:	string	:=	"avalon_access_from_uc";
		xdprio_aux_wrap_xdprio_aux_uc_channel_base_addr	:	integer	:=	0;
		ximpctrl_pm_aux_impctrl_sel_high_code	:	string	:=	"pm_aux_impctrl_tx_sel_high";
		ximpctrl_pm_aux_impctrl_tx_enable_eos_det	:	string	:=	"pm_aux_impctrl_tx_disable_eos_det";
		ximpctrl_pm_aux_impctrl_tx_ovwr_ncal	:	string	:=	"pm_aux_impctrl_tx_ovwr_pcal";
		ximpctrl_pm_aux_impctrl_tx_ovwr_state	:	string	:=	"pm_aux_impctrl_tx_ovwr_state_disable";
		ximpctrl_pm_aux_impctrl_tx_ovwr_state50	:	string	:=	"pm_aux_impctrl_tx_ovwr_state50";
		ximpctrl_pm_aux_impctrl_txcode_sel	:	string	:=	"pm_aux_impctrl_txcode_sel0"
	);
	port (
		-- Architecture ports
		dprio_addr	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		dprio_clk	:	in	std_logic	:=	'0';
		dprio_read	:	in	std_logic	:=	'0';
		dprio_rst_n	:	in	std_logic	:=	'0';
		dprio_write	:	in	std_logic	:=	'0';
		dprio_writedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		pld_scan_mode_n	:	in	std_logic	:=	'0';
		pld_scan_shift_n	:	in	std_logic	:=	'0';
		scan_clk_in_impctrl	:	in	std_logic	:=	'0';
		scan_in_impctrl	:	in	std_logic	:=	'0';
		dft_flag_down	:	out	std_logic	:=	'0';
		dft_flag_up	:	out	std_logic	:=	'0';
		scan_out_impctrl	:	out	std_logic	:=	'0';
		tstmux_out	:	out	std_logic_vector(7 downto 0)	:=	"00000000"
	);
end component;

begin



inst : twentynm_hssi_pma_aux_encrypted
	generic map (
		-- Instance parameters
		dprio_base_addr	=>	dprio_base_addr_int,
		dprio_broadcast_en	=>	dprio_broadcast_en,
		dprio_cvp_mdio_dis	=>	dprio_cvp_mdio_dis,
		dprio_force_mdio_dis	=>	dprio_force_mdio_dis,
		dprio_power_iso_en	=>	dprio_power_iso_en,
		initial_settings	=>	initial_settings,
		pm_aux_adc_vref_trim	=>	pm_aux_adc_vref_trim,
		pm_aux_atb_bgbyp	=>	pm_aux_atb_bgbyp,
		pm_aux_atb_en	=>	pm_aux_atb_en,
		pm_aux_atb_mode	=>	pm_aux_atb_mode,
		pm_aux_atbcmp_pdb	=>	pm_aux_atbcmp_pdb,
		pm_aux_atben0	=>	pm_aux_atben0,
		pm_aux_atben0_hssi	=>	pm_aux_atben0_hssi,
		pm_aux_atben0_io	=>	pm_aux_atben0_io,
		pm_aux_atben0_swap	=>	pm_aux_atben0_swap,
		pm_aux_atben1	=>	pm_aux_atben1,
		pm_aux_atben1_hssi	=>	pm_aux_atben1_hssi,
		pm_aux_atben1_io	=>	pm_aux_atben1_io,
		pm_aux_atben1_swap	=>	pm_aux_atben1_swap,
		pm_aux_bg_powerdown	=>	pm_aux_bg_powerdown,
		pm_aux_bypass_bg_voltage_to_iconstant	=>	pm_aux_bypass_bg_voltage_to_iconstant,
		pm_aux_bypass_bg_voltage_to_itrack	=>	pm_aux_bypass_bg_voltage_to_itrack,
		pm_aux_comp_minus	=>	pm_aux_comp_minus,
		pm_aux_comp_plus	=>	pm_aux_comp_plus,
		pm_aux_dac_atb_outsel	=>	pm_aux_dac_atb_outsel,
		pm_aux_dac_data	=>	pm_aux_dac_data_int,
		pm_aux_dac_data_sel	=>	pm_aux_dac_data_sel,
		pm_aux_dac_dmcn	=>	pm_aux_dac_dmcn_int,
		pm_aux_dac_dmcp	=>	pm_aux_dac_dmcp_int,
		pm_aux_dac_lst	=>	pm_aux_dac_lst,
		pm_aux_dac_neg_trigger	=>	pm_aux_dac_neg_trigger,
		pm_aux_dac_pdb	=>	pm_aux_dac_pdb,
		pm_aux_dac_resetb	=>	pm_aux_dac_resetb,
		pm_aux_dac_tstbus_sel	=>	pm_aux_dac_tstbus_sel,
		pm_aux_dac_vouten	=>	pm_aux_dac_vouten,
		pm_aux_dac_vref_sel	=>	pm_aux_dac_vref_sel,
		pm_aux_dac_vref_trim	=>	pm_aux_dac_vref_trim,
		pm_aux_dftcmp_pdb	=>	pm_aux_dftcmp_pdb,
		pm_aux_iconstant_opt	=>	pm_aux_iconstant_opt,
		pm_aux_impctrl_tstbus	=>	pm_aux_impctrl_tstbus,
		pm_aux_itracking_opt	=>	pm_aux_itracking_opt,
		pm_aux_lower_limit	=>	pm_aux_lower_limit_int,
		pm_aux_refclk_div	=>	pm_aux_refclk_div,
		pm_aux_rx_cal_override_value	=>	pm_aux_rx_cal_override_value,
		pm_aux_rx_cal_override_value_enable	=>	pm_aux_rx_cal_override_value_enable,
		pm_aux_rx_imp	=>	pm_aux_rx_imp,
		pm_aux_sar_atb_insel	=>	pm_aux_sar_atb_insel,
		pm_aux_sar_cal_b10	=>	pm_aux_sar_cal_b10,
		pm_aux_sar_cal_b11	=>	pm_aux_sar_cal_b11,
		pm_aux_sar_cal_b5	=>	pm_aux_sar_cal_b5,
		pm_aux_sar_cal_b6	=>	pm_aux_sar_cal_b6,
		pm_aux_sar_cal_b7	=>	pm_aux_sar_cal_b7,
		pm_aux_sar_cal_b8	=>	pm_aux_sar_cal_b8,
		pm_aux_sar_cal_b9	=>	pm_aux_sar_cal_b9,
		pm_aux_sar_cal_ctrl	=>	pm_aux_sar_cal_ctrl,
		pm_aux_sar_cal_mode	=>	pm_aux_sar_cal_mode,
		pm_aux_sar_cal_refn	=>	pm_aux_sar_cal_refn,
		pm_aux_sar_cal_refp	=>	pm_aux_sar_cal_refp,
		pm_aux_sar_cal_top	=>	pm_aux_sar_cal_top,
		pm_aux_sar_ckskew	=>	pm_aux_sar_ckskew,
		pm_aux_sar_cmp_curr	=>	pm_aux_sar_cmp_curr,
		pm_aux_sar_dmcn	=>	pm_aux_sar_dmcn_int,
		pm_aux_sar_dmcp	=>	pm_aux_sar_dmcp_int,
		pm_aux_sar_inbuf_byp	=>	pm_aux_sar_inbuf_byp,
		pm_aux_sar_insel	=>	pm_aux_sar_insel,
		pm_aux_sar_lowrate	=>	pm_aux_sar_lowrate,
		pm_aux_sar_lst	=>	pm_aux_sar_lst,
		pm_aux_sar_pdb	=>	pm_aux_sar_pdb,
		pm_aux_sar_resetb	=>	pm_aux_sar_resetb,
		pm_aux_sar_tstbus_sel	=>	pm_aux_sar_tstbus_sel,
		pm_aux_sar_vcm_ctrl	=>	pm_aux_sar_vcm_ctrl,
		pm_aux_sar_vcm_en	=>	pm_aux_sar_vcm_en,
		pm_aux_sel_fusetrim_cramtrim_adc_dac	=>	pm_aux_sel_fusetrim_cramtrim_adc_dac,
		pm_aux_termination_cal_ctrl	=>	pm_aux_termination_cal_ctrl,
		pm_aux_test_counter	=>	pm_aux_test_counter,
		pm_aux_tstmux_statreg	=>	pm_aux_tstmux_statreg,
		pm_aux_tx_cal_override_value	=>	pm_aux_tx_cal_override_value,
		pm_aux_tx_cal_override_value_enable	=>	pm_aux_tx_cal_override_value_enable,
		pm_aux_tx_imp	=>	pm_aux_tx_imp,
		pm_aux_upper_limit	=>	pm_aux_upper_limit_int,
		pm_aux_vgen_pdb	=>	pm_aux_vgen_pdb,
		pm_aux_vgen_sel	=>	pm_aux_vgen_sel_int,
		pm_aux_vrefen_minus	=>	pm_aux_vrefen_minus,
		pm_aux_vrefen_plus	=>	pm_aux_vrefen_plus,
		pma_aux_clock_select	=>	pma_aux_clock_select,
		powerdown_mode	=>	powerdown_mode,
		silicon_rev	=>	silicon_rev,
		sup_mode	=>	sup_mode,
		xdprio_aux_wrap_xdprio_aux_cfg_dprio_sel_core	=>	xdprio_aux_wrap_xdprio_aux_cfg_dprio_sel_core,
		xdprio_aux_wrap_xdprio_aux_uc_channel_base_addr	=>	xdprio_aux_wrap_xdprio_aux_uc_channel_base_addr_int,
		ximpctrl_pm_aux_impctrl_sel_high_code	=>	ximpctrl_pm_aux_impctrl_sel_high_code,
		ximpctrl_pm_aux_impctrl_tx_enable_eos_det	=>	ximpctrl_pm_aux_impctrl_tx_enable_eos_det,
		ximpctrl_pm_aux_impctrl_tx_ovwr_ncal	=>	ximpctrl_pm_aux_impctrl_tx_ovwr_ncal,
		ximpctrl_pm_aux_impctrl_tx_ovwr_state	=>	ximpctrl_pm_aux_impctrl_tx_ovwr_state,
		ximpctrl_pm_aux_impctrl_tx_ovwr_state50	=>	ximpctrl_pm_aux_impctrl_tx_ovwr_state50,
		ximpctrl_pm_aux_impctrl_txcode_sel	=>	ximpctrl_pm_aux_impctrl_txcode_sel
	)
	port map (
		-- Instance ports
		dprio_addr	=>	dprio_addr,
		dprio_clk	=>	dprio_clk,
		dprio_read	=>	dprio_read,
		dprio_rst_n	=>	dprio_rst_n,
		dprio_write	=>	dprio_write,
		dprio_writedata	=>	dprio_writedata,
		pld_scan_mode_n	=>	pld_scan_mode_n,
		pld_scan_shift_n	=>	pld_scan_shift_n,
		scan_clk_in_impctrl	=>	scan_clk_in_impctrl,
		scan_in_impctrl	=>	scan_in_impctrl,
		dft_flag_down	=>	dft_flag_down,
		dft_flag_up	=>	dft_flag_up,
		scan_out_impctrl	=>	scan_out_impctrl,
		tstmux_out	=>	tstmux_out
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_pma_cdr_refclk_select_mux	is
	generic (
		-- Entity parameters
		cdr_clkin_scratch0_src	:	string	:=	"cdr_clkin_scratch0_src_refclk_iqclk";
		cdr_clkin_scratch1_src	:	string	:=	"cdr_clkin_scratch1_src_refclk_iqclk";
		cdr_clkin_scratch2_src	:	string	:=	"cdr_clkin_scratch2_src_refclk_iqclk";
		cdr_clkin_scratch3_src	:	string	:=	"cdr_clkin_scratch3_src_refclk_iqclk";
		cdr_clkin_scratch4_src	:	string	:=	"cdr_clkin_scratch4_src_refclk_iqclk";
		inclk0_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		inclk1_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		inclk2_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		inclk3_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		inclk4_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		powerdown_mode	:	string	:=	"powerdown";
		receiver_detect_src	:	string	:=	"iqclk_src";
		refclk_select	:	string	:=	"ref_iqclk0";
		silicon_rev	:	string	:=	"20nm5es";
		xmux_refclk_src	:	string	:=	"refclk_iqclk";
		xpm_iqref_mux_iqclk_sel	:	string	:=	"power_down";
		xpm_iqref_mux_scratch0_src	:	string	:=	"scratch0_power_down";
		xpm_iqref_mux_scratch1_src	:	string	:=	"scratch1_power_down";
		xpm_iqref_mux_scratch2_src	:	string	:=	"scratch2_power_down";
		xpm_iqref_mux_scratch3_src	:	string	:=	"scratch3_power_down";
		xpm_iqref_mux_scratch4_src	:	string	:=	"scratch4_power_down"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		core_refclk	:	in	std_logic	:=	'0';
		iqtxrxclk	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		ref_iqclk	:	in	std_logic_vector(11 downto 0)	:=	"000000000000";
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		refclk	:	out	std_logic	:=	'0';
		rx_det_clk	:	out	std_logic	:=	'0'
	);
end twentynm_hssi_pma_cdr_refclk_select_mux;

architecture behavior of twentynm_hssi_pma_cdr_refclk_select_mux	is




component	twentynm_hssi_pma_cdr_refclk_select_mux_encrypted
	generic (
		-- Architecture parameters
		cdr_clkin_scratch0_src	:	string	:=	"cdr_clkin_scratch0_src_refclk_iqclk";
		cdr_clkin_scratch1_src	:	string	:=	"cdr_clkin_scratch1_src_refclk_iqclk";
		cdr_clkin_scratch2_src	:	string	:=	"cdr_clkin_scratch2_src_refclk_iqclk";
		cdr_clkin_scratch3_src	:	string	:=	"cdr_clkin_scratch3_src_refclk_iqclk";
		cdr_clkin_scratch4_src	:	string	:=	"cdr_clkin_scratch4_src_refclk_iqclk";
		inclk0_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		inclk1_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		inclk2_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		inclk3_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		inclk4_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		powerdown_mode	:	string	:=	"powerdown";
		receiver_detect_src	:	string	:=	"iqclk_src";
		refclk_select	:	string	:=	"ref_iqclk0";
		silicon_rev	:	string	:=	"20nm5es";
		xmux_refclk_src	:	string	:=	"refclk_iqclk";
		xpm_iqref_mux_iqclk_sel	:	string	:=	"power_down";
		xpm_iqref_mux_scratch0_src	:	string	:=	"scratch0_power_down";
		xpm_iqref_mux_scratch1_src	:	string	:=	"scratch1_power_down";
		xpm_iqref_mux_scratch2_src	:	string	:=	"scratch2_power_down";
		xpm_iqref_mux_scratch3_src	:	string	:=	"scratch3_power_down";
		xpm_iqref_mux_scratch4_src	:	string	:=	"scratch4_power_down"
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		core_refclk	:	in	std_logic	:=	'0';
		iqtxrxclk	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		ref_iqclk	:	in	std_logic_vector(11 downto 0)	:=	"000000000000";
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		refclk	:	out	std_logic	:=	'0';
		rx_det_clk	:	out	std_logic	:=	'0'
	);
end component;

begin



inst : twentynm_hssi_pma_cdr_refclk_select_mux_encrypted
	generic map (
		-- Instance parameters
		cdr_clkin_scratch0_src	=>	cdr_clkin_scratch0_src,
		cdr_clkin_scratch1_src	=>	cdr_clkin_scratch1_src,
		cdr_clkin_scratch2_src	=>	cdr_clkin_scratch2_src,
		cdr_clkin_scratch3_src	=>	cdr_clkin_scratch3_src,
		cdr_clkin_scratch4_src	=>	cdr_clkin_scratch4_src,
		inclk0_logical_to_physical_mapping	=>	inclk0_logical_to_physical_mapping,
		inclk1_logical_to_physical_mapping	=>	inclk1_logical_to_physical_mapping,
		inclk2_logical_to_physical_mapping	=>	inclk2_logical_to_physical_mapping,
		inclk3_logical_to_physical_mapping	=>	inclk3_logical_to_physical_mapping,
		inclk4_logical_to_physical_mapping	=>	inclk4_logical_to_physical_mapping,
		powerdown_mode	=>	powerdown_mode,
		receiver_detect_src	=>	receiver_detect_src,
		refclk_select	=>	refclk_select,
		silicon_rev	=>	silicon_rev,
		xmux_refclk_src	=>	xmux_refclk_src,
		xpm_iqref_mux_iqclk_sel	=>	xpm_iqref_mux_iqclk_sel,
		xpm_iqref_mux_scratch0_src	=>	xpm_iqref_mux_scratch0_src,
		xpm_iqref_mux_scratch1_src	=>	xpm_iqref_mux_scratch1_src,
		xpm_iqref_mux_scratch2_src	=>	xpm_iqref_mux_scratch2_src,
		xpm_iqref_mux_scratch3_src	=>	xpm_iqref_mux_scratch3_src,
		xpm_iqref_mux_scratch4_src	=>	xpm_iqref_mux_scratch4_src
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		core_refclk	=>	core_refclk,
		iqtxrxclk	=>	iqtxrxclk,
		ref_iqclk	=>	ref_iqclk,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		refclk	=>	refclk,
		rx_det_clk	=>	rx_det_clk
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_pma_cgb_master	is
	generic (
		-- Entity parameters
		bonding_reset_enable	:	string	:=	"allow_bonding_reset";
		cgb_enable_iqtxrxclk	:	string	:=	"enable_iqtxrxclk";
		cgb_power_down	:	string	:=	"power_down_cgb";
		datarate	:	string	:=	"0 bps";
		dft_iqtxrxclk_control	:	string	:=	"dft_iqtxrxclk_drv_low";
		initial_settings	:	string	:=	"false";
		input_select	:	string	:=	"unused";
		input_select_gen3	:	string	:=	"unused";
		master_cgb_clock_control0	:	string	:=	"master_cgb_no_dft_control0";
		master_cgb_clock_control1	:	string	:=	"master_cgb_no_dft_control1";
		master_cgb_clock_control2	:	string	:=	"master_cgb_no_dft_control2";
		master_cgb_clock_control3	:	string	:=	"master_cgb_no_dft_control3";
		master_cgb_clock_control4	:	string	:=	"master_cgb_no_dft_control4";
		master_cgb_clock_control5	:	string	:=	"master_cgb_no_dft_control5";
		mcgb_high_perf_datarate_limit	:	string	:=	"000000000000000000000000000000000000";
		mcgb_high_perf_voltage	:	bit_vector	:=	B"000000000000";
		mcgb_low_power_datarate_limit	:	string	:=	"000000000000000000000000000000000000";
		mcgb_low_power_voltage	:	bit_vector	:=	B"000000000000";
		mcgb_mid_power_datarate_limit	:	string	:=	"000000000000000000000000000000000000";
		mcgb_mid_power_voltage	:	bit_vector	:=	B"000000000000";
		observe_cgb_clocks	:	string	:=	"observe_nothing";
		optimal	:	string	:=	"true";
		pcie_gen3_bitwidth	:	string	:=	"pciegen3_wide";
		powerdown_mode	:	string	:=	"powerup";
		prot_mode	:	string	:=	"unused";
		scratch0_x1_clock_src	:	string	:=	"unused";
		scratch1_x1_clock_src	:	string	:=	"unused";
		scratch2_x1_clock_src	:	string	:=	"unused";
		scratch3_x1_clock_src	:	string	:=	"unused";
		ser_mode	:	string	:=	"sixty_four_bit";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode";
		tx_ucontrol_en	:	string	:=	"disable";
		tx_ucontrol_pcie	:	string	:=	"gen1";
		tx_ucontrol_reset	:	string	:=	"disable";
		vccdreg_output	:	string	:=	"vccdreg_nominal";
		x1_clock_source_sel	:	string	:=	"fpll_top";
		x1_div_m_sel	:	string	:=	"divbypass"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		cgb_rstb	:	in	std_logic	:=	'0';
		clk_fpll_b	:	in	std_logic	:=	'0';
		clk_fpll_t	:	in	std_logic	:=	'0';
		clk_lc_b	:	in	std_logic	:=	'0';
		clk_lc_t	:	in	std_logic	:=	'0';
		clkb_fpll_b	:	in	std_logic	:=	'0';
		clkb_fpll_t	:	in	std_logic	:=	'0';
		clkb_lc_b	:	in	std_logic	:=	'0';
		clkb_lc_t	:	in	std_logic	:=	'0';
		pcie_sw	:	in	std_logic_vector(1 downto 0)	:=	"00";
		tx_bonding_rstb	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		cpulse_out_bus	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		mstcgb_core	:	out	std_logic_vector(1 downto 0)	:=	"00";
		pcie_sw_done	:	out	std_logic_vector(1 downto 0)	:=	"00";
		tx_iqtxrxclk_out	:	out	std_logic	:=	'0'
	);
end twentynm_hssi_pma_cgb_master;

architecture behavior of twentynm_hssi_pma_cgb_master	is

constant mcgb_high_perf_voltage_int	:	integer	:=	bin2int(mcgb_high_perf_voltage);
constant mcgb_low_power_voltage_int	:	integer	:=	bin2int(mcgb_low_power_voltage);
constant mcgb_mid_power_voltage_int	:	integer	:=	bin2int(mcgb_mid_power_voltage);



component	twentynm_hssi_pma_cgb_master_encrypted
	generic (
		-- Architecture parameters
		bonding_reset_enable	:	string	:=	"allow_bonding_reset";
		cgb_enable_iqtxrxclk	:	string	:=	"enable_iqtxrxclk";
		cgb_power_down	:	string	:=	"power_down_cgb";
		datarate	:	string	:=	"0 bps";
		dft_iqtxrxclk_control	:	string	:=	"dft_iqtxrxclk_drv_low";
		initial_settings	:	string	:=	"false";
		input_select	:	string	:=	"unused";
		input_select_gen3	:	string	:=	"unused";
		master_cgb_clock_control0	:	string	:=	"master_cgb_no_dft_control0";
		master_cgb_clock_control1	:	string	:=	"master_cgb_no_dft_control1";
		master_cgb_clock_control2	:	string	:=	"master_cgb_no_dft_control2";
		master_cgb_clock_control3	:	string	:=	"master_cgb_no_dft_control3";
		master_cgb_clock_control4	:	string	:=	"master_cgb_no_dft_control4";
		master_cgb_clock_control5	:	string	:=	"master_cgb_no_dft_control5";
		mcgb_high_perf_datarate_limit	:	string	:=	"000000000000000000000000000000000000";
		mcgb_high_perf_voltage	:	integer	:=	0;
		mcgb_low_power_datarate_limit	:	string	:=	"000000000000000000000000000000000000";
		mcgb_low_power_voltage	:	integer	:=	0;
		mcgb_mid_power_datarate_limit	:	string	:=	"000000000000000000000000000000000000";
		mcgb_mid_power_voltage	:	integer	:=	0;
		observe_cgb_clocks	:	string	:=	"observe_nothing";
		optimal	:	string	:=	"true";
		pcie_gen3_bitwidth	:	string	:=	"pciegen3_wide";
		powerdown_mode	:	string	:=	"powerup";
		prot_mode	:	string	:=	"unused";
		scratch0_x1_clock_src	:	string	:=	"unused";
		scratch1_x1_clock_src	:	string	:=	"unused";
		scratch2_x1_clock_src	:	string	:=	"unused";
		scratch3_x1_clock_src	:	string	:=	"unused";
		ser_mode	:	string	:=	"sixty_four_bit";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode";
		tx_ucontrol_en	:	string	:=	"disable";
		tx_ucontrol_pcie	:	string	:=	"gen1";
		tx_ucontrol_reset	:	string	:=	"disable";
		vccdreg_output	:	string	:=	"vccdreg_nominal";
		x1_clock_source_sel	:	string	:=	"fpll_top";
		x1_div_m_sel	:	string	:=	"divbypass"
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		cgb_rstb	:	in	std_logic	:=	'0';
		clk_fpll_b	:	in	std_logic	:=	'0';
		clk_fpll_t	:	in	std_logic	:=	'0';
		clk_lc_b	:	in	std_logic	:=	'0';
		clk_lc_t	:	in	std_logic	:=	'0';
		clkb_fpll_b	:	in	std_logic	:=	'0';
		clkb_fpll_t	:	in	std_logic	:=	'0';
		clkb_lc_b	:	in	std_logic	:=	'0';
		clkb_lc_t	:	in	std_logic	:=	'0';
		pcie_sw	:	in	std_logic_vector(1 downto 0)	:=	"00";
		tx_bonding_rstb	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		cpulse_out_bus	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		mstcgb_core	:	out	std_logic_vector(1 downto 0)	:=	"00";
		pcie_sw_done	:	out	std_logic_vector(1 downto 0)	:=	"00";
		tx_iqtxrxclk_out	:	out	std_logic	:=	'0'
	);
end component;

begin



inst : twentynm_hssi_pma_cgb_master_encrypted
	generic map (
		-- Instance parameters
		bonding_reset_enable	=>	bonding_reset_enable,
		cgb_enable_iqtxrxclk	=>	cgb_enable_iqtxrxclk,
		cgb_power_down	=>	cgb_power_down,
		datarate	=>	datarate,
		dft_iqtxrxclk_control	=>	dft_iqtxrxclk_control,
		initial_settings	=>	initial_settings,
		input_select	=>	input_select,
		input_select_gen3	=>	input_select_gen3,
		master_cgb_clock_control0	=>	master_cgb_clock_control0,
		master_cgb_clock_control1	=>	master_cgb_clock_control1,
		master_cgb_clock_control2	=>	master_cgb_clock_control2,
		master_cgb_clock_control3	=>	master_cgb_clock_control3,
		master_cgb_clock_control4	=>	master_cgb_clock_control4,
		master_cgb_clock_control5	=>	master_cgb_clock_control5,
		mcgb_high_perf_datarate_limit	=>	mcgb_high_perf_datarate_limit,
		mcgb_high_perf_voltage	=>	mcgb_high_perf_voltage_int,
		mcgb_low_power_datarate_limit	=>	mcgb_low_power_datarate_limit,
		mcgb_low_power_voltage	=>	mcgb_low_power_voltage_int,
		mcgb_mid_power_datarate_limit	=>	mcgb_mid_power_datarate_limit,
		mcgb_mid_power_voltage	=>	mcgb_mid_power_voltage_int,
		observe_cgb_clocks	=>	observe_cgb_clocks,
		optimal	=>	optimal,
		pcie_gen3_bitwidth	=>	pcie_gen3_bitwidth,
		powerdown_mode	=>	powerdown_mode,
		prot_mode	=>	prot_mode,
		scratch0_x1_clock_src	=>	scratch0_x1_clock_src,
		scratch1_x1_clock_src	=>	scratch1_x1_clock_src,
		scratch2_x1_clock_src	=>	scratch2_x1_clock_src,
		scratch3_x1_clock_src	=>	scratch3_x1_clock_src,
		ser_mode	=>	ser_mode,
		silicon_rev	=>	silicon_rev,
		sup_mode	=>	sup_mode,
		tx_ucontrol_en	=>	tx_ucontrol_en,
		tx_ucontrol_pcie	=>	tx_ucontrol_pcie,
		tx_ucontrol_reset	=>	tx_ucontrol_reset,
		vccdreg_output	=>	vccdreg_output,
		x1_clock_source_sel	=>	x1_clock_source_sel,
		x1_div_m_sel	=>	x1_div_m_sel
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		cgb_rstb	=>	cgb_rstb,
		clk_fpll_b	=>	clk_fpll_b,
		clk_fpll_t	=>	clk_fpll_t,
		clk_lc_b	=>	clk_lc_b,
		clk_lc_t	=>	clk_lc_t,
		clkb_fpll_b	=>	clkb_fpll_b,
		clkb_fpll_t	=>	clkb_fpll_t,
		clkb_lc_b	=>	clkb_lc_b,
		clkb_lc_t	=>	clkb_lc_t,
		pcie_sw	=>	pcie_sw,
		tx_bonding_rstb	=>	tx_bonding_rstb,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		cpulse_out_bus	=>	cpulse_out_bus,
		mstcgb_core	=>	mstcgb_core,
		pcie_sw_done	=>	pcie_sw_done,
		tx_iqtxrxclk_out	=>	tx_iqtxrxclk_out
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_pma_channel_pll	is
	generic (
		-- Entity parameters
		analog_mode	:	string	:=	"user_custom";
		atb_select_control	:	string	:=	"atb_off";
		auto_reset_on	:	string	:=	"auto_reset_on";
		bandwidth_range_high	:	string	:=	"0 hz";
		bandwidth_range_low	:	string	:=	"0 hz";
		bbpd_data_pattern_filter_select	:	string	:=	"bbpd_data_pat_off";
		bw_sel	:	string	:=	"low";
		cal_vco_count_length	:	string	:=	"sel_8b_count";
		cdr_odi_select	:	string	:=	"sel_cdr";
		cdr_phaselock_mode	:	string	:=	"no_ignore_lock";
		cdr_powerdown_mode	:	string	:=	"power_down";
		cgb_div	:	integer	:=	1;
		chgpmp_current_dn_pd	:	string	:=	"cp_current_pd_dn_setting0";
		chgpmp_current_dn_trim	:	string	:=	"cp_current_trimming_dn_setting0";
		chgpmp_current_pd	:	string	:=	"cp_current_pd_setting0";
		chgpmp_current_pfd	:	string	:=	"cp_current_pfd_setting0";
		chgpmp_current_up_pd	:	string	:=	"cp_current_pd_up_setting0";
		chgpmp_current_up_trim	:	string	:=	"cp_current_trimming_up_setting0";
		chgpmp_dn_pd_trim_double	:	string	:=	"normal_dn_trim_current";
		chgpmp_replicate	:	string	:=	"false";
		chgpmp_testmode	:	string	:=	"cp_test_disable";
		chgpmp_up_pd_trim_double	:	string	:=	"normal_up_trim_current";
		chgpmp_vccreg	:	string	:=	"vreg_fw0";
		clklow_mux_select	:	string	:=	"clklow_mux_cdr_fbclk";
		datarate	:	string	:=	"0 bps";
		diag_loopback_enable	:	string	:=	"false";
		disable_up_dn	:	string	:=	"true";
		enable_idle_rx_channel_support	:	string	:=	"false";
		f_max_cmu_out_freq	:	string	:=	"000000000000000000000000000000000001";
		f_max_m_counter	:	string	:=	"000000000000000000000000000000000001";
		f_max_pfd	:	string	:=	"0 hz";
		f_max_ref	:	string	:=	"0 hz";
		f_max_vco	:	string	:=	"0 hz";
		f_min_gt_channel	:	string	:=	"0 hz";
		f_min_pfd	:	string	:=	"0 hz";
		f_min_ref	:	string	:=	"0 hz";
		f_min_vco	:	string	:=	"0 hz";
		fb_select	:	string	:=	"direct_fb";
		fref_clklow_div	:	integer	:=	1;
		fref_mux_select	:	string	:=	"fref_mux_cdr_refclk";
		gpon_lck2ref_control	:	string	:=	"gpon_lck2ref_off";
		initial_settings	:	string	:=	"false";
		iqclk_mux_sel	:	string	:=	"power_down";
		is_cascaded_pll	:	string	:=	"false";
		lck2ref_delay_control	:	string	:=	"lck2ref_delay_off";
		lf_resistor_pd	:	string	:=	"lf_pd_setting0";
		lf_resistor_pfd	:	string	:=	"lf_pfd_setting0";
		lf_ripple_cap	:	string	:=	"lf_no_ripple";
		loop_filter_bias_select	:	string	:=	"lpflt_bias_off";
		loopback_mode	:	string	:=	"loopback_disabled";
		lpd_counter	:	bit_vector	:=	B"00001";
		lpfd_counter	:	bit_vector	:=	B"00001";
		ltd_ltr_micro_controller_select	:	string	:=	"ltd_ltr_pcs";
		m_counter	:	integer	:=	16;
		n_counter	:	integer	:=	1;
		n_counter_scratch	:	bit_vector	:=	B"000001";
		optimal	:	string	:=	"true";
		output_clock_frequency	:	string	:=	"0 hz";
		pcie_gen	:	string	:=	"non_pcie";
		pd_fastlock_mode	:	string	:=	"false";
		pd_l_counter	:	integer	:=	1;
		pfd_l_counter	:	integer	:=	1;
		pm_speed_grade	:	string	:=	"e2";
		pma_width	:	integer	:=	8;
		position	:	string	:=	"position_unknown";
		power_mode	:	string	:=	"low_power";
		primary_use	:	string	:=	"cmu";
		prot_mode	:	string	:=	"unused";
		reference_clock_frequency	:	string	:=	"0 hz";
		requires_gt_capable_channel	:	string	:=	"false";
		reverse_serial_loopback	:	string	:=	"no_loopback";
		set_cdr_input_freq_range	:	bit_vector	:=	B"00000000";
		set_cdr_v2i_enable	:	string	:=	"true";
		set_cdr_vco_reset	:	string	:=	"false";
		set_cdr_vco_speed	:	bit_vector	:=	B"00001";
		set_cdr_vco_speed_fix	:	bit_vector	:=	B"00000000";
		set_cdr_vco_speed_pciegen3	:	string	:=	"cdr_vco_max_speedbin_pciegen3";
		side	:	string	:=	"side_unknown";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode";
		top_or_bottom	:	string	:=	"tb_unknown";
		tx_pll_prot_mode	:	string	:=	"txpll_unused";
		txpll_hclk_driver_enable	:	string	:=	"false";
		uc_cru_rstb	:	string	:=	"cdr_lf_reset_off";
		uc_ro_cal	:	string	:=	"uc_ro_cal_off";
		uc_ro_cal_status	:	string	:=	"uc_ro_cal_notdone";
		vco_freq	:	string	:=	"0 hz";
		vco_overrange_voltage	:	string	:=	"vco_overrange_off";
		vco_underrange_voltage	:	string	:=	"vco_underange_off"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		adapt_en	:	in	std_logic	:=	'0';
		atbsel	:	in	std_logic_vector(62 downto 0)	:=	"000000000000000000000000000000000000000000000000000000000000000";
		clk0_bbpd	:	in	std_logic	:=	'0';
		clk180_bbpd	:	in	std_logic	:=	'0';
		clk270_bbpd	:	in	std_logic	:=	'0';
		clk90_bbpd	:	in	std_logic	:=	'0';
		deven	:	in	std_logic	:=	'0';
		devenb	:	in	std_logic	:=	'0';
		dfe_test	:	in	std_logic	:=	'0';
		dodd	:	in	std_logic	:=	'0';
		doddb	:	in	std_logic	:=	'0';
		e270	:	in	std_logic	:=	'0';
		e270b	:	in	std_logic	:=	'0';
		e90	:	in	std_logic	:=	'0';
		e90b	:	in	std_logic	:=	'0';
		early_eios	:	in	std_logic	:=	'0';
		error_even	:	in	std_logic	:=	'0';
		error_evenb	:	in	std_logic	:=	'0';
		error_odd	:	in	std_logic	:=	'0';
		error_oddb	:	in	std_logic	:=	'0';
		fpll_test0	:	in	std_logic	:=	'0';
		fpll_test1	:	in	std_logic	:=	'0';
		iqtxrxclk	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		ltd_b	:	in	std_logic	:=	'0';
		ltr	:	in	std_logic	:=	'0';
		odi_clk	:	in	std_logic	:=	'0';
		odi_clkb	:	in	std_logic	:=	'0';
		pcie_sw_ret	:	in	std_logic_vector(1 downto 0)	:=	"00";
		ppm_lock	:	in	std_logic	:=	'0';
		refclk	:	in	std_logic	:=	'0';
		rst_n	:	in	std_logic	:=	'0';
		rx_deser_pclk_test	:	in	std_logic	:=	'0';
		rx_lpbkn	:	in	std_logic	:=	'0';
		rx_lpbkp	:	in	std_logic	:=	'0';
		rxp	:	in	std_logic	:=	'0';
		sd	:	in	std_logic	:=	'0';
		tx_ser_pclk_test	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		cdr_cnt_done	:	out	std_logic	:=	'0';
		cdr_lpbkdp	:	out	std_logic	:=	'0';
		cdr_lpbkp	:	out	std_logic	:=	'0';
		cdr_refclk_cal_out	:	out	std_logic_vector(11 downto 0)	:=	"000000000000";
		cdr_vco_cal_out	:	out	std_logic_vector(11 downto 0)	:=	"000000000000";
		clk0_des	:	out	std_logic	:=	'0';
		clk0_odi	:	out	std_logic	:=	'0';
		clk0_pd	:	out	std_logic	:=	'0';
		clk0_pfd	:	out	std_logic	:=	'0';
		clk180_des	:	out	std_logic	:=	'0';
		clk180_odi	:	out	std_logic	:=	'0';
		clk180_pd	:	out	std_logic	:=	'0';
		clk180_pfd	:	out	std_logic	:=	'0';
		clk270_des	:	out	std_logic	:=	'0';
		clk270_odi	:	out	std_logic	:=	'0';
		clk270_pd	:	out	std_logic	:=	'0';
		clk90_des	:	out	std_logic	:=	'0';
		clk90_odi	:	out	std_logic	:=	'0';
		clk90_pd	:	out	std_logic	:=	'0';
		clklow	:	out	std_logic	:=	'0';
		deven_des	:	out	std_logic	:=	'0';
		devenb_des	:	out	std_logic	:=	'0';
		dodd_des	:	out	std_logic	:=	'0';
		doddb_des	:	out	std_logic	:=	'0';
		error_even_des	:	out	std_logic	:=	'0';
		error_evenb_des	:	out	std_logic	:=	'0';
		error_odd_des	:	out	std_logic	:=	'0';
		error_oddb_des	:	out	std_logic	:=	'0';
		fref	:	out	std_logic	:=	'0';
		lock2ref	:	out	std_logic	:=	'0';
		overrange	:	out	std_logic	:=	'0';
		pfdmode_lock	:	out	std_logic	:=	'0';
		rlpbkdn	:	out	std_logic	:=	'0';
		rlpbkdp	:	out	std_logic	:=	'0';
		rlpbkn	:	out	std_logic	:=	'0';
		rlpbkp	:	out	std_logic	:=	'0';
		rx_signal_ok	:	out	std_logic	:=	'0';
		rxpll_lock	:	out	std_logic	:=	'0';
		tx_rlpbk	:	out	std_logic	:=	'0';
		underrange	:	out	std_logic	:=	'0';
		von_lp	:	out	std_logic	:=	'0';
		vop_lp	:	out	std_logic	:=	'0'
	);
end twentynm_hssi_pma_channel_pll;

architecture behavior of twentynm_hssi_pma_channel_pll	is

constant lpd_counter_int	:	integer	:=	bin2int(lpd_counter);
constant lpfd_counter_int	:	integer	:=	bin2int(lpfd_counter);
constant n_counter_scratch_int	:	integer	:=	bin2int(n_counter_scratch);
constant set_cdr_input_freq_range_int	:	integer	:=	bin2int(set_cdr_input_freq_range);
constant set_cdr_vco_speed_int	:	integer	:=	bin2int(set_cdr_vco_speed);
constant set_cdr_vco_speed_fix_int	:	integer	:=	bin2int(set_cdr_vco_speed_fix);

signal clk180_des_temp : std_logic;
signal clk0_des_temp : std_logic;


component	twentynm_hssi_pma_channel_pll_encrypted
	generic (
		-- Architecture parameters
		analog_mode	:	string	:=	"user_custom";
		atb_select_control	:	string	:=	"atb_off";
		auto_reset_on	:	string	:=	"auto_reset_on";
		bandwidth_range_high	:	string	:=	"0 hz";
		bandwidth_range_low	:	string	:=	"0 hz";
		bbpd_data_pattern_filter_select	:	string	:=	"bbpd_data_pat_off";
		bw_sel	:	string	:=	"low";
		cal_vco_count_length	:	string	:=	"sel_8b_count";
		cdr_odi_select	:	string	:=	"sel_cdr";
		cdr_phaselock_mode	:	string	:=	"no_ignore_lock";
		cdr_powerdown_mode	:	string	:=	"power_down";
		cgb_div	:	integer	:=	1;
		chgpmp_current_dn_pd	:	string	:=	"cp_current_pd_dn_setting0";
		chgpmp_current_dn_trim	:	string	:=	"cp_current_trimming_dn_setting0";
		chgpmp_current_pfd	:	string	:=	"cp_current_pfd_setting0";
		chgpmp_current_up_pd	:	string	:=	"cp_current_pd_up_setting0";
		chgpmp_current_up_trim	:	string	:=	"cp_current_trimming_up_setting0";
		chgpmp_dn_pd_trim_double	:	string	:=	"normal_dn_trim_current";
		chgpmp_replicate	:	string	:=	"false";
		chgpmp_testmode	:	string	:=	"cp_test_disable";
		chgpmp_up_pd_trim_double	:	string	:=	"normal_up_trim_current";
		chgpmp_vccreg	:	string	:=	"vreg_fw0";
		clklow_mux_select	:	string	:=	"clklow_mux_cdr_fbclk";
		datarate	:	string	:=	"0 bps";
		diag_loopback_enable	:	string	:=	"false";
		disable_up_dn	:	string	:=	"true";
		enable_idle_rx_channel_support	:	string	:=	"false";
		f_max_cmu_out_freq	:	string	:=	"000000000000000000000000000000000001";
		f_max_m_counter	:	string	:=	"000000000000000000000000000000000001";
		f_max_pfd	:	string	:=	"0 hz";
		f_max_ref	:	string	:=	"0 hz";
		f_max_vco	:	string	:=	"0 hz";
		f_min_gt_channel	:	string	:=	"0 hz";
		f_min_pfd	:	string	:=	"0 hz";
		f_min_ref	:	string	:=	"0 hz";
		f_min_vco	:	string	:=	"0 hz";
		fb_select	:	string	:=	"direct_fb";
		fref_clklow_div	:	integer	:=	1;
		fref_mux_select	:	string	:=	"fref_mux_cdr_refclk";
		gpon_lck2ref_control	:	string	:=	"gpon_lck2ref_off";
		initial_settings	:	string	:=	"false";
		iqclk_mux_sel	:	string	:=	"power_down";
		is_cascaded_pll	:	string	:=	"false";
		lck2ref_delay_control	:	string	:=	"lck2ref_delay_off";
		lf_resistor_pd	:	string	:=	"lf_pd_setting0";
		lf_resistor_pfd	:	string	:=	"lf_pfd_setting0";
		lf_ripple_cap	:	string	:=	"lf_no_ripple";
		loop_filter_bias_select	:	string	:=	"lpflt_bias_off";
		loopback_mode	:	string	:=	"loopback_disabled";
		lpd_counter	:	integer	:=	1;
		lpfd_counter	:	integer	:=	1;
		ltd_ltr_micro_controller_select	:	string	:=	"ltd_ltr_pcs";
		m_counter	:	integer	:=	16;
		n_counter	:	integer	:=	1;
		n_counter_scratch	:	integer	:=	1;
		optimal	:	string	:=	"true";
		output_clock_frequency	:	string	:=	"0 hz";
		pcie_gen	:	string	:=	"non_pcie";
		pd_fastlock_mode	:	string	:=	"false";
		pd_l_counter	:	integer	:=	1;
		pfd_l_counter	:	integer	:=	1;
		pm_speed_grade	:	string	:=	"e2";
		pma_width	:	integer	:=	8;
		position	:	string	:=	"position_unknown";
		power_mode	:	string	:=	"low_power";
		primary_use	:	string	:=	"cmu";
		prot_mode	:	string	:=	"unused";
		reference_clock_frequency	:	string	:=	"0 hz";
		requires_gt_capable_channel	:	string	:=	"false";
		reverse_serial_loopback	:	string	:=	"no_loopback";
		set_cdr_input_freq_range	:	integer	:=	0;
		set_cdr_v2i_enable	:	string	:=	"true";
		set_cdr_vco_reset	:	string	:=	"false";
		set_cdr_vco_speed	:	integer	:=	1;
		set_cdr_vco_speed_fix	:	integer	:=	0;
		set_cdr_vco_speed_pciegen3	:	string	:=	"cdr_vco_max_speedbin_pciegen3";
		side	:	string	:=	"side_unknown";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode";
		top_or_bottom	:	string	:=	"tb_unknown";
		tx_pll_prot_mode	:	string	:=	"txpll_unused";
		txpll_hclk_driver_enable	:	string	:=	"false";
		uc_cru_rstb	:	string	:=	"cdr_lf_reset_off";
		uc_ro_cal	:	string	:=	"uc_ro_cal_off";
		uc_ro_cal_status	:	string	:=	"uc_ro_cal_notdone";
		vco_freq	:	string	:=	"0 hz";
		vco_overrange_voltage	:	string	:=	"vco_overrange_off";
		vco_underrange_voltage	:	string	:=	"vco_underange_off"
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		adapt_en	:	in	std_logic	:=	'0';
		atbsel	:	in	std_logic_vector(62 downto 0)	:=	"000000000000000000000000000000000000000000000000000000000000000";
		clk0_bbpd	:	in	std_logic	:=	'0';
		clk180_bbpd	:	in	std_logic	:=	'0';
		clk270_bbpd	:	in	std_logic	:=	'0';
		clk90_bbpd	:	in	std_logic	:=	'0';
		deven	:	in	std_logic	:=	'0';
		devenb	:	in	std_logic	:=	'0';
		dfe_test	:	in	std_logic	:=	'0';
		dodd	:	in	std_logic	:=	'0';
		doddb	:	in	std_logic	:=	'0';
		e270	:	in	std_logic	:=	'0';
		e270b	:	in	std_logic	:=	'0';
		e90	:	in	std_logic	:=	'0';
		e90b	:	in	std_logic	:=	'0';
		early_eios	:	in	std_logic	:=	'0';
		error_even	:	in	std_logic	:=	'0';
		error_evenb	:	in	std_logic	:=	'0';
		error_odd	:	in	std_logic	:=	'0';
		error_oddb	:	in	std_logic	:=	'0';
		fpll_test0	:	in	std_logic	:=	'0';
		fpll_test1	:	in	std_logic	:=	'0';
		iqtxrxclk	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		ltd_b	:	in	std_logic	:=	'0';
		ltr	:	in	std_logic	:=	'0';
		odi_clk	:	in	std_logic	:=	'0';
		odi_clkb	:	in	std_logic	:=	'0';
		pcie_sw_ret	:	in	std_logic_vector(1 downto 0)	:=	"00";
		ppm_lock	:	in	std_logic	:=	'0';
		refclk	:	in	std_logic	:=	'0';
		rst_n	:	in	std_logic	:=	'0';
		rx_deser_pclk_test	:	in	std_logic	:=	'0';
		rx_lpbkn	:	in	std_logic	:=	'0';
		rx_lpbkp	:	in	std_logic	:=	'0';
		rxp	:	in	std_logic	:=	'0';
		sd	:	in	std_logic	:=	'0';
		tx_ser_pclk_test	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		cdr_cnt_done	:	out	std_logic	:=	'0';
		cdr_lpbkdp	:	out	std_logic	:=	'0';
		cdr_lpbkp	:	out	std_logic	:=	'0';
		cdr_refclk_cal_out	:	out	std_logic_vector(11 downto 0)	:=	"000000000000";
		cdr_vco_cal_out	:	out	std_logic_vector(11 downto 0)	:=	"000000000000";
		clk0_des	:	out	std_logic	:=	'0';
		clk0_odi	:	out	std_logic	:=	'0';
		clk0_pd	:	out	std_logic	:=	'0';
		clk0_pfd	:	out	std_logic	:=	'0';
		clk180_des	:	out	std_logic	:=	'0';
		clk180_odi	:	out	std_logic	:=	'0';
		clk180_pd	:	out	std_logic	:=	'0';
		clk180_pfd	:	out	std_logic	:=	'0';
		clk270_odi	:	out	std_logic	:=	'0';
		clk270_pd	:	out	std_logic	:=	'0';
		clk90_odi	:	out	std_logic	:=	'0';
		clk90_pd	:	out	std_logic	:=	'0';
		clklow	:	out	std_logic	:=	'0';
		deven_des	:	out	std_logic	:=	'0';
		devenb_des	:	out	std_logic	:=	'0';
		dodd_des	:	out	std_logic	:=	'0';
		doddb_des	:	out	std_logic	:=	'0';
		error_even_des	:	out	std_logic	:=	'0';
		error_evenb_des	:	out	std_logic	:=	'0';
		error_odd_des	:	out	std_logic	:=	'0';
		error_oddb_des	:	out	std_logic	:=	'0';
		fref	:	out	std_logic	:=	'0';
		lock2ref	:	out	std_logic	:=	'0';
		overrange	:	out	std_logic	:=	'0';
		pfdmode_lock	:	out	std_logic	:=	'0';
		rlpbkdn	:	out	std_logic	:=	'0';
		rlpbkdp	:	out	std_logic	:=	'0';
		rlpbkn	:	out	std_logic	:=	'0';
		rlpbkp	:	out	std_logic	:=	'0';
		rx_signal_ok	:	out	std_logic	:=	'0';
		rxpll_lock	:	out	std_logic	:=	'0';
		tx_rlpbk	:	out	std_logic	:=	'0';
		underrange	:	out	std_logic	:=	'0';
		von_lp	:	out	std_logic	:=	'0';
		vop_lp	:	out	std_logic	:=	'0'
	);
end component;

begin

clk270_des <= clk180_des_temp;
clk180_des <= clk180_des_temp;
clk90_des <= clk0_des_temp;
clk0_des <= clk0_des_temp;


inst : twentynm_hssi_pma_channel_pll_encrypted
	generic map (
		-- Instance parameters
		analog_mode	=>	analog_mode,
		atb_select_control	=>	atb_select_control,
		auto_reset_on	=>	auto_reset_on,
		bandwidth_range_high	=>	bandwidth_range_high,
		bandwidth_range_low	=>	bandwidth_range_low,
		bbpd_data_pattern_filter_select	=>	bbpd_data_pattern_filter_select,
		bw_sel	=>	bw_sel,
		cal_vco_count_length	=>	cal_vco_count_length,
		cdr_odi_select	=>	cdr_odi_select,
		cdr_phaselock_mode	=>	cdr_phaselock_mode,
		cdr_powerdown_mode	=>	cdr_powerdown_mode,
		cgb_div	=>	cgb_div,
		chgpmp_current_dn_pd	=>	chgpmp_current_dn_pd,
		chgpmp_current_dn_trim	=>	chgpmp_current_dn_trim,
		chgpmp_current_pfd	=>	chgpmp_current_pfd,
		chgpmp_current_up_pd	=>	chgpmp_current_up_pd,
		chgpmp_current_up_trim	=>	chgpmp_current_up_trim,
		chgpmp_dn_pd_trim_double	=>	chgpmp_dn_pd_trim_double,
		chgpmp_replicate	=>	chgpmp_replicate,
		chgpmp_testmode	=>	chgpmp_testmode,
		chgpmp_up_pd_trim_double	=>	chgpmp_up_pd_trim_double,
		chgpmp_vccreg	=>	chgpmp_vccreg,
		clklow_mux_select	=>	clklow_mux_select,
		datarate	=>	datarate,
		diag_loopback_enable	=>	diag_loopback_enable,
		disable_up_dn	=>	disable_up_dn,
		enable_idle_rx_channel_support	=>	enable_idle_rx_channel_support,
		f_max_cmu_out_freq	=>	f_max_cmu_out_freq,
		f_max_m_counter	=>	f_max_m_counter,
		f_max_pfd	=>	f_max_pfd,
		f_max_ref	=>	f_max_ref,
		f_max_vco	=>	f_max_vco,
		f_min_gt_channel	=>	f_min_gt_channel,
		f_min_pfd	=>	f_min_pfd,
		f_min_ref	=>	f_min_ref,
		f_min_vco	=>	f_min_vco,
		fb_select	=>	fb_select,
		fref_clklow_div	=>	fref_clklow_div,
		fref_mux_select	=>	fref_mux_select,
		gpon_lck2ref_control	=>	gpon_lck2ref_control,
		initial_settings	=>	initial_settings,
		iqclk_mux_sel	=>	iqclk_mux_sel,
		is_cascaded_pll	=>	is_cascaded_pll,
		lck2ref_delay_control	=>	lck2ref_delay_control,
		lf_resistor_pd	=>	lf_resistor_pd,
		lf_resistor_pfd	=>	lf_resistor_pfd,
		lf_ripple_cap	=>	lf_ripple_cap,
		loop_filter_bias_select	=>	loop_filter_bias_select,
		loopback_mode	=>	loopback_mode,
		lpd_counter	=>	lpd_counter_int,
		lpfd_counter	=>	lpfd_counter_int,
		ltd_ltr_micro_controller_select	=>	ltd_ltr_micro_controller_select,
		m_counter	=>	m_counter,
		n_counter	=>	n_counter,
		n_counter_scratch	=>	n_counter_scratch_int,
		optimal	=>	optimal,
		output_clock_frequency	=>	output_clock_frequency,
		pcie_gen	=>	pcie_gen,
		pd_fastlock_mode	=>	pd_fastlock_mode,
		pd_l_counter	=>	pd_l_counter,
		pfd_l_counter	=>	pfd_l_counter,
		pm_speed_grade	=>	pm_speed_grade,
		pma_width	=>	pma_width,
		position	=>	position,
		power_mode	=>	power_mode,
		primary_use	=>	primary_use,
		prot_mode	=>	prot_mode,
		reference_clock_frequency	=>	reference_clock_frequency,
		requires_gt_capable_channel	=>	requires_gt_capable_channel,
		reverse_serial_loopback	=>	reverse_serial_loopback,
		set_cdr_input_freq_range	=>	set_cdr_input_freq_range_int,
		set_cdr_v2i_enable	=>	set_cdr_v2i_enable,
		set_cdr_vco_reset	=>	set_cdr_vco_reset,
		set_cdr_vco_speed	=>	set_cdr_vco_speed_int,
		set_cdr_vco_speed_fix	=>	set_cdr_vco_speed_fix_int,
		set_cdr_vco_speed_pciegen3	=>	set_cdr_vco_speed_pciegen3,
		side	=>	side,
		silicon_rev	=>	silicon_rev,
		sup_mode	=>	sup_mode,
		top_or_bottom	=>	top_or_bottom,
		tx_pll_prot_mode	=>	tx_pll_prot_mode,
		txpll_hclk_driver_enable	=>	txpll_hclk_driver_enable,
		uc_cru_rstb	=>	uc_cru_rstb,
		uc_ro_cal	=>	uc_ro_cal,
		uc_ro_cal_status	=>	uc_ro_cal_status,
		vco_freq	=>	vco_freq,
		vco_overrange_voltage	=>	vco_overrange_voltage,
		vco_underrange_voltage	=>	vco_underrange_voltage
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		adapt_en	=>	adapt_en,
		atbsel	=>	atbsel,
		clk0_bbpd	=>	clk0_bbpd,
		clk180_bbpd	=>	clk180_bbpd,
		clk270_bbpd	=>	clk270_bbpd,
		clk90_bbpd	=>	clk90_bbpd,
		deven	=>	deven,
		devenb	=>	devenb,
		dfe_test	=>	dfe_test,
		dodd	=>	dodd,
		doddb	=>	doddb,
		e270	=>	e270,
		e270b	=>	e270b,
		e90	=>	e90,
		e90b	=>	e90b,
		early_eios	=>	early_eios,
		error_even	=>	error_even,
		error_evenb	=>	error_evenb,
		error_odd	=>	error_odd,
		error_oddb	=>	error_oddb,
		fpll_test0	=>	fpll_test0,
		fpll_test1	=>	fpll_test1,
		iqtxrxclk	=>	iqtxrxclk,
		ltd_b	=>	ltd_b,
		ltr	=>	ltr,
		odi_clk	=>	odi_clk,
		odi_clkb	=>	odi_clkb,
		pcie_sw_ret	=>	pcie_sw_ret,
		ppm_lock	=>	ppm_lock,
		refclk	=>	refclk,
		rst_n	=>	rst_n,
		rx_deser_pclk_test	=>	rx_deser_pclk_test,
		rx_lpbkn	=>	rx_lpbkn,
		rx_lpbkp	=>	rx_lpbkp,
		rxp	=>	rxp,
		sd	=>	sd,
		tx_ser_pclk_test	=>	tx_ser_pclk_test,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		cdr_cnt_done	=>	cdr_cnt_done,
		cdr_lpbkdp	=>	cdr_lpbkdp,
		cdr_lpbkp	=>	cdr_lpbkp,
		cdr_refclk_cal_out	=>	cdr_refclk_cal_out,
		cdr_vco_cal_out	=>	cdr_vco_cal_out,
		clk0_des	=>	clk0_des_temp,
		clk0_odi	=>	clk0_odi,
		clk0_pd	=>	clk0_pd,
		clk0_pfd	=>	clk0_pfd,
		clk180_des	=>	clk180_des_temp,
		clk180_odi	=>	clk180_odi,
		clk180_pd	=>	clk180_pd,
		clk180_pfd	=>	clk180_pfd,
		clk270_odi	=>	clk270_odi,
		clk270_pd	=>	clk270_pd,
		clk90_odi	=>	clk90_odi,
		clk90_pd	=>	clk90_pd,
		clklow	=>	clklow,
		deven_des	=>	deven_des,
		devenb_des	=>	devenb_des,
		dodd_des	=>	dodd_des,
		doddb_des	=>	doddb_des,
		error_even_des	=>	error_even_des,
		error_evenb_des	=>	error_evenb_des,
		error_odd_des	=>	error_odd_des,
		error_oddb_des	=>	error_oddb_des,
		fref	=>	fref,
		lock2ref	=>	lock2ref,
		overrange	=>	overrange,
		pfdmode_lock	=>	pfdmode_lock,
		rlpbkdn	=>	rlpbkdn,
		rlpbkdp	=>	rlpbkdp,
		rlpbkn	=>	rlpbkn,
		rlpbkp	=>	rlpbkp,
		rx_signal_ok	=>	rx_signal_ok,
		rxpll_lock	=>	rxpll_lock,
		tx_rlpbk	=>	tx_rlpbk,
		underrange	=>	underrange,
		von_lp	=>	von_lp,
		vop_lp	=>	vop_lp
	);
end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_pma_lc_refclk_select_mux	is
	generic (
		-- Entity parameters
		inclk0_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		inclk1_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		inclk2_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		inclk3_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		inclk4_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		powerdown_mode	:	string	:=	"powerup";
		refclk_select	:	string	:=	"ref_iqclk0";
		silicon_rev	:	string	:=	"20nm5es";
		xmux_lc_scratch0_src	:	string	:=	"scratch0_src_lvpecl";
		xmux_lc_scratch1_src	:	string	:=	"scratch1_src_lvpecl";
		xmux_lc_scratch2_src	:	string	:=	"scratch2_src_lvpecl";
		xmux_lc_scratch3_src	:	string	:=	"scratch3_src_lvpecl";
		xmux_lc_scratch4_src	:	string	:=	"scratch4_src_lvpecl";
		xmux_refclk_src	:	string	:=	"src_lvpecl";
		xpm_iqref_mux_iqclk_sel	:	string	:=	"power_down";
		xpm_iqref_mux_scratch0_src	:	string	:=	"scratch0_power_down";
		xpm_iqref_mux_scratch1_src	:	string	:=	"scratch1_power_down";
		xpm_iqref_mux_scratch2_src	:	string	:=	"scratch2_power_down";
		xpm_iqref_mux_scratch3_src	:	string	:=	"scratch3_power_down";
		xpm_iqref_mux_scratch4_src	:	string	:=	"scratch4_power_down"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		core_refclk	:	in	std_logic	:=	'0';
		cr_pdb	:	in	std_logic	:=	'0';
		iqtxrxclk	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		lvpecl_in	:	in	std_logic	:=	'0';
		ref_iqclk	:	in	std_logic_vector(11 downto 0)	:=	"000000000000";
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		refclk	:	out	std_logic	:=	'0'
	);
end twentynm_hssi_pma_lc_refclk_select_mux;

architecture behavior of twentynm_hssi_pma_lc_refclk_select_mux	is




component	twentynm_hssi_pma_lc_refclk_select_mux_encrypted
	generic (
		-- Architecture parameters
		inclk0_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		inclk1_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		inclk2_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		inclk3_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		inclk4_logical_to_physical_mapping	:	string	:=	"ref_iqclk0";
		powerdown_mode	:	string	:=	"powerup";
		refclk_select	:	string	:=	"ref_iqclk0";
		silicon_rev	:	string	:=	"20nm5es";
		xmux_lc_scratch0_src	:	string	:=	"scratch0_src_lvpecl";
		xmux_lc_scratch1_src	:	string	:=	"scratch1_src_lvpecl";
		xmux_lc_scratch2_src	:	string	:=	"scratch2_src_lvpecl";
		xmux_lc_scratch3_src	:	string	:=	"scratch3_src_lvpecl";
		xmux_lc_scratch4_src	:	string	:=	"scratch4_src_lvpecl";
		xmux_refclk_src	:	string	:=	"src_lvpecl";
		xpm_iqref_mux_iqclk_sel	:	string	:=	"power_down";
		xpm_iqref_mux_scratch0_src	:	string	:=	"scratch0_power_down";
		xpm_iqref_mux_scratch1_src	:	string	:=	"scratch1_power_down";
		xpm_iqref_mux_scratch2_src	:	string	:=	"scratch2_power_down";
		xpm_iqref_mux_scratch3_src	:	string	:=	"scratch3_power_down";
		xpm_iqref_mux_scratch4_src	:	string	:=	"scratch4_power_down"
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		core_refclk	:	in	std_logic	:=	'0';
		cr_pdb	:	in	std_logic	:=	'0';
		iqtxrxclk	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		lvpecl_in	:	in	std_logic	:=	'0';
		ref_iqclk	:	in	std_logic_vector(11 downto 0)	:=	"000000000000";
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		refclk	:	out	std_logic	:=	'0'
	);
end component;

begin



inst : twentynm_hssi_pma_lc_refclk_select_mux_encrypted
	generic map (
		-- Instance parameters
		inclk0_logical_to_physical_mapping	=>	inclk0_logical_to_physical_mapping,
		inclk1_logical_to_physical_mapping	=>	inclk1_logical_to_physical_mapping,
		inclk2_logical_to_physical_mapping	=>	inclk2_logical_to_physical_mapping,
		inclk3_logical_to_physical_mapping	=>	inclk3_logical_to_physical_mapping,
		inclk4_logical_to_physical_mapping	=>	inclk4_logical_to_physical_mapping,
		powerdown_mode	=>	powerdown_mode,
		refclk_select	=>	refclk_select,
		silicon_rev	=>	silicon_rev,
		xmux_lc_scratch0_src	=>	xmux_lc_scratch0_src,
		xmux_lc_scratch1_src	=>	xmux_lc_scratch1_src,
		xmux_lc_scratch2_src	=>	xmux_lc_scratch2_src,
		xmux_lc_scratch3_src	=>	xmux_lc_scratch3_src,
		xmux_lc_scratch4_src	=>	xmux_lc_scratch4_src,
		xmux_refclk_src	=>	xmux_refclk_src,
		xpm_iqref_mux_iqclk_sel	=>	xpm_iqref_mux_iqclk_sel,
		xpm_iqref_mux_scratch0_src	=>	xpm_iqref_mux_scratch0_src,
		xpm_iqref_mux_scratch1_src	=>	xpm_iqref_mux_scratch1_src,
		xpm_iqref_mux_scratch2_src	=>	xpm_iqref_mux_scratch2_src,
		xpm_iqref_mux_scratch3_src	=>	xpm_iqref_mux_scratch3_src,
		xpm_iqref_mux_scratch4_src	=>	xpm_iqref_mux_scratch4_src
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		core_refclk	=>	core_refclk,
		cr_pdb	=>	cr_pdb,
		iqtxrxclk	=>	iqtxrxclk,
		lvpecl_in	=>	lvpecl_in,
		ref_iqclk	=>	ref_iqclk,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		refclk	=>	refclk
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_pma_rx_buf	is
	generic (
		-- Entity parameters
		act_isource_disable	:	string	:=	"isrc_en";
		bodybias_enable	:	string	:=	"bodybias_en";
		bodybias_select	:	string	:=	"bodybias_sel1";
		bypass_eqz_stages_234	:	string	:=	"bypass_off";
		cdrclk_to_cgb	:	string	:=	"cdrclk_2cgb_dis";
		cgm_bias_disable	:	string	:=	"cgmbias_en";
		datarate	:	string	:=	"0 bps";
		diag_lp_en	:	string	:=	"dlp_off";
		eq_bw_sel	:	string	:=	"eq_bw_1";
		eq_dc_gain_trim	:	string	:=	"no_dc_gain";
		initial_settings	:	string	:=	"false";
		input_vcm_sel	:	string	:=	"high_vcm";
		iostandard	:	string	:=	"hssi_diffio";
		lfeq_enable	:	string	:=	"non_lfeq_mode";
		lfeq_zero_control	:	string	:=	"lfeq_setting_2";
		link	:	string	:=	"sr";
		link_rx	:	string	:=	"sr";
		loopback_modes	:	string	:=	"lpbk_disable";
		offset_cal_pd	:	string	:=	"eqz1_en";
		offset_cancellation_coarse	:	string	:=	"coarse_setting_00";
		offset_cancellation_ctrl	:	string	:=	"volt_0mv";
		offset_cancellation_fine	:	string	:=	"fine_setting_00";
		offset_pd	:	string	:=	"oc_en";
		one_stage_enable	:	string	:=	"non_s1_mode";
		optimal	:	string	:=	"true";
		pdb_rx	:	string	:=	"power_down_rx";
		pm_speed_grade	:	string	:=	"e2";
		pm_tx_rx_cvp_mode	:	string	:=	"cvp_off";
		pm_tx_rx_pcie_gen	:	string	:=	"non_pcie";
		pm_tx_rx_pcie_gen_bitwidth	:	string	:=	"pcie_gen3_32b";
		pm_tx_rx_testmux_select	:	string	:=	"setting0";
		power_mode	:	string	:=	"low_power";
		power_mode_rx	:	string	:=	"low_power";
		power_rail_eht	:	integer	:=	0;
		power_rail_er	:	integer	:=	0;
		prot_mode	:	string	:=	"basic_rx";
		qpi_enable	:	string	:=	"non_qpi_mode";
		refclk_en	:	string	:=	"enable";
		rx_atb_select	:	string	:=	"atb_disable";
		rx_refclk_divider	:	string	:=	"bypass_divider";
		rx_sel_bias_source	:	string	:=	"bias_vcmdrv";
		rx_vga_oc_en	:	string	:=	"vga_cal_off";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode";
		term_sel	:	string	:=	"r_r1";
		term_tri_enable	:	string	:=	"disable_tri";
		vccela_supply_voltage	:	string	:=	"vccela_1p1v";
		vcm_current_add	:	string	:=	"vcm_current_default";
		vcm_sel	:	string	:=	"vcm_setting_10";
		vga_bandwidth_select	:	string	:=	"vga_bw_1";
		xrx_path_analog_mode	:	string	:=	"user_custom";
		xrx_path_datarate	:	string	:=	"0 bps";
		xrx_path_datawidth	:	bit_vector	:=	B"00000000";
		xrx_path_gt_enabled	:	string	:=	"disable";
		xrx_path_initial_settings	:	string	:=	"false";
		xrx_path_jtag_hys	:	string	:=	"hys_increase_disable";
		xrx_path_jtag_lp	:	string	:=	"lp_off";
		xrx_path_optimal	:	string	:=	"true";
		xrx_path_pma_rx_divclk_hz	:	string	:=	"00000000000000000000000000000000";
		xrx_path_prot_mode	:	string	:=	"unused";
		xrx_path_sup_mode	:	string	:=	"user_mode";
		xrx_path_uc_cal_enable	:	string	:=	"rx_cal_off";
		xrx_path_uc_cru_rstb	:	string	:=	"cdr_lf_reset_off";
		xrx_path_uc_pcie_sw	:	string	:=	"uc_pcie_gen1";
		xrx_path_uc_rx_rstb	:	string	:=	"rx_reset_on"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		clk_divrx	:	in	std_logic	:=	'0';
		lpbkn	:	in	std_logic	:=	'0';
		lpbkp	:	in	std_logic	:=	'0';
		rx_qpi_pulldn	:	in	std_logic	:=	'0';
		rx_rstn	:	in	std_logic	:=	'0';
		rx_sel_b50	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		rxn	:	in	std_logic	:=	'0';
		rxp	:	in	std_logic	:=	'0';
		s_lpbk_b	:	in	std_logic	:=	'0';
		vcz	:	in	std_logic_vector(27 downto 0)	:=	"0000000000000000000000000000";
		vds_eqz_s1_set	:	in	std_logic_vector(14 downto 0)	:=	"000000000000000";
		vds_lfeqz_czero	:	in	std_logic_vector(1 downto 0)	:=	"00";
		vds_lfeqz_fb_set	:	in	std_logic_vector(6 downto 0)	:=	"0000000";
		vds_vga_set	:	in	std_logic_vector(6 downto 0)	:=	"0000000";
		vga_cm_bidir_in	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		inn	:	out	std_logic	:=	'0';
		inp	:	out	std_logic	:=	'0';
		outn	:	out	std_logic	:=	'0';
		outp	:	out	std_logic	:=	'0';
		pull_dn	:	out	std_logic	:=	'0';
		rdlpbkn	:	out	std_logic	:=	'0';
		rdlpbkp	:	out	std_logic	:=	'0';
		rx_refclk	:	out	std_logic	:=	'0';
		vga_cm_bidir_out	:	out	std_logic	:=	'0'
	);
end twentynm_hssi_pma_rx_buf;

architecture behavior of twentynm_hssi_pma_rx_buf	is

constant xrx_path_datawidth_int	:	integer	:=	bin2int(xrx_path_datawidth);



component	twentynm_hssi_pma_rx_buf_encrypted
	generic (
		-- Architecture parameters
		act_isource_disable	:	string	:=	"isrc_en";
		bodybias_enable	:	string	:=	"bodybias_en";
		bodybias_select	:	string	:=	"bodybias_sel1";
		bypass_eqz_stages_234	:	string	:=	"bypass_off";
		cdrclk_to_cgb	:	string	:=	"cdrclk_2cgb_dis";
		cgm_bias_disable	:	string	:=	"cgmbias_en";
		datarate	:	string	:=	"0 bps";
		diag_lp_en	:	string	:=	"dlp_off";
		eq_bw_sel	:	string	:=	"eq_bw_1";
		eq_dc_gain_trim	:	string	:=	"no_dc_gain";
		initial_settings	:	string	:=	"false";
		input_vcm_sel	:	string	:=	"high_vcm";
		iostandard	:	string	:=	"hssi_diffio";
		lfeq_enable	:	string	:=	"non_lfeq_mode";
		lfeq_zero_control	:	string	:=	"lfeq_setting_2";
		link	:	string	:=	"sr";
		link_rx	:	string	:=	"sr";
		loopback_modes	:	string	:=	"lpbk_disable";
		offset_cal_pd	:	string	:=	"eqz1_en";
		offset_cancellation_coarse	:	string	:=	"coarse_setting_00";
		offset_cancellation_ctrl	:	string	:=	"volt_0mv";
		offset_cancellation_fine	:	string	:=	"fine_setting_00";
		offset_pd	:	string	:=	"oc_en";
		one_stage_enable	:	string	:=	"non_s1_mode";
		optimal	:	string	:=	"true";
		pdb_rx	:	string	:=	"power_down_rx";
		pm_speed_grade	:	string	:=	"e2";
		pm_tx_rx_cvp_mode	:	string	:=	"cvp_off";
		pm_tx_rx_pcie_gen	:	string	:=	"non_pcie";
		pm_tx_rx_pcie_gen_bitwidth	:	string	:=	"pcie_gen3_32b";
		pm_tx_rx_testmux_select	:	string	:=	"setting0";
		power_mode	:	string	:=	"low_power";
		power_mode_rx	:	string	:=	"low_power";
		power_rail_eht	:	integer	:=	0;
		power_rail_er	:	integer	:=	0;
		prot_mode	:	string	:=	"basic_rx";
		qpi_enable	:	string	:=	"non_qpi_mode";
		refclk_en	:	string	:=	"enable";
		rx_atb_select	:	string	:=	"atb_disable";
		rx_refclk_divider	:	string	:=	"bypass_divider";
		rx_sel_bias_source	:	string	:=	"bias_vcmdrv";
		rx_vga_oc_en	:	string	:=	"vga_cal_off";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode";
		term_sel	:	string	:=	"r_r1";
		term_tri_enable	:	string	:=	"disable_tri";
		vccela_supply_voltage	:	string	:=	"vccela_1p1v";
		vcm_current_add	:	string	:=	"vcm_current_default";
		vcm_sel	:	string	:=	"vcm_setting_10";
		vga_bandwidth_select	:	string	:=	"vga_bw_1";
		xrx_path_analog_mode	:	string	:=	"user_custom";
		xrx_path_datarate	:	string	:=	"0 bps";
		xrx_path_datawidth	:	integer	:=	0;
		xrx_path_gt_enabled	:	string	:=	"disable";
		xrx_path_initial_settings	:	string	:=	"false";
		xrx_path_jtag_hys	:	string	:=	"hys_increase_disable";
		xrx_path_jtag_lp	:	string	:=	"lp_off";
		xrx_path_optimal	:	string	:=	"true";
		xrx_path_pma_rx_divclk_hz	:	string	:=	"00000000000000000000000000000000";
		xrx_path_prot_mode	:	string	:=	"unused";
		xrx_path_sup_mode	:	string	:=	"user_mode";
		xrx_path_uc_cal_enable	:	string	:=	"rx_cal_off";
		xrx_path_uc_cru_rstb	:	string	:=	"cdr_lf_reset_off";
		xrx_path_uc_pcie_sw	:	string	:=	"uc_pcie_gen1";
		xrx_path_uc_rx_rstb	:	string	:=	"rx_reset_on"
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		clk_divrx	:	in	std_logic	:=	'0';
		lpbkn	:	in	std_logic	:=	'0';
		lpbkp	:	in	std_logic	:=	'0';
		rx_qpi_pulldn	:	in	std_logic	:=	'0';
		rx_rstn	:	in	std_logic	:=	'0';
		rx_sel_b50	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		rxn	:	in	std_logic	:=	'0';
		rxp	:	in	std_logic	:=	'0';
		s_lpbk_b	:	in	std_logic	:=	'0';
		vcz	:	in	std_logic_vector(27 downto 0)	:=	"0000000000000000000000000000";
		vds_eqz_s1_set	:	in	std_logic_vector(14 downto 0)	:=	"000000000000000";
		vds_lfeqz_czero	:	in	std_logic_vector(1 downto 0)	:=	"00";
		vds_lfeqz_fb_set	:	in	std_logic_vector(6 downto 0)	:=	"0000000";
		vds_vga_set	:	in	std_logic_vector(6 downto 0)	:=	"0000000";
		vga_cm_bidir_in	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		inn	:	out	std_logic	:=	'0';
		inp	:	out	std_logic	:=	'0';
		outn	:	out	std_logic	:=	'0';
		outp	:	out	std_logic	:=	'0';
		pull_dn	:	out	std_logic	:=	'0';
		rdlpbkn	:	out	std_logic	:=	'0';
		rdlpbkp	:	out	std_logic	:=	'0';
		rx_refclk	:	out	std_logic	:=	'0';
		vga_cm_bidir_out	:	out	std_logic	:=	'0'
	);
end component;

begin



inst : twentynm_hssi_pma_rx_buf_encrypted
	generic map (
		-- Instance parameters
		act_isource_disable	=>	act_isource_disable,
		bodybias_enable	=>	bodybias_enable,
		bodybias_select	=>	bodybias_select,
		bypass_eqz_stages_234	=>	bypass_eqz_stages_234,
		cdrclk_to_cgb	=>	cdrclk_to_cgb,
		cgm_bias_disable	=>	cgm_bias_disable,
		datarate	=>	datarate,
		diag_lp_en	=>	diag_lp_en,
		eq_bw_sel	=>	eq_bw_sel,
		eq_dc_gain_trim	=>	eq_dc_gain_trim,
		initial_settings	=>	initial_settings,
		input_vcm_sel	=>	input_vcm_sel,
		iostandard	=>	iostandard,
		lfeq_enable	=>	lfeq_enable,
		lfeq_zero_control	=>	lfeq_zero_control,
		link	=>	link,
		link_rx	=>	link_rx,
		loopback_modes	=>	loopback_modes,
		offset_cal_pd	=>	offset_cal_pd,
		offset_cancellation_coarse	=>	offset_cancellation_coarse,
		offset_cancellation_ctrl	=>	offset_cancellation_ctrl,
		offset_cancellation_fine	=>	offset_cancellation_fine,
		offset_pd	=>	offset_pd,
		one_stage_enable	=>	one_stage_enable,
		optimal	=>	optimal,
		pdb_rx	=>	pdb_rx,
		pm_speed_grade	=>	pm_speed_grade,
		pm_tx_rx_cvp_mode	=>	pm_tx_rx_cvp_mode,
		pm_tx_rx_pcie_gen	=>	pm_tx_rx_pcie_gen,
		pm_tx_rx_pcie_gen_bitwidth	=>	pm_tx_rx_pcie_gen_bitwidth,
		pm_tx_rx_testmux_select	=>	pm_tx_rx_testmux_select,
		power_mode	=>	power_mode,
		power_mode_rx	=>	power_mode_rx,
		power_rail_eht	=>	power_rail_eht,
		power_rail_er	=>	power_rail_er,
		prot_mode	=>	prot_mode,
		qpi_enable	=>	qpi_enable,
		refclk_en	=>	refclk_en,
		rx_atb_select	=>	rx_atb_select,
		rx_refclk_divider	=>	rx_refclk_divider,
		rx_sel_bias_source	=>	rx_sel_bias_source,
		rx_vga_oc_en	=>	rx_vga_oc_en,
		silicon_rev	=>	silicon_rev,
		sup_mode	=>	sup_mode,
		term_sel	=>	term_sel,
		term_tri_enable	=>	term_tri_enable,
		vccela_supply_voltage	=>	vccela_supply_voltage,
		vcm_current_add	=>	vcm_current_add,
		vcm_sel	=>	vcm_sel,
		vga_bandwidth_select	=>	vga_bandwidth_select,
		xrx_path_analog_mode	=>	xrx_path_analog_mode,
		xrx_path_datarate	=>	xrx_path_datarate,
		xrx_path_datawidth	=>	xrx_path_datawidth_int,
		xrx_path_gt_enabled	=>	xrx_path_gt_enabled,
		xrx_path_initial_settings	=>	xrx_path_initial_settings,
		xrx_path_jtag_hys	=>	xrx_path_jtag_hys,
		xrx_path_jtag_lp	=>	xrx_path_jtag_lp,
		xrx_path_optimal	=>	xrx_path_optimal,
		xrx_path_pma_rx_divclk_hz	=>	xrx_path_pma_rx_divclk_hz,
		xrx_path_prot_mode	=>	xrx_path_prot_mode,
		xrx_path_sup_mode	=>	xrx_path_sup_mode,
		xrx_path_uc_cal_enable	=>	xrx_path_uc_cal_enable,
		xrx_path_uc_cru_rstb	=>	xrx_path_uc_cru_rstb,
		xrx_path_uc_pcie_sw	=>	xrx_path_uc_pcie_sw,
		xrx_path_uc_rx_rstb	=>	xrx_path_uc_rx_rstb
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		clk_divrx	=>	clk_divrx,
		lpbkn	=>	lpbkn,
		lpbkp	=>	lpbkp,
		rx_qpi_pulldn	=>	rx_qpi_pulldn,
		rx_rstn	=>	rx_rstn,
		rx_sel_b50	=>	rx_sel_b50,
		rxn	=>	rxn,
		rxp	=>	rxp,
		s_lpbk_b	=>	s_lpbk_b,
		vcz	=>	vcz,
		vds_eqz_s1_set	=>	vds_eqz_s1_set,
		vds_lfeqz_czero	=>	vds_lfeqz_czero,
		vds_lfeqz_fb_set	=>	vds_lfeqz_fb_set,
		vds_vga_set	=>	vds_vga_set,
		vga_cm_bidir_in	=>	vga_cm_bidir_in,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		inn	=>	inn,
		inp	=>	inp,
		outn	=>	outn,
		outp	=>	outp,
		pull_dn	=>	pull_dn,
		rdlpbkn	=>	rdlpbkn,
		rdlpbkp	=>	rdlpbkp,
		rx_refclk	=>	rx_refclk,
		vga_cm_bidir_out	=>	vga_cm_bidir_out
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_pma_rx_deser	is
	generic (
		-- Entity parameters
		bitslip_bypass	:	string	:=	"bs_bypass_no";
		clkdiv_source	:	string	:=	"vco_bypass_normal";
		clkdivrx_user_mode	:	string	:=	"clkdivrx_user_disabled";
		datarate	:	string	:=	"0 bps";
		deser_factor	:	integer	:=	8;
		deser_powerdown	:	string	:=	"deser_power_up";
		force_adaptation_outputs	:	string	:=	"normal_outputs";
		force_clkdiv_for_testing	:	string	:=	"normal_clkdiv";
		optimal	:	string	:=	"true";
		pcie_gen	:	string	:=	"non_pcie";
		pcie_gen_bitwidth	:	string	:=	"pcie_gen3_32b";
		prot_mode	:	string	:=	"basic_rx";
		rst_n_adapt_odi	:	string	:=	"no_rst_adapt_odi";
		sdclk_enable	:	string	:=	"false";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode";
		tdr_mode	:	string	:=	"select_bbpd_data"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		adapt_en	:	in	std_logic	:=	'0';
		bitslip	:	in	std_logic	:=	'0';
		clk0	:	in	std_logic	:=	'0';
		clk0_odi	:	in	std_logic	:=	'0';
		clk180	:	in	std_logic	:=	'0';
		clk180_odi	:	in	std_logic	:=	'0';
		clk270	:	in	std_logic	:=	'0';
		clk90	:	in	std_logic	:=	'0';
		clklow	:	in	std_logic	:=	'0';
		deven	:	in	std_logic	:=	'0';
		deven_odi	:	in	std_logic	:=	'0';
		devenb	:	in	std_logic	:=	'0';
		devenb_odi	:	in	std_logic	:=	'0';
		dodd	:	in	std_logic	:=	'0';
		dodd_odi	:	in	std_logic	:=	'0';
		doddb	:	in	std_logic	:=	'0';
		doddb_odi	:	in	std_logic	:=	'0';
		error_even	:	in	std_logic	:=	'0';
		error_evenb	:	in	std_logic	:=	'0';
		error_odd	:	in	std_logic	:=	'0';
		error_oddb	:	in	std_logic	:=	'0';
		fref	:	in	std_logic	:=	'0';
		odi_en	:	in	std_logic	:=	'0';
		pcie_sw	:	in	std_logic_vector(1 downto 0)	:=	"00";
		pfdmode_lock	:	in	std_logic	:=	'0';
		rst_n	:	in	std_logic	:=	'0';
		tdr_en	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		adapt_clk	:	out	std_logic	:=	'0';
		clkdiv	:	out	std_logic	:=	'0';
		clkdiv_user	:	out	std_logic	:=	'0';
		clkdivrx_rx	:	out	std_logic	:=	'0';
		data	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		dout	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		error_deser	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		odi_clkout	:	out	std_logic	:=	'0';
		odi_dout	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		pcie_sw_ret	:	out	std_logic_vector(1 downto 0)	:=	"00";
		tstmx_deser	:	out	std_logic_vector(7 downto 0)	:=	"00000000"
	);
end twentynm_hssi_pma_rx_deser;

architecture behavior of twentynm_hssi_pma_rx_deser	is

function padder(s: string) return string is
	variable s0: string(1 to s'length) := s;
	variable RetVal: string(1 to 8);
	begin
		RetVal := (others => ' ');
		RetVal(s0'range) := s0;
		return RetVal;
end function padder;

signal silicon_rev_local : string(1 to 8) := (padder(silicon_rev));



signal clk0_temp : std_logic;
signal clk180_temp : std_logic;

component	twentynm_hssi_pma_rx_deser_encrypted
	generic (
		-- Architecture parameters
		bitslip_bypass	:	string	:=	"bs_bypass_no";
		clkdiv_source	:	string	:=	"vco_bypass_normal";
		clkdivrx_user_mode	:	string	:=	"clkdivrx_user_disabled";
		datarate	:	string	:=	"0 bps";
		deser_factor	:	integer	:=	8;
		deser_powerdown	:	string	:=	"deser_power_up";
		force_adaptation_outputs	:	string	:=	"normal_outputs";
		force_clkdiv_for_testing	:	string	:=	"normal_clkdiv";
		optimal	:	string	:=	"true";
		pcie_gen	:	string	:=	"non_pcie";
		pcie_gen_bitwidth	:	string	:=	"pcie_gen3_32b";
		prot_mode	:	string	:=	"basic_rx";
		rst_n_adapt_odi	:	string	:=	"no_rst_adapt_odi";
		sdclk_enable	:	string	:=	"false";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode";
		tdr_mode	:	string	:=	"select_bbpd_data"
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		adapt_en	:	in	std_logic	:=	'0';
		bitslip	:	in	std_logic	:=	'0';
		clk0	:	in	std_logic	:=	'0';
		clk0_odi	:	in	std_logic	:=	'0';
		clk180	:	in	std_logic	:=	'0';
		clk180_odi	:	in	std_logic	:=	'0';
		clklow	:	in	std_logic	:=	'0';
		deven	:	in	std_logic	:=	'0';
		deven_odi	:	in	std_logic	:=	'0';
		devenb	:	in	std_logic	:=	'0';
		devenb_odi	:	in	std_logic	:=	'0';
		dodd	:	in	std_logic	:=	'0';
		dodd_odi	:	in	std_logic	:=	'0';
		doddb	:	in	std_logic	:=	'0';
		doddb_odi	:	in	std_logic	:=	'0';
		error_even	:	in	std_logic	:=	'0';
		error_evenb	:	in	std_logic	:=	'0';
		error_odd	:	in	std_logic	:=	'0';
		error_oddb	:	in	std_logic	:=	'0';
		fref	:	in	std_logic	:=	'0';
		odi_en	:	in	std_logic	:=	'0';
		pcie_sw	:	in	std_logic_vector(1 downto 0)	:=	"00";
		pfdmode_lock	:	in	std_logic	:=	'0';
		rst_n	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		adapt_clk	:	out	std_logic	:=	'0';
		clkdiv	:	out	std_logic	:=	'0';
		clkdiv_user	:	out	std_logic	:=	'0';
		clkdivrx_rx	:	out	std_logic	:=	'0';
		data	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		dout	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		error_deser	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		odi_dout	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		pcie_sw_ret	:	out	std_logic_vector(1 downto 0)	:=	"00";
		tstmx_deser	:	out	std_logic_vector(7 downto 0)	:=	"00000000"
	);
end component;

begin


input_diffs:PROCESS(clk90,clk0,clk270,clk180)
BEGIN

CASE silicon_rev_local IS
	WHEN "20nm5es " => clk0_temp <= clk90;
	WHEN OTHERS => clk0_temp <= clk0;
END CASE;

CASE silicon_rev_local IS
	WHEN "20nm5es " => clk180_temp <= clk270;
	WHEN OTHERS => clk180_temp <= clk180;
END CASE;

END PROCESS input_diffs;

inst : twentynm_hssi_pma_rx_deser_encrypted
	generic map (
		-- Instance parameters
		bitslip_bypass	=>	bitslip_bypass,
		clkdiv_source	=>	clkdiv_source,
		clkdivrx_user_mode	=>	clkdivrx_user_mode,
		datarate	=>	datarate,
		deser_factor	=>	deser_factor,
		deser_powerdown	=>	deser_powerdown,
		force_adaptation_outputs	=>	force_adaptation_outputs,
		force_clkdiv_for_testing	=>	force_clkdiv_for_testing,
		optimal	=>	optimal,
		pcie_gen	=>	pcie_gen,
		pcie_gen_bitwidth	=>	pcie_gen_bitwidth,
		prot_mode	=>	prot_mode,
		rst_n_adapt_odi	=>	rst_n_adapt_odi,
		sdclk_enable	=>	sdclk_enable,
		silicon_rev	=>	silicon_rev,
		sup_mode	=>	sup_mode,
		tdr_mode	=>	tdr_mode
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		adapt_en	=>	adapt_en,
		bitslip	=>	bitslip,
		clk0	=>	clk0_temp,
		clk0_odi	=>	clk0_odi,
		clk180	=>	clk180_temp,
		clk180_odi	=>	clk180_odi,
		clklow	=>	clklow,
		deven	=>	deven,
		deven_odi	=>	deven_odi,
		devenb	=>	devenb,
		devenb_odi	=>	devenb_odi,
		dodd	=>	dodd,
		dodd_odi	=>	dodd_odi,
		doddb	=>	doddb,
		doddb_odi	=>	doddb_odi,
		error_even	=>	error_even,
		error_evenb	=>	error_evenb,
		error_odd	=>	error_odd,
		error_oddb	=>	error_oddb,
		fref	=>	fref,
		odi_en	=>	odi_en,
		pcie_sw	=>	pcie_sw,
		pfdmode_lock	=>	pfdmode_lock,
		rst_n	=>	rst_n,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		adapt_clk	=>	adapt_clk,
		clkdiv	=>	clkdiv,
		clkdiv_user	=>	clkdiv_user,
		clkdivrx_rx	=>	clkdivrx_rx,
		data	=>	data,
		dout	=>	dout,
		error_deser	=>	error_deser,
		odi_dout	=>	odi_dout,
		pcie_sw_ret	=>	pcie_sw_ret,
		tstmx_deser	=>	tstmx_deser
	);
end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_pma_rx_dfe	is
	generic (
		-- Entity parameters
		atb_select	:	string	:=	"atb_disable";
		datarate	:	string	:=	"0 bps";
		dft_en	:	string	:=	"dft_disable";
		initial_settings	:	string	:=	"true";
		oc_sa_adp1	:	bit_vector	:=	B"00000000";
		oc_sa_adp2	:	bit_vector	:=	B"00000000";
		oc_sa_c270	:	bit_vector	:=	B"00000000";
		oc_sa_c90	:	bit_vector	:=	B"00000000";
		oc_sa_d0c0	:	bit_vector	:=	B"00000000";
		oc_sa_d0c180	:	bit_vector	:=	B"00000000";
		oc_sa_d1c0	:	bit_vector	:=	B"00000000";
		oc_sa_d1c180	:	bit_vector	:=	B"00000000";
		optimal	:	string	:=	"true";
		pdb	:	string	:=	"dfe_enable";
		pdb_fixedtap	:	string	:=	"fixtap_dfe_powerdown";
		pdb_floattap	:	string	:=	"floattap_dfe_powerdown";
		pdb_fxtap4t7	:	string	:=	"fxtap4t7_powerdown";
		power_mode	:	string	:=	"low_power";
		prot_mode	:	string	:=	"basic_rx";
		sel_fltapstep_dec	:	string	:=	"fltap_step_no_dec";
		sel_fltapstep_inc	:	string	:=	"fltap_step_no_inc";
		sel_fxtapstep_dec	:	string	:=	"fxtap_step_no_dec";
		sel_fxtapstep_inc	:	string	:=	"fxtap_step_no_inc";
		sel_oc_en	:	string	:=	"off_canc_disable";
		sel_probe_tstmx	:	string	:=	"probe_tstmx_none";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode";
		uc_rx_dfe_cal	:	string	:=	"uc_rx_dfe_cal_off";
		uc_rx_dfe_cal_status	:	string	:=	"uc_rx_dfe_cal_notdone"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		adapt_en	:	in	std_logic	:=	'0';
		adp_clk	:	in	std_logic	:=	'0';
		clk0	:	in	std_logic	:=	'0';
		clk180	:	in	std_logic	:=	'0';
		clk270	:	in	std_logic	:=	'0';
		clk90	:	in	std_logic	:=	'0';
		dfe_fltap1_coeff	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		dfe_fltap1_sgn	:	in	std_logic	:=	'0';
		dfe_fltap2_coeff	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		dfe_fltap2_sgn	:	in	std_logic	:=	'0';
		dfe_fltap3_coeff	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		dfe_fltap3_sgn	:	in	std_logic	:=	'0';
		dfe_fltap4_coeff	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		dfe_fltap4_sgn	:	in	std_logic	:=	'0';
		dfe_fltap_bypdeser	:	in	std_logic	:=	'0';
		dfe_fltap_position	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		dfe_fxtap1_coeff	:	in	std_logic_vector(6 downto 0)	:=	"0000000";
		dfe_fxtap2_coeff	:	in	std_logic_vector(6 downto 0)	:=	"0000000";
		dfe_fxtap2_sgn	:	in	std_logic	:=	'0';
		dfe_fxtap3_coeff	:	in	std_logic_vector(6 downto 0)	:=	"0000000";
		dfe_fxtap3_sgn	:	in	std_logic	:=	'0';
		dfe_fxtap4_coeff	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		dfe_fxtap4_sgn	:	in	std_logic	:=	'0';
		dfe_fxtap5_coeff	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		dfe_fxtap5_sgn	:	in	std_logic	:=	'0';
		dfe_fxtap6_coeff	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		dfe_fxtap6_sgn	:	in	std_logic	:=	'0';
		dfe_fxtap7_coeff	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		dfe_fxtap7_sgn	:	in	std_logic	:=	'0';
		dfe_rstn	:	in	std_logic	:=	'0';
		dfe_spec_disable	:	in	std_logic	:=	'0';
		dfe_spec_sgn_sel	:	in	std_logic	:=	'0';
		dfe_vref_sgn_sel	:	in	std_logic	:=	'0';
		rxn	:	in	std_logic	:=	'0';
		rxp	:	in	std_logic	:=	'0';
		vga_vcm	:	in	std_logic	:=	'0';
		vref_level_coeff	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		clk0_bbpd	:	out	std_logic	:=	'0';
		clk180_bbpd	:	out	std_logic	:=	'0';
		clk270_bbpd	:	out	std_logic	:=	'0';
		clk90_bbpd	:	out	std_logic	:=	'0';
		deven	:	out	std_logic	:=	'0';
		devenb	:	out	std_logic	:=	'0';
		dfe_oc_tstmx	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		dodd	:	out	std_logic	:=	'0';
		doddb	:	out	std_logic	:=	'0';
		edge270	:	out	std_logic	:=	'0';
		edge270b	:	out	std_logic	:=	'0';
		edge90	:	out	std_logic	:=	'0';
		edge90b	:	out	std_logic	:=	'0';
		err_ev	:	out	std_logic	:=	'0';
		err_evb	:	out	std_logic	:=	'0';
		err_od	:	out	std_logic	:=	'0';
		err_odb	:	out	std_logic	:=	'0';
		spec_vrefh	:	out	std_logic	:=	'0';
		spec_vrefl	:	out	std_logic	:=	'0'
	);
end twentynm_hssi_pma_rx_dfe;

architecture behavior of twentynm_hssi_pma_rx_dfe	is

constant oc_sa_adp1_int	:	integer	:=	bin2int(oc_sa_adp1);
constant oc_sa_adp2_int	:	integer	:=	bin2int(oc_sa_adp2);
constant oc_sa_c270_int	:	integer	:=	bin2int(oc_sa_c270);
constant oc_sa_c90_int	:	integer	:=	bin2int(oc_sa_c90);
constant oc_sa_d0c0_int	:	integer	:=	bin2int(oc_sa_d0c0);
constant oc_sa_d0c180_int	:	integer	:=	bin2int(oc_sa_d0c180);
constant oc_sa_d1c0_int	:	integer	:=	bin2int(oc_sa_d1c0);
constant oc_sa_d1c180_int	:	integer	:=	bin2int(oc_sa_d1c180);



component	twentynm_hssi_pma_rx_dfe_encrypted
	generic (
		-- Architecture parameters
		atb_select	:	string	:=	"atb_disable";
		datarate	:	string	:=	"0 bps";
		dft_en	:	string	:=	"dft_disable";
		initial_settings	:	string	:=	"true";
		oc_sa_adp1	:	integer	:=	0;
		oc_sa_adp2	:	integer	:=	0;
		oc_sa_c270	:	integer	:=	0;
		oc_sa_c90	:	integer	:=	0;
		oc_sa_d0c0	:	integer	:=	0;
		oc_sa_d0c180	:	integer	:=	0;
		oc_sa_d1c0	:	integer	:=	0;
		oc_sa_d1c180	:	integer	:=	0;
		optimal	:	string	:=	"true";
		pdb	:	string	:=	"dfe_enable";
		pdb_fixedtap	:	string	:=	"fixtap_dfe_powerdown";
		pdb_floattap	:	string	:=	"floattap_dfe_powerdown";
		pdb_fxtap4t7	:	string	:=	"fxtap4t7_powerdown";
		power_mode	:	string	:=	"low_power";
		prot_mode	:	string	:=	"basic_rx";
		sel_fltapstep_dec	:	string	:=	"fltap_step_no_dec";
		sel_fltapstep_inc	:	string	:=	"fltap_step_no_inc";
		sel_fxtapstep_dec	:	string	:=	"fxtap_step_no_dec";
		sel_fxtapstep_inc	:	string	:=	"fxtap_step_no_inc";
		sel_oc_en	:	string	:=	"off_canc_disable";
		sel_probe_tstmx	:	string	:=	"probe_tstmx_none";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode";
		uc_rx_dfe_cal	:	string	:=	"uc_rx_dfe_cal_off";
		uc_rx_dfe_cal_status	:	string	:=	"uc_rx_dfe_cal_notdone"
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		adapt_en	:	in	std_logic	:=	'0';
		adp_clk	:	in	std_logic	:=	'0';
		clk0	:	in	std_logic	:=	'0';
		clk180	:	in	std_logic	:=	'0';
		clk270	:	in	std_logic	:=	'0';
		clk90	:	in	std_logic	:=	'0';
		dfe_fltap1_coeff	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		dfe_fltap1_sgn	:	in	std_logic	:=	'0';
		dfe_fltap2_coeff	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		dfe_fltap2_sgn	:	in	std_logic	:=	'0';
		dfe_fltap3_coeff	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		dfe_fltap3_sgn	:	in	std_logic	:=	'0';
		dfe_fltap4_coeff	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		dfe_fltap4_sgn	:	in	std_logic	:=	'0';
		dfe_fltap_bypdeser	:	in	std_logic	:=	'0';
		dfe_fltap_position	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		dfe_fxtap1_coeff	:	in	std_logic_vector(6 downto 0)	:=	"0000000";
		dfe_fxtap2_coeff	:	in	std_logic_vector(6 downto 0)	:=	"0000000";
		dfe_fxtap2_sgn	:	in	std_logic	:=	'0';
		dfe_fxtap3_coeff	:	in	std_logic_vector(6 downto 0)	:=	"0000000";
		dfe_fxtap3_sgn	:	in	std_logic	:=	'0';
		dfe_fxtap4_coeff	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		dfe_fxtap4_sgn	:	in	std_logic	:=	'0';
		dfe_fxtap5_coeff	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		dfe_fxtap5_sgn	:	in	std_logic	:=	'0';
		dfe_fxtap6_coeff	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		dfe_fxtap6_sgn	:	in	std_logic	:=	'0';
		dfe_fxtap7_coeff	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		dfe_fxtap7_sgn	:	in	std_logic	:=	'0';
		dfe_rstn	:	in	std_logic	:=	'0';
		dfe_spec_disable	:	in	std_logic	:=	'0';
		dfe_spec_sgn_sel	:	in	std_logic	:=	'0';
		dfe_vref_sgn_sel	:	in	std_logic	:=	'0';
		rxn	:	in	std_logic	:=	'0';
		rxp	:	in	std_logic	:=	'0';
		vga_vcm	:	in	std_logic	:=	'0';
		vref_level_coeff	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		clk0_bbpd	:	out	std_logic	:=	'0';
		clk180_bbpd	:	out	std_logic	:=	'0';
		clk270_bbpd	:	out	std_logic	:=	'0';
		clk90_bbpd	:	out	std_logic	:=	'0';
		deven	:	out	std_logic	:=	'0';
		devenb	:	out	std_logic	:=	'0';
		dfe_oc_tstmx	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		dodd	:	out	std_logic	:=	'0';
		doddb	:	out	std_logic	:=	'0';
		edge270	:	out	std_logic	:=	'0';
		edge270b	:	out	std_logic	:=	'0';
		edge90	:	out	std_logic	:=	'0';
		edge90b	:	out	std_logic	:=	'0';
		err_ev	:	out	std_logic	:=	'0';
		err_evb	:	out	std_logic	:=	'0';
		err_od	:	out	std_logic	:=	'0';
		err_odb	:	out	std_logic	:=	'0';
		spec_vrefh	:	out	std_logic	:=	'0';
		spec_vrefl	:	out	std_logic	:=	'0'
	);
end component;

begin



inst : twentynm_hssi_pma_rx_dfe_encrypted
	generic map (
		-- Instance parameters
		atb_select	=>	atb_select,
		datarate	=>	datarate,
		dft_en	=>	dft_en,
		initial_settings	=>	initial_settings,
		oc_sa_adp1	=>	oc_sa_adp1_int,
		oc_sa_adp2	=>	oc_sa_adp2_int,
		oc_sa_c270	=>	oc_sa_c270_int,
		oc_sa_c90	=>	oc_sa_c90_int,
		oc_sa_d0c0	=>	oc_sa_d0c0_int,
		oc_sa_d0c180	=>	oc_sa_d0c180_int,
		oc_sa_d1c0	=>	oc_sa_d1c0_int,
		oc_sa_d1c180	=>	oc_sa_d1c180_int,
		optimal	=>	optimal,
		pdb	=>	pdb,
		pdb_fixedtap	=>	pdb_fixedtap,
		pdb_floattap	=>	pdb_floattap,
		pdb_fxtap4t7	=>	pdb_fxtap4t7,
		power_mode	=>	power_mode,
		prot_mode	=>	prot_mode,
		sel_fltapstep_dec	=>	sel_fltapstep_dec,
		sel_fltapstep_inc	=>	sel_fltapstep_inc,
		sel_fxtapstep_dec	=>	sel_fxtapstep_dec,
		sel_fxtapstep_inc	=>	sel_fxtapstep_inc,
		sel_oc_en	=>	sel_oc_en,
		sel_probe_tstmx	=>	sel_probe_tstmx,
		silicon_rev	=>	silicon_rev,
		sup_mode	=>	sup_mode,
		uc_rx_dfe_cal	=>	uc_rx_dfe_cal,
		uc_rx_dfe_cal_status	=>	uc_rx_dfe_cal_status
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		adapt_en	=>	adapt_en,
		adp_clk	=>	adp_clk,
		clk0	=>	clk0,
		clk180	=>	clk180,
		clk270	=>	clk270,
		clk90	=>	clk90,
		dfe_fltap1_coeff	=>	dfe_fltap1_coeff,
		dfe_fltap1_sgn	=>	dfe_fltap1_sgn,
		dfe_fltap2_coeff	=>	dfe_fltap2_coeff,
		dfe_fltap2_sgn	=>	dfe_fltap2_sgn,
		dfe_fltap3_coeff	=>	dfe_fltap3_coeff,
		dfe_fltap3_sgn	=>	dfe_fltap3_sgn,
		dfe_fltap4_coeff	=>	dfe_fltap4_coeff,
		dfe_fltap4_sgn	=>	dfe_fltap4_sgn,
		dfe_fltap_bypdeser	=>	dfe_fltap_bypdeser,
		dfe_fltap_position	=>	dfe_fltap_position,
		dfe_fxtap1_coeff	=>	dfe_fxtap1_coeff,
		dfe_fxtap2_coeff	=>	dfe_fxtap2_coeff,
		dfe_fxtap2_sgn	=>	dfe_fxtap2_sgn,
		dfe_fxtap3_coeff	=>	dfe_fxtap3_coeff,
		dfe_fxtap3_sgn	=>	dfe_fxtap3_sgn,
		dfe_fxtap4_coeff	=>	dfe_fxtap4_coeff,
		dfe_fxtap4_sgn	=>	dfe_fxtap4_sgn,
		dfe_fxtap5_coeff	=>	dfe_fxtap5_coeff,
		dfe_fxtap5_sgn	=>	dfe_fxtap5_sgn,
		dfe_fxtap6_coeff	=>	dfe_fxtap6_coeff,
		dfe_fxtap6_sgn	=>	dfe_fxtap6_sgn,
		dfe_fxtap7_coeff	=>	dfe_fxtap7_coeff,
		dfe_fxtap7_sgn	=>	dfe_fxtap7_sgn,
		dfe_rstn	=>	dfe_rstn,
		dfe_spec_disable	=>	dfe_spec_disable,
		dfe_spec_sgn_sel	=>	dfe_spec_sgn_sel,
		dfe_vref_sgn_sel	=>	dfe_vref_sgn_sel,
		rxn	=>	rxn,
		rxp	=>	rxp,
		vga_vcm	=>	vga_vcm,
		vref_level_coeff	=>	vref_level_coeff,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		clk0_bbpd	=>	clk0_bbpd,
		clk180_bbpd	=>	clk180_bbpd,
		clk270_bbpd	=>	clk270_bbpd,
		clk90_bbpd	=>	clk90_bbpd,
		deven	=>	deven,
		devenb	=>	devenb,
		dfe_oc_tstmx	=>	dfe_oc_tstmx,
		dodd	=>	dodd,
		doddb	=>	doddb,
		edge270	=>	edge270,
		edge270b	=>	edge270b,
		edge90	=>	edge90,
		edge90b	=>	edge90b,
		err_ev	=>	err_ev,
		err_evb	=>	err_evb,
		err_od	=>	err_od,
		err_odb	=>	err_odb,
		spec_vrefh	=>	spec_vrefh,
		spec_vrefl	=>	spec_vrefl
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_pma_rx_odi	is
	generic (
		-- Entity parameters
		clk_dcd_bypass	:	string	:=	"no_bypass";
		datarate	:	string	:=	"0 bps";
		enable_odi	:	string	:=	"power_down_eye";
		initial_settings	:	string	:=	"false";
		invert_dfe_vref	:	string	:=	"no_inversion";
		monitor_bw_sel	:	string	:=	"bw_1";
		oc_sa_c0	:	bit_vector	:=	B"00000000";
		oc_sa_c180	:	bit_vector	:=	B"00000000";
		optimal	:	string	:=	"true";
		phase_steps_64_vs_128	:	string	:=	"phase_steps_64";
		phase_steps_sel	:	string	:=	"step40";
		power_mode	:	string	:=	"low_power";
		prot_mode	:	string	:=	"basic_rx";
		sel_oc_en	:	string	:=	"off_canc_disable";
		silicon_rev	:	string	:=	"20nm5es";
		step_ctrl_sel	:	string	:=	"feedback_mode";
		sup_mode	:	string	:=	"user_mode";
		v_vert_sel	:	string	:=	"plus";
		v_vert_threshold_scaling	:	string	:=	"scale_3";
		vert_threshold	:	string	:=	"vert_0"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		clk0	:	in	std_logic	:=	'0';
		clk180	:	in	std_logic	:=	'0';
		clk270	:	in	std_logic	:=	'0';
		clk90	:	in	std_logic	:=	'0';
		it50u	:	in	std_logic	:=	'0';
		it50u2	:	in	std_logic	:=	'0';
		it50u4	:	in	std_logic	:=	'0';
		odi_atb_sel	:	in	std_logic_vector(2 downto 0)	:=	"000";
		odi_dft_clr	:	in	std_logic	:=	'0';
		odi_latch_clk	:	in	std_logic	:=	'0';
		odi_shift_clk	:	in	std_logic	:=	'0';
		odi_shift_in	:	in	std_logic	:=	'0';
		rx_n	:	in	std_logic	:=	'0';
		rx_p	:	in	std_logic	:=	'0';
		rxn_sum	:	in	std_logic	:=	'0';
		rxp_sum	:	in	std_logic	:=	'0';
		spec_vrefh	:	in	std_logic	:=	'0';
		spec_vrefl	:	in	std_logic	:=	'0';
		vcm_vref	:	in	std_logic	:=	'0';
		vertical_fb	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		atb0	:	out	std_logic	:=	'0';
		atb1	:	out	std_logic	:=	'0';
		clk0_eye	:	out	std_logic	:=	'0';
		clk0_eye_lb	:	out	std_logic	:=	'0';
		clk180_eye	:	out	std_logic	:=	'0';
		clk180_eye_lb	:	out	std_logic	:=	'0';
		de_eye	:	out	std_logic	:=	'0';
		deb_eye	:	out	std_logic	:=	'0';
		do_eye	:	out	std_logic	:=	'0';
		dob_eye	:	out	std_logic	:=	'0';
		odi_en	:	out	std_logic	:=	'0';
		odi_oc_tstmx	:	out	std_logic_vector(1 downto 0)	:=	"00";
		tdr_en	:	out	std_logic	:=	'0';
		vref_sel_out	:	out	std_logic	:=	'0'
	);
end twentynm_hssi_pma_rx_odi;

architecture behavior of twentynm_hssi_pma_rx_odi	is

constant oc_sa_c0_int	:	integer	:=	bin2int(oc_sa_c0);
constant oc_sa_c180_int	:	integer	:=	bin2int(oc_sa_c180);



component	twentynm_hssi_pma_rx_odi_encrypted
	generic (
		-- Architecture parameters
		clk_dcd_bypass	:	string	:=	"no_bypass";
		datarate	:	string	:=	"0 bps";
		enable_odi	:	string	:=	"power_down_eye";
		initial_settings	:	string	:=	"false";
		invert_dfe_vref	:	string	:=	"no_inversion";
		monitor_bw_sel	:	string	:=	"bw_1";
		oc_sa_c0	:	integer	:=	0;
		oc_sa_c180	:	integer	:=	0;
		optimal	:	string	:=	"true";
		phase_steps_64_vs_128	:	string	:=	"phase_steps_64";
		phase_steps_sel	:	string	:=	"step40";
		power_mode	:	string	:=	"low_power";
		prot_mode	:	string	:=	"basic_rx";
		sel_oc_en	:	string	:=	"off_canc_disable";
		silicon_rev	:	string	:=	"20nm5es";
		step_ctrl_sel	:	string	:=	"feedback_mode";
		sup_mode	:	string	:=	"user_mode";
		v_vert_sel	:	string	:=	"plus";
		v_vert_threshold_scaling	:	string	:=	"scale_3";
		vert_threshold	:	string	:=	"vert_0"
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		clk0	:	in	std_logic	:=	'0';
		clk180	:	in	std_logic	:=	'0';
		clk270	:	in	std_logic	:=	'0';
		clk90	:	in	std_logic	:=	'0';
		it50u	:	in	std_logic	:=	'0';
		it50u2	:	in	std_logic	:=	'0';
		it50u4	:	in	std_logic	:=	'0';
		odi_atb_sel	:	in	std_logic_vector(2 downto 0)	:=	"000";
		odi_dft_clr	:	in	std_logic	:=	'0';
		odi_latch_clk	:	in	std_logic	:=	'0';
		odi_shift_clk	:	in	std_logic	:=	'0';
		odi_shift_in	:	in	std_logic	:=	'0';
		rx_n	:	in	std_logic	:=	'0';
		rx_p	:	in	std_logic	:=	'0';
		rxn_sum	:	in	std_logic	:=	'0';
		rxp_sum	:	in	std_logic	:=	'0';
		spec_vrefh	:	in	std_logic	:=	'0';
		spec_vrefl	:	in	std_logic	:=	'0';
		vcm_vref	:	in	std_logic	:=	'0';
		vertical_fb	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		atb0	:	out	std_logic	:=	'0';
		atb1	:	out	std_logic	:=	'0';
		clk0_eye	:	out	std_logic	:=	'0';
		clk0_eye_lb	:	out	std_logic	:=	'0';
		clk180_eye	:	out	std_logic	:=	'0';
		clk180_eye_lb	:	out	std_logic	:=	'0';
		de_eye	:	out	std_logic	:=	'0';
		deb_eye	:	out	std_logic	:=	'0';
		do_eye	:	out	std_logic	:=	'0';
		dob_eye	:	out	std_logic	:=	'0';
		odi_en	:	out	std_logic	:=	'0';
		odi_oc_tstmx	:	out	std_logic_vector(1 downto 0)	:=	"00";
		tdr_en	:	out	std_logic	:=	'0';
		vref_sel_out	:	out	std_logic	:=	'0'
	);
end component;

begin



inst : twentynm_hssi_pma_rx_odi_encrypted
	generic map (
		-- Instance parameters
		clk_dcd_bypass	=>	clk_dcd_bypass,
		datarate	=>	datarate,
		enable_odi	=>	enable_odi,
		initial_settings	=>	initial_settings,
		invert_dfe_vref	=>	invert_dfe_vref,
		monitor_bw_sel	=>	monitor_bw_sel,
		oc_sa_c0	=>	oc_sa_c0_int,
		oc_sa_c180	=>	oc_sa_c180_int,
		optimal	=>	optimal,
		phase_steps_64_vs_128	=>	phase_steps_64_vs_128,
		phase_steps_sel	=>	phase_steps_sel,
		power_mode	=>	power_mode,
		prot_mode	=>	prot_mode,
		sel_oc_en	=>	sel_oc_en,
		silicon_rev	=>	silicon_rev,
		step_ctrl_sel	=>	step_ctrl_sel,
		sup_mode	=>	sup_mode,
		v_vert_sel	=>	v_vert_sel,
		v_vert_threshold_scaling	=>	v_vert_threshold_scaling,
		vert_threshold	=>	vert_threshold
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		clk0	=>	clk0,
		clk180	=>	clk180,
		clk270	=>	clk270,
		clk90	=>	clk90,
		it50u	=>	it50u,
		it50u2	=>	it50u2,
		it50u4	=>	it50u4,
		odi_atb_sel	=>	odi_atb_sel,
		odi_dft_clr	=>	odi_dft_clr,
		odi_latch_clk	=>	odi_latch_clk,
		odi_shift_clk	=>	odi_shift_clk,
		odi_shift_in	=>	odi_shift_in,
		rx_n	=>	rx_n,
		rx_p	=>	rx_p,
		rxn_sum	=>	rxn_sum,
		rxp_sum	=>	rxp_sum,
		spec_vrefh	=>	spec_vrefh,
		spec_vrefl	=>	spec_vrefl,
		vcm_vref	=>	vcm_vref,
		vertical_fb	=>	vertical_fb,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		atb0	=>	atb0,
		atb1	=>	atb1,
		clk0_eye	=>	clk0_eye,
		clk0_eye_lb	=>	clk0_eye_lb,
		clk180_eye	=>	clk180_eye,
		clk180_eye_lb	=>	clk180_eye_lb,
		de_eye	=>	de_eye,
		deb_eye	=>	deb_eye,
		do_eye	=>	do_eye,
		dob_eye	=>	dob_eye,
		odi_en	=>	odi_en,
		odi_oc_tstmx	=>	odi_oc_tstmx,
		tdr_en	=>	tdr_en,
		vref_sel_out	=>	vref_sel_out
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_pma_rx_sd	is
	generic (
		-- Entity parameters
		link	:	string	:=	"sr";
		optimal	:	string	:=	"true";
		power_mode	:	string	:=	"low_power";
		prot_mode	:	string	:=	"basic_rx";
		sd_output_off	:	integer	:=	1;
		sd_output_on	:	integer	:=	1;
		sd_pdb	:	string	:=	"sd_off";
		sd_threshold	:	string	:=	"sdlv_3";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		clk	:	in	std_logic	:=	'0';
		qpi	:	in	std_logic	:=	'0';
		rstn_sd	:	in	std_logic	:=	'0';
		s_lpbk_b	:	in	std_logic	:=	'0';
		vin	:	in	std_logic	:=	'0';
		vip	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		sd	:	out	std_logic	:=	'0'
	);
end twentynm_hssi_pma_rx_sd;

architecture behavior of twentynm_hssi_pma_rx_sd	is




component	twentynm_hssi_pma_rx_sd_encrypted
	generic (
		-- Architecture parameters
		link	:	string	:=	"sr";
		optimal	:	string	:=	"true";
		power_mode	:	string	:=	"low_power";
		prot_mode	:	string	:=	"basic_rx";
		sd_output_off	:	integer	:=	1;
		sd_output_on	:	integer	:=	1;
		sd_pdb	:	string	:=	"sd_off";
		sd_threshold	:	string	:=	"sdlv_3";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode"
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		clk	:	in	std_logic	:=	'0';
		qpi	:	in	std_logic	:=	'0';
		rstn_sd	:	in	std_logic	:=	'0';
		s_lpbk_b	:	in	std_logic	:=	'0';
		vin	:	in	std_logic	:=	'0';
		vip	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		sd	:	out	std_logic	:=	'0'
	);
end component;

begin



inst : twentynm_hssi_pma_rx_sd_encrypted
	generic map (
		-- Instance parameters
		link	=>	link,
		optimal	=>	optimal,
		power_mode	=>	power_mode,
		prot_mode	=>	prot_mode,
		sd_output_off	=>	sd_output_off,
		sd_output_on	=>	sd_output_on,
		sd_pdb	=>	sd_pdb,
		sd_threshold	=>	sd_threshold,
		silicon_rev	=>	silicon_rev,
		sup_mode	=>	sup_mode
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		clk	=>	clk,
		qpi	=>	qpi,
		rstn_sd	=>	rstn_sd,
		s_lpbk_b	=>	s_lpbk_b,
		vin	=>	vin,
		vip	=>	vip,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		sd	=>	sd
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_pma_tx_buf	is
	generic (
		-- Entity parameters
		calibration_en	:	string	:=	"false";
		calibration_resistor_value	:	string	:=	"res_setting0";
		cdr_cp_calibration_en	:	string	:=	"cdr_cp_cal_disable";
		chgpmp_current_dn_trim	:	string	:=	"cp_current_trimming_dn_setting0";
		chgpmp_current_up_trim	:	string	:=	"cp_current_trimming_up_setting0";
		chgpmp_dn_trim_double	:	string	:=	"normal_dn_trim_current";
		chgpmp_up_trim_double	:	string	:=	"normal_up_trim_current";
		compensation_driver_en	:	string	:=	"disable";
		compensation_en	:	string	:=	"enable";
		cpen_ctrl	:	string	:=	"cp_l0";
		datarate	:	string	:=	"0 bps";
		dcd_clk_div_ctrl	:	string	:=	"dcd_ck_div128";
		dcd_detection_en	:	string	:=	"enable";
		dft_sel	:	string	:=	"dft_disabled";
		duty_cycle_correction_bandwidth	:	string	:=	"dcc_bw_12";
		duty_cycle_correction_bandwidth_dn	:	string	:=	"dcd_bw_dn_0";
		duty_cycle_correction_mode_ctrl	:	string	:=	"dcc_disable";
		duty_cycle_correction_reference1	:	string	:=	"dcc_ref1_3";
		duty_cycle_correction_reference2	:	string	:=	"dcc_ref2_3";
		duty_cycle_correction_reset_n	:	string	:=	"reset_n";
		duty_cycle_cp_comp_en	:	string	:=	"cp_comp_off";
		duty_cycle_detector_cp_cal	:	string	:=	"dcd_cp_cal_disable";
		duty_cycle_detector_sa_cal	:	string	:=	"dcd_sa_cal_disable";
		duty_cycle_input_polarity	:	string	:=	"dcc_input_pos";
		duty_cycle_setting	:	string	:=	"dcc_t32";
		duty_cycle_setting_aux	:	string	:=	"dcc2_t32";
		enable_idle_tx_channel_support	:	string	:=	"false";
		initial_settings	:	string	:=	"false";
		jtag_drv_sel	:	string	:=	"drv1";
		jtag_lp	:	string	:=	"lp_off";
		link	:	string	:=	"sr";
		link_tx	:	string	:=	"sr";
		low_power_en	:	string	:=	"disable";
		lst	:	string	:=	"atb_disabled";
		mcgb_location_for_pcie	:	bit_vector	:=	B"0000";
		optimal	:	string	:=	"true";
		pm_speed_grade	:	string	:=	"e2";
		power_mode	:	string	:=	"low_power";
		power_rail_eht	:	integer	:=	0;
		power_rail_et	:	integer	:=	0;
		pre_emp_sign_1st_post_tap	:	string	:=	"fir_post_1t_neg";
		pre_emp_sign_2nd_post_tap	:	string	:=	"fir_post_2t_neg";
		pre_emp_sign_pre_tap_1t	:	string	:=	"fir_pre_1t_neg";
		pre_emp_sign_pre_tap_2t	:	string	:=	"fir_pre_2t_neg";
		pre_emp_switching_ctrl_1st_post_tap	:	bit_vector	:=	B"000000";
		pre_emp_switching_ctrl_2nd_post_tap	:	bit_vector	:=	B"0000";
		pre_emp_switching_ctrl_pre_tap_1t	:	bit_vector	:=	B"00000";
		pre_emp_switching_ctrl_pre_tap_2t	:	bit_vector	:=	B"000";
		prot_mode	:	string	:=	"basic_tx";
		res_cal_local	:	string	:=	"non_local";
		rx_det	:	string	:=	"mode_0";
		rx_det_output_sel	:	string	:=	"rx_det_pcie_out";
		rx_det_pdb	:	string	:=	"rx_det_off";
		sense_amp_offset_cal_curr_n	:	string	:=	"sa_os_cal_in_0";
		sense_amp_offset_cal_curr_p	:	bit_vector	:=	B"00000";
		ser_powerdown	:	string	:=	"power_down_ser";
		silicon_rev	:	string	:=	"20nm5es";
		slew_rate_ctrl	:	string	:=	"slew_r7";
		sup_mode	:	string	:=	"user_mode";
		swing_level	:	string	:=	"lv";
		term_code	:	string	:=	"rterm_code7";
		term_n_tune	:	string	:=	"rterm_n0";
		term_p_tune	:	string	:=	"rterm_p0";
		term_sel	:	string	:=	"r_r1";
		tri_driver	:	string	:=	"tri_driver_disable";
		tx_powerdown	:	string	:=	"normal_tx_on";
		uc_dcd_cal	:	string	:=	"uc_dcd_cal_off";
		uc_dcd_cal_status	:	string	:=	"uc_dcd_cal_notdone";
		uc_gen3	:	string	:=	"gen3_off";
		uc_gen4	:	string	:=	"gen4_off";
		uc_skew_cal	:	string	:=	"uc_skew_cal_off";
		uc_skew_cal_status	:	string	:=	"uc_skew_cal_notdone";
		uc_txvod_cal	:	string	:=	"uc_tx_vod_cal_off";
		uc_txvod_cal_cont	:	string	:=	"uc_tx_vod_cal_cont_off";
		uc_txvod_cal_status	:	string	:=	"uc_tx_vod_cal_notdone";
		uc_vcc_setting	:	string	:=	"vcc_setting0";
		user_fir_coeff_ctrl_sel	:	string	:=	"ram_ctl";
		vod_output_swing_ctrl	:	bit_vector	:=	B"00000";
		vreg_output	:	string	:=	"vccdreg_nominal";
		xtx_path_analog_mode	:	string	:=	"user_custom";
		xtx_path_bonding_mode	:	string	:=	"x1_non_bonded";
		xtx_path_calibration_en	:	string	:=	"false";
		xtx_path_clock_divider_ratio	:	bit_vector	:=	B"0000";
		xtx_path_datarate	:	string	:=	"0 bps";
		xtx_path_datawidth	:	bit_vector	:=	B"00000000";
		xtx_path_gt_enabled	:	string	:=	"disable";
		xtx_path_initial_settings	:	string	:=	"false";
		xtx_path_optimal	:	string	:=	"true";
		xtx_path_pma_tx_divclk_hz	:	string	:=	"00000000000000000000000000000000";
		xtx_path_prot_mode	:	string	:=	"basic_tx";
		xtx_path_sup_mode	:	string	:=	"user_mode";
		xtx_path_swing_level	:	string	:=	"lv";
		xtx_path_tx_pll_clk_hz	:	string	:=	"0 hz"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		bsmode	:	in	std_logic	:=	'0';
		bsoeb	:	in	std_logic	:=	'0';
		bstxn_in	:	in	std_logic	:=	'0';
		bstxp_in	:	in	std_logic	:=	'0';
		clk0_tx	:	in	std_logic	:=	'0';
		clk180_tx	:	in	std_logic	:=	'0';
		clk_dcd	:	in	std_logic	:=	'0';
		clksn	:	in	std_logic	:=	'0';
		clksp	:	in	std_logic	:=	'0';
		cr_rdynamic_sw	:	in	std_logic	:=	'0';
		i_coeff	:	in	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		oe	:	in	std_logic	:=	'0';
		oeb	:	in	std_logic	:=	'0';
		oo	:	in	std_logic	:=	'0';
		oob	:	in	std_logic	:=	'0';
		pcie_sw_master	:	in	std_logic	:=	'0';
		rx_det_clk	:	in	std_logic	:=	'0';
		rx_n_bidir_in	:	in	std_logic	:=	'0';
		rx_p_bidir_in	:	in	std_logic	:=	'0';
		s_lpbk_b	:	in	std_logic	:=	'0';
		tx50	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		tx_det_rx	:	in	std_logic	:=	'0';
		tx_elec_idle	:	in	std_logic	:=	'0';
		tx_qpi_pulldn	:	in	std_logic	:=	'0';
		tx_qpi_pullup	:	in	std_logic	:=	'0';
		tx_rlpbk	:	in	std_logic	:=	'0';
		vrlpbkn	:	in	std_logic	:=	'0';
		vrlpbkn_1t	:	in	std_logic	:=	'0';
		vrlpbkp	:	in	std_logic	:=	'0';
		vrlpbkp_1t	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		atbsel	:	out	std_logic_vector(2 downto 0)	:=	"000";
		ckn	:	out	std_logic	:=	'0';
		ckp	:	out	std_logic	:=	'0';
		dcd_out1	:	out	std_logic	:=	'0';
		dcd_out2	:	out	std_logic	:=	'0';
		dcd_out_ready	:	out	std_logic	:=	'0';
		detect_on	:	out	std_logic_vector(1 downto 0)	:=	"00";
		lbvon	:	out	std_logic	:=	'0';
		lbvop	:	out	std_logic	:=	'0';
		rx_detect_valid	:	out	std_logic	:=	'0';
		rx_found	:	out	std_logic	:=	'0';
		rx_found_pcie_spl_test	:	out	std_logic	:=	'0';
		sel_vreg	:	out	std_logic	:=	'0';
		spl_clk_test	:	out	std_logic	:=	'0';
		tx_dftout	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		vlptxn	:	out	std_logic	:=	'0';
		vlptxp	:	out	std_logic	:=	'0';
		von	:	out	std_logic	:=	'0';
		vop	:	out	std_logic	:=	'0'
	);
end twentynm_hssi_pma_tx_buf;

architecture behavior of twentynm_hssi_pma_tx_buf	is

constant mcgb_location_for_pcie_int	:	integer	:=	bin2int(mcgb_location_for_pcie);
constant pre_emp_switching_ctrl_1st_post_tap_int	:	integer	:=	bin2int(pre_emp_switching_ctrl_1st_post_tap);
constant pre_emp_switching_ctrl_2nd_post_tap_int	:	integer	:=	bin2int(pre_emp_switching_ctrl_2nd_post_tap);
constant pre_emp_switching_ctrl_pre_tap_1t_int	:	integer	:=	bin2int(pre_emp_switching_ctrl_pre_tap_1t);
constant pre_emp_switching_ctrl_pre_tap_2t_int	:	integer	:=	bin2int(pre_emp_switching_ctrl_pre_tap_2t);
constant sense_amp_offset_cal_curr_p_int	:	integer	:=	bin2int(sense_amp_offset_cal_curr_p);
constant vod_output_swing_ctrl_int	:	integer	:=	bin2int(vod_output_swing_ctrl);
constant xtx_path_clock_divider_ratio_int	:	integer	:=	bin2int(xtx_path_clock_divider_ratio);
constant xtx_path_datawidth_int	:	integer	:=	bin2int(xtx_path_datawidth);



component	twentynm_hssi_pma_tx_buf_encrypted
	generic (
		-- Architecture parameters
		calibration_en	:	string	:=	"false";
		calibration_resistor_value	:	string	:=	"res_setting0";
		cdr_cp_calibration_en	:	string	:=	"cdr_cp_cal_disable";
		chgpmp_current_dn_trim	:	string	:=	"cp_current_trimming_dn_setting0";
		chgpmp_current_up_trim	:	string	:=	"cp_current_trimming_up_setting0";
		chgpmp_dn_trim_double	:	string	:=	"normal_dn_trim_current";
		chgpmp_up_trim_double	:	string	:=	"normal_up_trim_current";
		compensation_driver_en	:	string	:=	"disable";
		compensation_en	:	string	:=	"enable";
		cpen_ctrl	:	string	:=	"cp_l0";
		datarate	:	string	:=	"0 bps";
		dcd_clk_div_ctrl	:	string	:=	"dcd_ck_div128";
		dcd_detection_en	:	string	:=	"enable";
		dft_sel	:	string	:=	"dft_disabled";
		duty_cycle_correction_bandwidth	:	string	:=	"dcc_bw_12";
		duty_cycle_correction_bandwidth_dn	:	string	:=	"dcd_bw_dn_0";
		duty_cycle_correction_mode_ctrl	:	string	:=	"dcc_disable";
		duty_cycle_correction_reference1	:	string	:=	"dcc_ref1_3";
		duty_cycle_correction_reference2	:	string	:=	"dcc_ref2_3";
		duty_cycle_correction_reset_n	:	string	:=	"reset_n";
		duty_cycle_cp_comp_en	:	string	:=	"cp_comp_off";
		duty_cycle_detector_cp_cal	:	string	:=	"dcd_cp_cal_disable";
		duty_cycle_detector_sa_cal	:	string	:=	"dcd_sa_cal_disable";
		duty_cycle_input_polarity	:	string	:=	"dcc_input_pos";
		duty_cycle_setting	:	string	:=	"dcc_t32";
		duty_cycle_setting_aux	:	string	:=	"dcc2_t32";
		enable_idle_tx_channel_support	:	string	:=	"false";
		initial_settings	:	string	:=	"false";
		jtag_drv_sel	:	string	:=	"drv1";
		jtag_lp	:	string	:=	"lp_off";
		link	:	string	:=	"sr";
		link_tx	:	string	:=	"sr";
		low_power_en	:	string	:=	"disable";
		lst	:	string	:=	"atb_disabled";
		mcgb_location_for_pcie	:	integer	:=	0;
		optimal	:	string	:=	"true";
		pm_speed_grade	:	string	:=	"e2";
		power_mode	:	string	:=	"low_power";
		power_rail_eht	:	integer	:=	0;
		power_rail_et	:	integer	:=	0;
		pre_emp_sign_1st_post_tap	:	string	:=	"fir_post_1t_neg";
		pre_emp_sign_2nd_post_tap	:	string	:=	"fir_post_2t_neg";
		pre_emp_sign_pre_tap_1t	:	string	:=	"fir_pre_1t_neg";
		pre_emp_sign_pre_tap_2t	:	string	:=	"fir_pre_2t_neg";
		pre_emp_switching_ctrl_1st_post_tap	:	integer	:=	0;
		pre_emp_switching_ctrl_2nd_post_tap	:	integer	:=	0;
		pre_emp_switching_ctrl_pre_tap_1t	:	integer	:=	0;
		pre_emp_switching_ctrl_pre_tap_2t	:	integer	:=	0;
		prot_mode	:	string	:=	"basic_tx";
		res_cal_local	:	string	:=	"non_local";
		rx_det	:	string	:=	"mode_0";
		rx_det_output_sel	:	string	:=	"rx_det_pcie_out";
		rx_det_pdb	:	string	:=	"rx_det_off";
		sense_amp_offset_cal_curr_n	:	string	:=	"sa_os_cal_in_0";
		sense_amp_offset_cal_curr_p	:	integer	:=	0;
		ser_powerdown	:	string	:=	"power_down_ser";
		silicon_rev	:	string	:=	"20nm5es";
		slew_rate_ctrl	:	string	:=	"slew_r7";
		sup_mode	:	string	:=	"user_mode";
		swing_level	:	string	:=	"lv";
		term_code	:	string	:=	"rterm_code7";
		term_n_tune	:	string	:=	"rterm_n0";
		term_p_tune	:	string	:=	"rterm_p0";
		term_sel	:	string	:=	"r_r1";
		tri_driver	:	string	:=	"tri_driver_disable";
		tx_powerdown	:	string	:=	"normal_tx_on";
		uc_dcd_cal	:	string	:=	"uc_dcd_cal_off";
		uc_dcd_cal_status	:	string	:=	"uc_dcd_cal_notdone";
		uc_gen3	:	string	:=	"gen3_off";
		uc_gen4	:	string	:=	"gen4_off";
		uc_skew_cal	:	string	:=	"uc_skew_cal_off";
		uc_skew_cal_status	:	string	:=	"uc_skew_cal_notdone";
		uc_txvod_cal	:	string	:=	"uc_tx_vod_cal_off";
		uc_txvod_cal_cont	:	string	:=	"uc_tx_vod_cal_cont_off";
		uc_txvod_cal_status	:	string	:=	"uc_tx_vod_cal_notdone";
		uc_vcc_setting	:	string	:=	"vcc_setting0";
		user_fir_coeff_ctrl_sel	:	string	:=	"ram_ctl";
		vod_output_swing_ctrl	:	integer	:=	0;
		vreg_output	:	string	:=	"vccdreg_nominal";
		xtx_path_analog_mode	:	string	:=	"user_custom";
		xtx_path_bonding_mode	:	string	:=	"x1_non_bonded";
		xtx_path_calibration_en	:	string	:=	"false";
		xtx_path_clock_divider_ratio	:	integer	:=	0;
		xtx_path_datarate	:	string	:=	"0 bps";
		xtx_path_datawidth	:	integer	:=	0;
		xtx_path_gt_enabled	:	string	:=	"disable";
		xtx_path_initial_settings	:	string	:=	"false";
		xtx_path_optimal	:	string	:=	"true";
		xtx_path_pma_tx_divclk_hz	:	string	:=	"00000000000000000000000000000000";
		xtx_path_prot_mode	:	string	:=	"basic_tx";
		xtx_path_sup_mode	:	string	:=	"user_mode";
		xtx_path_swing_level	:	string	:=	"lv";
		xtx_path_tx_pll_clk_hz	:	string	:=	"0 hz"
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		bsmode	:	in	std_logic	:=	'0';
		bsoeb	:	in	std_logic	:=	'0';
		bstxn_in	:	in	std_logic	:=	'0';
		bstxp_in	:	in	std_logic	:=	'0';
		clk0_tx	:	in	std_logic	:=	'0';
		clk180_tx	:	in	std_logic	:=	'0';
		clk_dcd	:	in	std_logic	:=	'0';
		clksn	:	in	std_logic	:=	'0';
		clksp	:	in	std_logic	:=	'0';
		cr_rdynamic_sw	:	in	std_logic	:=	'0';
		i_coeff	:	in	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		oe	:	in	std_logic	:=	'0';
		oeb	:	in	std_logic	:=	'0';
		oo	:	in	std_logic	:=	'0';
		oob	:	in	std_logic	:=	'0';
		pcie_sw_master	:	in	std_logic	:=	'0';
		rx_det_clk	:	in	std_logic	:=	'0';
		rx_n_bidir_in	:	in	std_logic	:=	'0';
		rx_p_bidir_in	:	in	std_logic	:=	'0';
		s_lpbk_b	:	in	std_logic	:=	'0';
		tx50	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		tx_det_rx	:	in	std_logic	:=	'0';
		tx_elec_idle	:	in	std_logic	:=	'0';
		tx_qpi_pulldn	:	in	std_logic	:=	'0';
		tx_qpi_pullup	:	in	std_logic	:=	'0';
		tx_rlpbk	:	in	std_logic	:=	'0';
		vrlpbkn	:	in	std_logic	:=	'0';
		vrlpbkn_1t	:	in	std_logic	:=	'0';
		vrlpbkp	:	in	std_logic	:=	'0';
		vrlpbkp_1t	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		atbsel	:	out	std_logic_vector(2 downto 0)	:=	"000";
		ckn	:	out	std_logic	:=	'0';
		ckp	:	out	std_logic	:=	'0';
		dcd_out1	:	out	std_logic	:=	'0';
		dcd_out2	:	out	std_logic	:=	'0';
		dcd_out_ready	:	out	std_logic	:=	'0';
		detect_on	:	out	std_logic_vector(1 downto 0)	:=	"00";
		lbvon	:	out	std_logic	:=	'0';
		lbvop	:	out	std_logic	:=	'0';
		rx_detect_valid	:	out	std_logic	:=	'0';
		rx_found	:	out	std_logic	:=	'0';
		rx_found_pcie_spl_test	:	out	std_logic	:=	'0';
		sel_vreg	:	out	std_logic	:=	'0';
		spl_clk_test	:	out	std_logic	:=	'0';
		tx_dftout	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		vlptxn	:	out	std_logic	:=	'0';
		vlptxp	:	out	std_logic	:=	'0';
		von	:	out	std_logic	:=	'0';
		vop	:	out	std_logic	:=	'0'
	);
end component;

begin



inst : twentynm_hssi_pma_tx_buf_encrypted
	generic map (
		-- Instance parameters
		calibration_en	=>	calibration_en,
		calibration_resistor_value	=>	calibration_resistor_value,
		cdr_cp_calibration_en	=>	cdr_cp_calibration_en,
		chgpmp_current_dn_trim	=>	chgpmp_current_dn_trim,
		chgpmp_current_up_trim	=>	chgpmp_current_up_trim,
		chgpmp_dn_trim_double	=>	chgpmp_dn_trim_double,
		chgpmp_up_trim_double	=>	chgpmp_up_trim_double,
		compensation_driver_en	=>	compensation_driver_en,
		compensation_en	=>	compensation_en,
		cpen_ctrl	=>	cpen_ctrl,
		datarate	=>	datarate,
		dcd_clk_div_ctrl	=>	dcd_clk_div_ctrl,
		dcd_detection_en	=>	dcd_detection_en,
		dft_sel	=>	dft_sel,
		duty_cycle_correction_bandwidth	=>	duty_cycle_correction_bandwidth,
		duty_cycle_correction_bandwidth_dn	=>	duty_cycle_correction_bandwidth_dn,
		duty_cycle_correction_mode_ctrl	=>	duty_cycle_correction_mode_ctrl,
		duty_cycle_correction_reference1	=>	duty_cycle_correction_reference1,
		duty_cycle_correction_reference2	=>	duty_cycle_correction_reference2,
		duty_cycle_correction_reset_n	=>	duty_cycle_correction_reset_n,
		duty_cycle_cp_comp_en	=>	duty_cycle_cp_comp_en,
		duty_cycle_detector_cp_cal	=>	duty_cycle_detector_cp_cal,
		duty_cycle_detector_sa_cal	=>	duty_cycle_detector_sa_cal,
		duty_cycle_input_polarity	=>	duty_cycle_input_polarity,
		duty_cycle_setting	=>	duty_cycle_setting,
		duty_cycle_setting_aux	=>	duty_cycle_setting_aux,
		enable_idle_tx_channel_support	=>	enable_idle_tx_channel_support,
		initial_settings	=>	initial_settings,
		jtag_drv_sel	=>	jtag_drv_sel,
		jtag_lp	=>	jtag_lp,
		link	=>	link,
		link_tx	=>	link_tx,
		low_power_en	=>	low_power_en,
		lst	=>	lst,
		mcgb_location_for_pcie	=>	mcgb_location_for_pcie_int,
		optimal	=>	optimal,
		pm_speed_grade	=>	pm_speed_grade,
		power_mode	=>	power_mode,
		power_rail_eht	=>	power_rail_eht,
		power_rail_et	=>	power_rail_et,
		pre_emp_sign_1st_post_tap	=>	pre_emp_sign_1st_post_tap,
		pre_emp_sign_2nd_post_tap	=>	pre_emp_sign_2nd_post_tap,
		pre_emp_sign_pre_tap_1t	=>	pre_emp_sign_pre_tap_1t,
		pre_emp_sign_pre_tap_2t	=>	pre_emp_sign_pre_tap_2t,
		pre_emp_switching_ctrl_1st_post_tap	=>	pre_emp_switching_ctrl_1st_post_tap_int,
		pre_emp_switching_ctrl_2nd_post_tap	=>	pre_emp_switching_ctrl_2nd_post_tap_int,
		pre_emp_switching_ctrl_pre_tap_1t	=>	pre_emp_switching_ctrl_pre_tap_1t_int,
		pre_emp_switching_ctrl_pre_tap_2t	=>	pre_emp_switching_ctrl_pre_tap_2t_int,
		prot_mode	=>	prot_mode,
		res_cal_local	=>	res_cal_local,
		rx_det	=>	rx_det,
		rx_det_output_sel	=>	rx_det_output_sel,
		rx_det_pdb	=>	rx_det_pdb,
		sense_amp_offset_cal_curr_n	=>	sense_amp_offset_cal_curr_n,
		sense_amp_offset_cal_curr_p	=>	sense_amp_offset_cal_curr_p_int,
		ser_powerdown	=>	ser_powerdown,
		silicon_rev	=>	silicon_rev,
		slew_rate_ctrl	=>	slew_rate_ctrl,
		sup_mode	=>	sup_mode,
		swing_level	=>	swing_level,
		term_code	=>	term_code,
		term_n_tune	=>	term_n_tune,
		term_p_tune	=>	term_p_tune,
		term_sel	=>	term_sel,
		tri_driver	=>	tri_driver,
		tx_powerdown	=>	tx_powerdown,
		uc_dcd_cal	=>	uc_dcd_cal,
		uc_dcd_cal_status	=>	uc_dcd_cal_status,
		uc_gen3	=>	uc_gen3,
		uc_gen4	=>	uc_gen4,
		uc_skew_cal	=>	uc_skew_cal,
		uc_skew_cal_status	=>	uc_skew_cal_status,
		uc_txvod_cal	=>	uc_txvod_cal,
		uc_txvod_cal_cont	=>	uc_txvod_cal_cont,
		uc_txvod_cal_status	=>	uc_txvod_cal_status,
		uc_vcc_setting	=>	uc_vcc_setting,
		user_fir_coeff_ctrl_sel	=>	user_fir_coeff_ctrl_sel,
		vod_output_swing_ctrl	=>	vod_output_swing_ctrl_int,
		vreg_output	=>	vreg_output,
		xtx_path_analog_mode	=>	xtx_path_analog_mode,
		xtx_path_bonding_mode	=>	xtx_path_bonding_mode,
		xtx_path_calibration_en	=>	xtx_path_calibration_en,
		xtx_path_clock_divider_ratio	=>	xtx_path_clock_divider_ratio_int,
		xtx_path_datarate	=>	xtx_path_datarate,
		xtx_path_datawidth	=>	xtx_path_datawidth_int,
		xtx_path_gt_enabled	=>	xtx_path_gt_enabled,
		xtx_path_initial_settings	=>	xtx_path_initial_settings,
		xtx_path_optimal	=>	xtx_path_optimal,
		xtx_path_pma_tx_divclk_hz	=>	xtx_path_pma_tx_divclk_hz,
		xtx_path_prot_mode	=>	xtx_path_prot_mode,
		xtx_path_sup_mode	=>	xtx_path_sup_mode,
		xtx_path_swing_level	=>	xtx_path_swing_level,
		xtx_path_tx_pll_clk_hz	=>	xtx_path_tx_pll_clk_hz
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		bsmode	=>	bsmode,
		bsoeb	=>	bsoeb,
		bstxn_in	=>	bstxn_in,
		bstxp_in	=>	bstxp_in,
		clk0_tx	=>	clk0_tx,
		clk180_tx	=>	clk180_tx,
		clk_dcd	=>	clk_dcd,
		clksn	=>	clksn,
		clksp	=>	clksp,
		cr_rdynamic_sw	=>	cr_rdynamic_sw,
		i_coeff	=>	i_coeff,
		oe	=>	oe,
		oeb	=>	oeb,
		oo	=>	oo,
		oob	=>	oob,
		pcie_sw_master	=>	pcie_sw_master,
		rx_det_clk	=>	rx_det_clk,
		rx_n_bidir_in	=>	rx_n_bidir_in,
		rx_p_bidir_in	=>	rx_p_bidir_in,
		s_lpbk_b	=>	s_lpbk_b,
		tx50	=>	tx50,
		tx_det_rx	=>	tx_det_rx,
		tx_elec_idle	=>	tx_elec_idle,
		tx_qpi_pulldn	=>	tx_qpi_pulldn,
		tx_qpi_pullup	=>	tx_qpi_pullup,
		tx_rlpbk	=>	tx_rlpbk,
		vrlpbkn	=>	vrlpbkn,
		vrlpbkn_1t	=>	vrlpbkn_1t,
		vrlpbkp	=>	vrlpbkp,
		vrlpbkp_1t	=>	vrlpbkp_1t,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		atbsel	=>	atbsel,
		ckn	=>	ckn,
		ckp	=>	ckp,
		dcd_out1	=>	dcd_out1,
		dcd_out2	=>	dcd_out2,
		dcd_out_ready	=>	dcd_out_ready,
		detect_on	=>	detect_on,
		lbvon	=>	lbvon,
		lbvop	=>	lbvop,
		rx_detect_valid	=>	rx_detect_valid,
		rx_found	=>	rx_found,
		rx_found_pcie_spl_test	=>	rx_found_pcie_spl_test,
		sel_vreg	=>	sel_vreg,
		spl_clk_test	=>	spl_clk_test,
		tx_dftout	=>	tx_dftout,
		vlptxn	=>	vlptxn,
		vlptxp	=>	vlptxp,
		von	=>	von,
		vop	=>	vop
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_pma_tx_cgb	is
	generic (
		-- Entity parameters
		bitslip_enable	:	string	:=	"enable_bitslip";
		bonding_mode	:	string	:=	"x1_non_bonded";
		bonding_reset_enable	:	string	:=	"allow_bonding_reset";
		cgb_power_down	:	string	:=	"power_down_cgb";
		datarate	:	string	:=	"0 bps";
		dprio_cgb_vreg_boost	:	string	:=	"no_voltage_boost";
		initial_settings	:	string	:=	"false";
		input_select_gen3	:	string	:=	"unused";
		input_select_x1	:	string	:=	"unused";
		input_select_xn	:	string	:=	"unused";
		observe_cgb_clocks	:	string	:=	"observe_nothing";
		pcie_gen3_bitwidth	:	string	:=	"pciegen3_wide";
		prot_mode	:	string	:=	"basic_tx";
		scratch0_x1_clock_src	:	string	:=	"unused";
		scratch1_x1_clock_src	:	string	:=	"unused";
		scratch2_x1_clock_src	:	string	:=	"unused";
		scratch3_x1_clock_src	:	string	:=	"unused";
		select_done_master_or_slave	:	string	:=	"choose_slave_pcie_sw_done";
		ser_mode	:	string	:=	"eight_bit";
		ser_powerdown	:	string	:=	"normal_poweron_ser";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode";
		tx_ucontrol_en	:	string	:=	"disable";
		tx_ucontrol_pcie	:	string	:=	"gen1";
		tx_ucontrol_reset	:	string	:=	"disable";
		vccdreg_output	:	string	:=	"vccdreg_nominal";
		x1_clock_source_sel	:	string	:=	"cdr_txpll_t";
		x1_div_m_sel	:	string	:=	"divbypass";
		xn_clock_source_sel	:	string	:=	"sel_xn_up"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		ckdccn	:	in	std_logic	:=	'0';
		ckdccp	:	in	std_logic	:=	'0';
		clk_cdr_b	:	in	std_logic	:=	'0';
		clk_cdr_direct	:	in	std_logic	:=	'0';
		clk_cdr_t	:	in	std_logic	:=	'0';
		clk_fpll_b	:	in	std_logic	:=	'0';
		clk_fpll_t	:	in	std_logic	:=	'0';
		clk_lc_b	:	in	std_logic	:=	'0';
		clk_lc_hs	:	in	std_logic	:=	'0';
		clk_lc_t	:	in	std_logic	:=	'0';
		clkb_cdr_b	:	in	std_logic	:=	'0';
		clkb_cdr_direct	:	in	std_logic	:=	'0';
		clkb_cdr_t	:	in	std_logic	:=	'0';
		clkb_fpll_b	:	in	std_logic	:=	'0';
		clkb_fpll_t	:	in	std_logic	:=	'0';
		clkb_lc_b	:	in	std_logic	:=	'0';
		clkb_lc_hs	:	in	std_logic	:=	'0';
		clkb_lc_t	:	in	std_logic	:=	'0';
		cpulse_x6_dn_bus	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		cpulse_x6_up_bus	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		cpulse_xn_dn_bus	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		cpulse_xn_up_bus	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		pcie_sw	:	in	std_logic_vector(1 downto 0)	:=	"00";
		pcie_sw_done_master	:	in	std_logic_vector(1 downto 0)	:=	"00";
		tx_bitslip	:	in	std_logic	:=	'0';
		tx_bonding_rstb	:	in	std_logic	:=	'0';
		tx_pma_rstb	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		bitslipstate	:	out	std_logic	:=	'0';
		cpulse_out_bus	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		div2	:	out	std_logic	:=	'0';
		div4	:	out	std_logic	:=	'0';
		div5	:	out	std_logic	:=	'0';
		hifreqclkn	:	out	std_logic	:=	'0';
		hifreqclkp	:	out	std_logic	:=	'0';
		pcie_sw_done	:	out	std_logic_vector(1 downto 0)	:=	"00";
		pcie_sw_master	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rstb	:	out	std_logic	:=	'0'
	);
end twentynm_hssi_pma_tx_cgb;

architecture behavior of twentynm_hssi_pma_tx_cgb	is




component	twentynm_hssi_pma_tx_cgb_encrypted
	generic (
		-- Architecture parameters
		bitslip_enable	:	string	:=	"enable_bitslip";
		bonding_mode	:	string	:=	"x1_non_bonded";
		bonding_reset_enable	:	string	:=	"allow_bonding_reset";
		cgb_power_down	:	string	:=	"power_down_cgb";
		datarate	:	string	:=	"0 bps";
		dprio_cgb_vreg_boost	:	string	:=	"no_voltage_boost";
		initial_settings	:	string	:=	"false";
		input_select_gen3	:	string	:=	"unused";
		input_select_x1	:	string	:=	"unused";
		input_select_xn	:	string	:=	"unused";
		observe_cgb_clocks	:	string	:=	"observe_nothing";
		pcie_gen3_bitwidth	:	string	:=	"pciegen3_wide";
		prot_mode	:	string	:=	"basic_tx";
		scratch0_x1_clock_src	:	string	:=	"unused";
		scratch1_x1_clock_src	:	string	:=	"unused";
		scratch2_x1_clock_src	:	string	:=	"unused";
		scratch3_x1_clock_src	:	string	:=	"unused";
		select_done_master_or_slave	:	string	:=	"choose_slave_pcie_sw_done";
		ser_mode	:	string	:=	"eight_bit";
		ser_powerdown	:	string	:=	"normal_poweron_ser";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode";
		tx_ucontrol_en	:	string	:=	"disable";
		tx_ucontrol_pcie	:	string	:=	"gen1";
		tx_ucontrol_reset	:	string	:=	"disable";
		vccdreg_output	:	string	:=	"vccdreg_nominal";
		x1_clock_source_sel	:	string	:=	"cdr_txpll_t";
		x1_div_m_sel	:	string	:=	"divbypass";
		xn_clock_source_sel	:	string	:=	"sel_xn_up"
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		ckdccn	:	in	std_logic	:=	'0';
		ckdccp	:	in	std_logic	:=	'0';
		clk_cdr_b	:	in	std_logic	:=	'0';
		clk_cdr_direct	:	in	std_logic	:=	'0';
		clk_cdr_t	:	in	std_logic	:=	'0';
		clk_fpll_b	:	in	std_logic	:=	'0';
		clk_fpll_t	:	in	std_logic	:=	'0';
		clk_lc_b	:	in	std_logic	:=	'0';
		clk_lc_hs	:	in	std_logic	:=	'0';
		clk_lc_t	:	in	std_logic	:=	'0';
		clkb_cdr_b	:	in	std_logic	:=	'0';
		clkb_cdr_direct	:	in	std_logic	:=	'0';
		clkb_cdr_t	:	in	std_logic	:=	'0';
		clkb_fpll_b	:	in	std_logic	:=	'0';
		clkb_fpll_t	:	in	std_logic	:=	'0';
		clkb_lc_b	:	in	std_logic	:=	'0';
		clkb_lc_hs	:	in	std_logic	:=	'0';
		clkb_lc_t	:	in	std_logic	:=	'0';
		cpulse_x6_dn_bus	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		cpulse_x6_up_bus	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		cpulse_xn_dn_bus	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		cpulse_xn_up_bus	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		pcie_sw	:	in	std_logic_vector(1 downto 0)	:=	"00";
		pcie_sw_done_master	:	in	std_logic_vector(1 downto 0)	:=	"00";
		tx_bitslip	:	in	std_logic	:=	'0';
		tx_bonding_rstb	:	in	std_logic	:=	'0';
		tx_pma_rstb	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		bitslipstate	:	out	std_logic	:=	'0';
		cpulse_out_bus	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		div2	:	out	std_logic	:=	'0';
		div4	:	out	std_logic	:=	'0';
		div5	:	out	std_logic	:=	'0';
		hifreqclkn	:	out	std_logic	:=	'0';
		hifreqclkp	:	out	std_logic	:=	'0';
		pcie_sw_done	:	out	std_logic_vector(1 downto 0)	:=	"00";
		pcie_sw_master	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rstb	:	out	std_logic	:=	'0'
	);
end component;

begin



inst : twentynm_hssi_pma_tx_cgb_encrypted
	generic map (
		-- Instance parameters
		bitslip_enable	=>	bitslip_enable,
		bonding_mode	=>	bonding_mode,
		bonding_reset_enable	=>	bonding_reset_enable,
		cgb_power_down	=>	cgb_power_down,
		datarate	=>	datarate,
		dprio_cgb_vreg_boost	=>	dprio_cgb_vreg_boost,
		initial_settings	=>	initial_settings,
		input_select_gen3	=>	input_select_gen3,
		input_select_x1	=>	input_select_x1,
		input_select_xn	=>	input_select_xn,
		observe_cgb_clocks	=>	observe_cgb_clocks,
		pcie_gen3_bitwidth	=>	pcie_gen3_bitwidth,
		prot_mode	=>	prot_mode,
		scratch0_x1_clock_src	=>	scratch0_x1_clock_src,
		scratch1_x1_clock_src	=>	scratch1_x1_clock_src,
		scratch2_x1_clock_src	=>	scratch2_x1_clock_src,
		scratch3_x1_clock_src	=>	scratch3_x1_clock_src,
		select_done_master_or_slave	=>	select_done_master_or_slave,
		ser_mode	=>	ser_mode,
		ser_powerdown	=>	ser_powerdown,
		silicon_rev	=>	silicon_rev,
		sup_mode	=>	sup_mode,
		tx_ucontrol_en	=>	tx_ucontrol_en,
		tx_ucontrol_pcie	=>	tx_ucontrol_pcie,
		tx_ucontrol_reset	=>	tx_ucontrol_reset,
		vccdreg_output	=>	vccdreg_output,
		x1_clock_source_sel	=>	x1_clock_source_sel,
		x1_div_m_sel	=>	x1_div_m_sel,
		xn_clock_source_sel	=>	xn_clock_source_sel
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		ckdccn	=>	ckdccn,
		ckdccp	=>	ckdccp,
		clk_cdr_b	=>	clk_cdr_b,
		clk_cdr_direct	=>	clk_cdr_direct,
		clk_cdr_t	=>	clk_cdr_t,
		clk_fpll_b	=>	clk_fpll_b,
		clk_fpll_t	=>	clk_fpll_t,
		clk_lc_b	=>	clk_lc_b,
		clk_lc_hs	=>	clk_lc_hs,
		clk_lc_t	=>	clk_lc_t,
		clkb_cdr_b	=>	clkb_cdr_b,
		clkb_cdr_direct	=>	clkb_cdr_direct,
		clkb_cdr_t	=>	clkb_cdr_t,
		clkb_fpll_b	=>	clkb_fpll_b,
		clkb_fpll_t	=>	clkb_fpll_t,
		clkb_lc_b	=>	clkb_lc_b,
		clkb_lc_hs	=>	clkb_lc_hs,
		clkb_lc_t	=>	clkb_lc_t,
		cpulse_x6_dn_bus	=>	cpulse_x6_dn_bus,
		cpulse_x6_up_bus	=>	cpulse_x6_up_bus,
		cpulse_xn_dn_bus	=>	cpulse_xn_dn_bus,
		cpulse_xn_up_bus	=>	cpulse_xn_up_bus,
		pcie_sw	=>	pcie_sw,
		pcie_sw_done_master	=>	pcie_sw_done_master,
		tx_bitslip	=>	tx_bitslip,
		tx_bonding_rstb	=>	tx_bonding_rstb,
		tx_pma_rstb	=>	tx_pma_rstb,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		bitslipstate	=>	bitslipstate,
		cpulse_out_bus	=>	cpulse_out_bus,
		div2	=>	div2,
		div4	=>	div4,
		div5	=>	div5,
		hifreqclkn	=>	hifreqclkn,
		hifreqclkp	=>	hifreqclkp,
		pcie_sw_done	=>	pcie_sw_done,
		pcie_sw_master	=>	pcie_sw_master,
		rstb	=>	rstb
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_pma_tx_ser	is
	generic (
		-- Entity parameters
		bonding_mode	:	string	:=	"x1_non_bonded";
		clk_divtx_deskew	:	string	:=	"deskew_delay8";
		control_clk_divtx	:	string	:=	"no_dft_control_clkdivtx";
		duty_cycle_correction_mode_ctrl	:	string	:=	"dcc_disable";
		initial_settings	:	string	:=	"false";
		prot_mode	:	string	:=	"basic_tx";
		ser_clk_divtx_user_sel	:	string	:=	"divtx_user_33";
		ser_clk_mon	:	string	:=	"disable_clk_mon";
		ser_powerdown	:	string	:=	"normal_poweron_ser";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		bitslipstate	:	in	std_logic	:=	'0';
		cpulse	:	in	std_logic	:=	'0';
		data	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		hfclkn	:	in	std_logic	:=	'0';
		hfclkp	:	in	std_logic	:=	'0';
		lfclk	:	in	std_logic	:=	'0';
		lfclk2	:	in	std_logic	:=	'0';
		paraclk	:	in	std_logic	:=	'0';
		rser_div2	:	in	std_logic	:=	'0';
		rser_div4	:	in	std_logic	:=	'0';
		rser_div5	:	in	std_logic	:=	'0';
		rst_n	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		ckdrvn	:	out	std_logic	:=	'0';
		ckdrvp	:	out	std_logic	:=	'0';
		clk_divtx	:	out	std_logic	:=	'0';
		clk_divtx_user	:	out	std_logic	:=	'0';
		oe	:	out	std_logic	:=	'0';
		oeb	:	out	std_logic	:=	'0';
		oo	:	out	std_logic	:=	'0';
		oob	:	out	std_logic	:=	'0'
	);
end twentynm_hssi_pma_tx_ser;

architecture behavior of twentynm_hssi_pma_tx_ser	is




component	twentynm_hssi_pma_tx_ser_encrypted
	generic (
		-- Architecture parameters
		bonding_mode	:	string	:=	"x1_non_bonded";
		clk_divtx_deskew	:	string	:=	"deskew_delay8";
		control_clk_divtx	:	string	:=	"no_dft_control_clkdivtx";
		duty_cycle_correction_mode_ctrl	:	string	:=	"dcc_disable";
		initial_settings	:	string	:=	"false";
		prot_mode	:	string	:=	"basic_tx";
		ser_clk_divtx_user_sel	:	string	:=	"divtx_user_33";
		ser_clk_mon	:	string	:=	"disable_clk_mon";
		ser_powerdown	:	string	:=	"normal_poweron_ser";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode"
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		bitslipstate	:	in	std_logic	:=	'0';
		cpulse	:	in	std_logic	:=	'0';
		data	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		hfclkn	:	in	std_logic	:=	'0';
		hfclkp	:	in	std_logic	:=	'0';
		lfclk	:	in	std_logic	:=	'0';
		lfclk2	:	in	std_logic	:=	'0';
		paraclk	:	in	std_logic	:=	'0';
		rser_div2	:	in	std_logic	:=	'0';
		rser_div4	:	in	std_logic	:=	'0';
		rser_div5	:	in	std_logic	:=	'0';
		rst_n	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		ckdrvn	:	out	std_logic	:=	'0';
		ckdrvp	:	out	std_logic	:=	'0';
		clk_divtx	:	out	std_logic	:=	'0';
		clk_divtx_user	:	out	std_logic	:=	'0';
		oe	:	out	std_logic	:=	'0';
		oeb	:	out	std_logic	:=	'0';
		oo	:	out	std_logic	:=	'0';
		oob	:	out	std_logic	:=	'0'
	);
end component;

begin



inst : twentynm_hssi_pma_tx_ser_encrypted
	generic map (
		-- Instance parameters
		bonding_mode	=>	bonding_mode,
		clk_divtx_deskew	=>	clk_divtx_deskew,
		control_clk_divtx	=>	control_clk_divtx,
		duty_cycle_correction_mode_ctrl	=>	duty_cycle_correction_mode_ctrl,
		initial_settings	=>	initial_settings,
		prot_mode	=>	prot_mode,
		ser_clk_divtx_user_sel	=>	ser_clk_divtx_user_sel,
		ser_clk_mon	=>	ser_clk_mon,
		ser_powerdown	=>	ser_powerdown,
		silicon_rev	=>	silicon_rev,
		sup_mode	=>	sup_mode
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		bitslipstate	=>	bitslipstate,
		cpulse	=>	cpulse,
		data	=>	data,
		hfclkn	=>	hfclkn,
		hfclkp	=>	hfclkp,
		lfclk	=>	lfclk,
		lfclk2	=>	lfclk2,
		paraclk	=>	paraclk,
		rser_div2	=>	rser_div2,
		rser_div4	=>	rser_div4,
		rser_div5	=>	rser_div5,
		rst_n	=>	rst_n,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		ckdrvn	=>	ckdrvn,
		ckdrvp	=>	ckdrvp,
		clk_divtx	=>	clk_divtx,
		clk_divtx_user	=>	clk_divtx_user,
		oe	=>	oe,
		oeb	=>	oeb,
		oo	=>	oo,
		oob	=>	oob
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_pma_uc	is
	generic (
		-- Entity parameters
		a_break_vector_word_addr	:	bit_vector	:=	B"0000000000001000";
		a_exception_vector_word_addr	:	bit_vector	:=	B"0000000000001000";
		a_reset_vector_word_addr	:	bit_vector	:=	B"0000000000000000";
		cal_mode	:	string	:=	"cal_en";
		pm_uc_aux_base_addr	:	bit_vector	:=	B"00000000";
		pm_uc_cal_clk_div	:	bit_vector	:=	B"00100";
		pm_uc_cal_clk_inv	:	string	:=	"disable_inv";
		pm_uc_cal_clk_ph	:	bit_vector	:=	B"00010";
		pm_uc_clkdiv_sel	:	string	:=	"div2";
		pm_uc_clksel_core	:	string	:=	"disable_core_clk";
		pm_uc_clksel_osc	:	string	:=	"cb_clkusr";
		pm_uc_core_jtg_rst_disable	:	string	:=	"disable_jtg_rst";
		pm_uc_core_sys_rst_disable	:	string	:=	"disable_core_rst";
		pm_uc_ecc_rst_disable	:	string	:=	"enable_ecc_rst";
		pm_uc_engg_opt	:	string	:=	"reserved";
		pm_uc_family_device_info	:	bit_vector	:=	B"000000000000000000000000";
		pm_uc_hssi_base_addr	:	bit_vector	:=	B"00000001";
		pm_uc_pcs_dft_out	:	bit_vector	:=	B"0000000000";
		pm_uc_pcs_dft_sel	:	string	:=	"disable_pcs_dft";
		pm_uc_pcs_rd_lat	:	bit_vector	:=	B"010";
		pm_uc_pcs_slave_count	:	bit_vector	:=	B"00000000";
		pm_uc_ram	:	string	:=	"00000000000000000000000000000000000000";
		pm_uc_rmw_dis	:	string	:=	"enable_rmw";
		pm_uc_soft_nios	:	string	:=	"disable_soft";
		pm_uc_sys_enable	:	string	:=	"enable_sys";
		pmu_cal_bin_fname	:	string	:=	"nf_hssi_cal_v10.hex'";
		pmu_qparam_fname	:	string	:=	"nf_qparam_nf1.hex'";
		powerdown_mode	:	string	:=	"powerdown";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode"
	);
	port (
		-- Entity ports
		cb_clkusr	:	in	std_logic	:=	'0';
		cb_intosc	:	in	std_logic	:=	'0';
		core_avl_clk	:	in	std_logic	:=	'0';
		core_avl_readdata	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		core_avl_readdatavalid	:	in	std_logic	:=	'0';
		core_avl_rst_n	:	in	std_logic	:=	'0';
		core_avl_waitrequest	:	in	std_logic	:=	'0';
		core_interrupt_in	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		core_uc_rst_n	:	in	std_logic	:=	'0';
		dbg_dfx_clk	:	in	std_logic	:=	'0';
		dbg_dfx_sel	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		dbg_jtg_cdr	:	in	std_logic	:=	'0';
		dbg_jtg_ir_in	:	in	std_logic_vector(1 downto 0)	:=	"00";
		dbg_jtg_rti	:	in	std_logic	:=	'0';
		dbg_jtg_sdr	:	in	std_logic	:=	'0';
		dbg_jtg_tck	:	in	std_logic	:=	'0';
		dbg_jtg_tdi	:	in	std_logic	:=	'0';
		dbg_jtg_udr	:	in	std_logic	:=	'0';
		dbg_jtg_uir	:	in	std_logic	:=	'0';
		dft_clk	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		partial_reconfig	:	in	std_logic	:=	'0';
		soft_nios_addr	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		soft_nios_clk	:	in	std_logic	:=	'0';
		soft_nios_read	:	in	std_logic	:=	'0';
		soft_nios_write	:	in	std_logic	:=	'0';
		soft_nios_writedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		core_avl_addr	:	out	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		core_avl_burstcount	:	out	std_logic	:=	'0';
		core_avl_byteenable	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		core_avl_debugaccess	:	out	std_logic	:=	'0';
		core_avl_read	:	out	std_logic	:=	'0';
		core_avl_write	:	out	std_logic	:=	'0';
		core_avl_writedata	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		core_interrupt_out	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		dbg_dfx_out	:	out	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		dbg_jtg_ir_out	:	out	std_logic_vector(1 downto 0)	:=	"00";
		dbg_jtg_tdo	:	out	std_logic	:=	'0';
		dft_flag_down	:	out	std_logic	:=	'0';
		dft_flag_up	:	out	std_logic	:=	'0';
		soft_nios_readdata	:	out	std_logic_vector(7 downto 0)	:=	"00000000"
	);
end twentynm_hssi_pma_uc;

architecture behavior of twentynm_hssi_pma_uc	is

constant a_break_vector_word_addr_int	:	integer	:=	bin2int(a_break_vector_word_addr);
constant a_exception_vector_word_addr_int	:	integer	:=	bin2int(a_exception_vector_word_addr);
constant a_reset_vector_word_addr_int	:	integer	:=	bin2int(a_reset_vector_word_addr);
constant pm_uc_aux_base_addr_int	:	integer	:=	bin2int(pm_uc_aux_base_addr);
constant pm_uc_cal_clk_div_int	:	integer	:=	bin2int(pm_uc_cal_clk_div);
constant pm_uc_cal_clk_ph_int	:	integer	:=	bin2int(pm_uc_cal_clk_ph);
constant pm_uc_family_device_info_int	:	integer	:=	bin2int(pm_uc_family_device_info);
constant pm_uc_hssi_base_addr_int	:	integer	:=	bin2int(pm_uc_hssi_base_addr);
constant pm_uc_pcs_dft_out_int	:	integer	:=	bin2int(pm_uc_pcs_dft_out);
constant pm_uc_pcs_rd_lat_int	:	integer	:=	bin2int(pm_uc_pcs_rd_lat);
constant pm_uc_pcs_slave_count_int	:	integer	:=	bin2int(pm_uc_pcs_slave_count);



component	twentynm_hssi_pma_uc_encrypted
	generic (
		-- Architecture parameters
		a_break_vector_word_addr	:	integer	:=	8;
		a_exception_vector_word_addr	:	integer	:=	8;
		a_reset_vector_word_addr	:	integer	:=	0;
		cal_mode	:	string	:=	"cal_en";
		pm_uc_aux_base_addr	:	integer	:=	0;
		pm_uc_cal_clk_div	:	integer	:=	4;
		pm_uc_cal_clk_inv	:	string	:=	"disable_inv";
		pm_uc_cal_clk_ph	:	integer	:=	2;
		pm_uc_clkdiv_sel	:	string	:=	"div2";
		pm_uc_clksel_core	:	string	:=	"disable_core_clk";
		pm_uc_clksel_osc	:	string	:=	"cb_clkusr";
		pm_uc_core_jtg_rst_disable	:	string	:=	"disable_jtg_rst";
		pm_uc_core_sys_rst_disable	:	string	:=	"disable_core_rst";
		pm_uc_ecc_rst_disable	:	string	:=	"enable_ecc_rst";
		pm_uc_engg_opt	:	string	:=	"reserved";
		pm_uc_family_device_info	:	integer	:=	0;
		pm_uc_hssi_base_addr	:	integer	:=	1;
		pm_uc_pcs_dft_out	:	integer	:=	0;
		pm_uc_pcs_dft_sel	:	string	:=	"disable_pcs_dft";
		pm_uc_pcs_rd_lat	:	integer	:=	2;
		pm_uc_pcs_slave_count	:	integer	:=	0;
		pm_uc_ram	:	string	:=	"00000000000000000000000000000000000000";
		pm_uc_rmw_dis	:	string	:=	"enable_rmw";
		pm_uc_soft_nios	:	string	:=	"disable_soft";
		pm_uc_sys_enable	:	string	:=	"enable_sys";
		pmu_cal_bin_fname	:	string	:=	"nf_hssi_cal_v10.hex'";
		pmu_qparam_fname	:	string	:=	"nf_qparam_nf1.hex'";
		powerdown_mode	:	string	:=	"powerdown";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode"
	);
	port (
		-- Architecture ports
		cb_clkusr	:	in	std_logic	:=	'0';
		cb_intosc	:	in	std_logic	:=	'0';
		core_avl_clk	:	in	std_logic	:=	'0';
		core_avl_readdata	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		core_avl_readdatavalid	:	in	std_logic	:=	'0';
		core_avl_rst_n	:	in	std_logic	:=	'0';
		core_avl_waitrequest	:	in	std_logic	:=	'0';
		core_interrupt_in	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		core_uc_rst_n	:	in	std_logic	:=	'0';
		dbg_dfx_clk	:	in	std_logic	:=	'0';
		dbg_dfx_sel	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		dbg_jtg_cdr	:	in	std_logic	:=	'0';
		dbg_jtg_ir_in	:	in	std_logic_vector(1 downto 0)	:=	"00";
		dbg_jtg_rti	:	in	std_logic	:=	'0';
		dbg_jtg_sdr	:	in	std_logic	:=	'0';
		dbg_jtg_tck	:	in	std_logic	:=	'0';
		dbg_jtg_tdi	:	in	std_logic	:=	'0';
		dbg_jtg_udr	:	in	std_logic	:=	'0';
		dbg_jtg_uir	:	in	std_logic	:=	'0';
		dft_clk	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		partial_reconfig	:	in	std_logic	:=	'0';
		soft_nios_addr	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		soft_nios_clk	:	in	std_logic	:=	'0';
		soft_nios_read	:	in	std_logic	:=	'0';
		soft_nios_write	:	in	std_logic	:=	'0';
		soft_nios_writedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		core_avl_addr	:	out	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		core_avl_burstcount	:	out	std_logic	:=	'0';
		core_avl_byteenable	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		core_avl_debugaccess	:	out	std_logic	:=	'0';
		core_avl_read	:	out	std_logic	:=	'0';
		core_avl_write	:	out	std_logic	:=	'0';
		core_avl_writedata	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		core_interrupt_out	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		dbg_dfx_out	:	out	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		dbg_jtg_ir_out	:	out	std_logic_vector(1 downto 0)	:=	"00";
		dbg_jtg_tdo	:	out	std_logic	:=	'0';
		dft_flag_down	:	out	std_logic	:=	'0';
		dft_flag_up	:	out	std_logic	:=	'0';
		soft_nios_readdata	:	out	std_logic_vector(7 downto 0)	:=	"00000000"
	);
end component;

begin



inst : twentynm_hssi_pma_uc_encrypted
	generic map (
		-- Instance parameters
		a_break_vector_word_addr	=>	a_break_vector_word_addr_int,
		a_exception_vector_word_addr	=>	a_exception_vector_word_addr_int,
		a_reset_vector_word_addr	=>	a_reset_vector_word_addr_int,
		cal_mode	=>	cal_mode,
		pm_uc_aux_base_addr	=>	pm_uc_aux_base_addr_int,
		pm_uc_cal_clk_div	=>	pm_uc_cal_clk_div_int,
		pm_uc_cal_clk_inv	=>	pm_uc_cal_clk_inv,
		pm_uc_cal_clk_ph	=>	pm_uc_cal_clk_ph_int,
		pm_uc_clkdiv_sel	=>	pm_uc_clkdiv_sel,
		pm_uc_clksel_core	=>	pm_uc_clksel_core,
		pm_uc_clksel_osc	=>	pm_uc_clksel_osc,
		pm_uc_core_jtg_rst_disable	=>	pm_uc_core_jtg_rst_disable,
		pm_uc_core_sys_rst_disable	=>	pm_uc_core_sys_rst_disable,
		pm_uc_ecc_rst_disable	=>	pm_uc_ecc_rst_disable,
		pm_uc_engg_opt	=>	pm_uc_engg_opt,
		pm_uc_family_device_info	=>	pm_uc_family_device_info_int,
		pm_uc_hssi_base_addr	=>	pm_uc_hssi_base_addr_int,
		pm_uc_pcs_dft_out	=>	pm_uc_pcs_dft_out_int,
		pm_uc_pcs_dft_sel	=>	pm_uc_pcs_dft_sel,
		pm_uc_pcs_rd_lat	=>	pm_uc_pcs_rd_lat_int,
		pm_uc_pcs_slave_count	=>	pm_uc_pcs_slave_count_int,
		pm_uc_ram	=>	pm_uc_ram,
		pm_uc_rmw_dis	=>	pm_uc_rmw_dis,
		pm_uc_soft_nios	=>	pm_uc_soft_nios,
		pm_uc_sys_enable	=>	pm_uc_sys_enable,
		pmu_cal_bin_fname	=>	pmu_cal_bin_fname,
		pmu_qparam_fname	=>	pmu_qparam_fname,
		powerdown_mode	=>	powerdown_mode,
		silicon_rev	=>	silicon_rev,
		sup_mode	=>	sup_mode
	)
	port map (
		-- Instance ports
		cb_clkusr	=>	cb_clkusr,
		cb_intosc	=>	cb_intosc,
		core_avl_clk	=>	core_avl_clk,
		core_avl_readdata	=>	core_avl_readdata,
		core_avl_readdatavalid	=>	core_avl_readdatavalid,
		core_avl_rst_n	=>	core_avl_rst_n,
		core_avl_waitrequest	=>	core_avl_waitrequest,
		core_interrupt_in	=>	core_interrupt_in,
		core_uc_rst_n	=>	core_uc_rst_n,
		dbg_dfx_clk	=>	dbg_dfx_clk,
		dbg_dfx_sel	=>	dbg_dfx_sel,
		dbg_jtg_cdr	=>	dbg_jtg_cdr,
		dbg_jtg_ir_in	=>	dbg_jtg_ir_in,
		dbg_jtg_rti	=>	dbg_jtg_rti,
		dbg_jtg_sdr	=>	dbg_jtg_sdr,
		dbg_jtg_tck	=>	dbg_jtg_tck,
		dbg_jtg_tdi	=>	dbg_jtg_tdi,
		dbg_jtg_udr	=>	dbg_jtg_udr,
		dbg_jtg_uir	=>	dbg_jtg_uir,
		dft_clk	=>	dft_clk,
		partial_reconfig	=>	partial_reconfig,
		soft_nios_addr	=>	soft_nios_addr,
		soft_nios_clk	=>	soft_nios_clk,
		soft_nios_read	=>	soft_nios_read,
		soft_nios_write	=>	soft_nios_write,
		soft_nios_writedata	=>	soft_nios_writedata,
		core_avl_addr	=>	core_avl_addr,
		core_avl_burstcount	=>	core_avl_burstcount,
		core_avl_byteenable	=>	core_avl_byteenable,
		core_avl_debugaccess	=>	core_avl_debugaccess,
		core_avl_read	=>	core_avl_read,
		core_avl_write	=>	core_avl_write,
		core_avl_writedata	=>	core_avl_writedata,
		core_interrupt_out	=>	core_interrupt_out,
		dbg_dfx_out	=>	dbg_dfx_out,
		dbg_jtg_ir_out	=>	dbg_jtg_ir_out,
		dbg_jtg_tdo	=>	dbg_jtg_tdo,
		dft_flag_down	=>	dft_flag_down,
		dft_flag_up	=>	dft_flag_up,
		soft_nios_readdata	=>	soft_nios_readdata
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_refclk_divider	is
	generic (
		-- Entity parameters
		clk_divider	:	string	:=	"div2_off";
		clkbuf_sel	:	string	:=	"high_vcm";
		core_clk_lvpecl	:	string	:=	"core_clk_lvpecl_off";
		enable_lvpecl	:	string	:=	"lvpecl_enable";
		iostandard	:	string	:=	"lvpecl";
		optimal	:	string	:=	"true";
		powerdown_mode	:	string	:=	"powerup";
		sel_pldclk	:	string	:=	"iqclk_sel_lvpecl";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode";
		term_tristate	:	string	:=	"tristate_off";
		vcm_pup	:	string	:=	"pup_off"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		ac_mode	:	in	std_logic	:=	'0';
		atb_0_bidir_in	:	in	std_logic	:=	'0';
		atb_1_bidir_in	:	in	std_logic	:=	'0';
		atbsel_lvpecl	:	in	std_logic	:=	'0';
		clkbuf_b50	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		highz	:	in	std_logic	:=	'0';
		hotsckt	:	in	std_logic	:=	'0';
		mem_init	:	in	std_logic	:=	'0';
		mode	:	in	std_logic	:=	'0';
		pldclk	:	in	std_logic	:=	'0';
		refclk_inn	:	in	std_logic	:=	'0';
		refclk_inp	:	in	std_logic	:=	'0';
		refclk_n	:	in	std_logic	:=	'0';
		refclk_p	:	in	std_logic	:=	'0';
		rjdrv_sel	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rjhys_sel	:	in	std_logic	:=	'0';
		rjtaglp	:	in	std_logic	:=	'0';
		vlprxn	:	in	std_logic	:=	'0';
		vlprxp	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		bsrefclkn	:	out	std_logic	:=	'0';
		bsrefclkp	:	out	std_logic	:=	'0';
		refclk_a	:	out	std_logic	:=	'0'
	);
end twentynm_hssi_refclk_divider;

architecture behavior of twentynm_hssi_refclk_divider	is




component	twentynm_hssi_refclk_divider_encrypted
	generic (
		-- Architecture parameters
		clk_divider	:	string	:=	"div2_off";
		clkbuf_sel	:	string	:=	"high_vcm";
		core_clk_lvpecl	:	string	:=	"core_clk_lvpecl_off";
		enable_lvpecl	:	string	:=	"lvpecl_enable";
		iostandard	:	string	:=	"lvpecl";
		optimal	:	string	:=	"true";
		powerdown_mode	:	string	:=	"powerup";
		sel_pldclk	:	string	:=	"iqclk_sel_lvpecl";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode";
		term_tristate	:	string	:=	"tristate_off";
		vcm_pup	:	string	:=	"pup_off"
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		ac_mode	:	in	std_logic	:=	'0';
		atb_0_bidir_in	:	in	std_logic	:=	'0';
		atb_1_bidir_in	:	in	std_logic	:=	'0';
		atbsel_lvpecl	:	in	std_logic	:=	'0';
		clkbuf_b50	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		highz	:	in	std_logic	:=	'0';
		hotsckt	:	in	std_logic	:=	'0';
		mem_init	:	in	std_logic	:=	'0';
		mode	:	in	std_logic	:=	'0';
		pldclk	:	in	std_logic	:=	'0';
		refclk_inn	:	in	std_logic	:=	'0';
		refclk_inp	:	in	std_logic	:=	'0';
		refclk_n	:	in	std_logic	:=	'0';
		refclk_p	:	in	std_logic	:=	'0';
		rjdrv_sel	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rjhys_sel	:	in	std_logic	:=	'0';
		rjtaglp	:	in	std_logic	:=	'0';
		vlprxn	:	in	std_logic	:=	'0';
		vlprxp	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		bsrefclkn	:	out	std_logic	:=	'0';
		bsrefclkp	:	out	std_logic	:=	'0';
		refclk_a	:	out	std_logic	:=	'0'
	);
end component;

begin



inst : twentynm_hssi_refclk_divider_encrypted
	generic map (
		-- Instance parameters
		clk_divider	=>	clk_divider,
		clkbuf_sel	=>	clkbuf_sel,
		core_clk_lvpecl	=>	core_clk_lvpecl,
		enable_lvpecl	=>	enable_lvpecl,
		iostandard	=>	iostandard,
		optimal	=>	optimal,
		powerdown_mode	=>	powerdown_mode,
		sel_pldclk	=>	sel_pldclk,
		silicon_rev	=>	silicon_rev,
		sup_mode	=>	sup_mode,
		term_tristate	=>	term_tristate,
		vcm_pup	=>	vcm_pup
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		ac_mode	=>	ac_mode,
		atb_0_bidir_in	=>	atb_0_bidir_in,
		atb_1_bidir_in	=>	atb_1_bidir_in,
		atbsel_lvpecl	=>	atbsel_lvpecl,
		clkbuf_b50	=>	clkbuf_b50,
		highz	=>	highz,
		hotsckt	=>	hotsckt,
		mem_init	=>	mem_init,
		mode	=>	mode,
		pldclk	=>	pldclk,
		refclk_inn	=>	refclk_inn,
		refclk_inp	=>	refclk_inp,
		refclk_n	=>	refclk_n,
		refclk_p	=>	refclk_p,
		rjdrv_sel	=>	rjdrv_sel,
		rjhys_sel	=>	rjhys_sel,
		rjtaglp	=>	rjtaglp,
		vlprxn	=>	vlprxn,
		vlprxp	=>	vlprxp,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		bsrefclkn	=>	bsrefclkn,
		bsrefclkp	=>	bsrefclkp,
		refclk_a	=>	refclk_a
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_rx_pcs_pma_interface	is
	generic (
		-- Entity parameters
		block_sel	:	string	:=	"eight_g_pcs";
		channel_operation_mode	:	string	:=	"tx_rx_pair_enabled";
		clkslip_sel	:	string	:=	"pld";
		lpbk_en	:	string	:=	"disable";
		master_clk_sel	:	string	:=	"master_rx_pma_clk";
		pldif_datawidth_mode	:	string	:=	"pldif_data_10bit";
		pma_dw_rx	:	string	:=	"pma_8b_rx";
		pma_if_dft_en	:	string	:=	"dft_dis";
		pma_if_dft_val	:	string	:=	"dft_0";
		prbs9_dwidth	:	string	:=	"prbs9_64b";
		prbs_clken	:	string	:=	"prbs_clk_dis";
		prbs_ver	:	string	:=	"prbs_off";
		prot_mode_rx	:	string	:=	"disabled_prot_mode_rx";
		reconfig_settings	:	string	:=	"{}";
		rx_dyn_polarity_inversion	:	string	:=	"rx_dyn_polinv_dis";
		rx_lpbk_en	:	string	:=	"lpbk_dis";
		rx_prbs_force_signal_ok	:	string	:=	"unforce_sig_ok";
		rx_prbs_mask	:	string	:=	"prbsmask128";
		rx_prbs_mode	:	string	:=	"teng_mode";
		rx_signalok_signaldet_sel	:	string	:=	"sel_sig_det";
		rx_static_polarity_inversion	:	string	:=	"rx_stat_polinv_dis";
		rx_uhsif_lpbk_en	:	string	:=	"uhsif_lpbk_dis";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		int_pmaif_10g_random_err	:	in	std_logic	:=	'0';
		int_pmaif_8g_rx_clkslip	:	in	std_logic	:=	'0';
		int_pmaif_pldif_eye_monitor	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		int_pmaif_pldif_pmaif_rx_pld_rst_n	:	in	std_logic	:=	'0';
		int_pmaif_pldif_polinv_rx	:	in	std_logic	:=	'0';
		int_pmaif_pldif_prbs_err_clr	:	in	std_logic	:=	'0';
		int_pmaif_pldif_rx_clkslip	:	in	std_logic	:=	'0';
		int_pmaif_pldif_rxpma_rstb	:	in	std_logic	:=	'0';
		pma_rx_clkdiv_user	:	in	std_logic	:=	'0';
		pma_rx_detect_valid	:	in	std_logic	:=	'0';
		pma_rx_found	:	in	std_logic	:=	'0';
		pma_rx_pma_clk	:	in	std_logic	:=	'0';
		pma_rx_pma_data	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		pma_rx_signal_ok	:	in	std_logic	:=	'0';
		pma_rxpll_lock	:	in	std_logic	:=	'0';
		pma_signal_det	:	in	std_logic	:=	'0';
		pma_tx_pma_clk	:	in	std_logic	:=	'0';
		refclk_dig	:	in	std_logic	:=	'0';
		scan_mode_n	:	in	std_logic	:=	'0';
		tx_pma_data_loopback	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		tx_pma_uhsif_data_loopback	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		int_pmaif_10g_rx_pma_clk	:	out	std_logic	:=	'0';
		int_pmaif_10g_rx_pma_data	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		int_pmaif_10g_signal_ok	:	out	std_logic	:=	'0';
		int_pmaif_8g_pudi	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		int_pmaif_8g_rcvd_clk_pma	:	out	std_logic	:=	'0';
		int_pmaif_8g_rx_detect_valid	:	out	std_logic	:=	'0';
		int_pmaif_8g_rx_found	:	out	std_logic	:=	'0';
		int_pmaif_8g_sigdetni	:	out	std_logic	:=	'0';
		int_pmaif_g3_pma_data_in	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		int_pmaif_g3_pma_rx_detect_valid	:	out	std_logic	:=	'0';
		int_pmaif_g3_pma_rx_found	:	out	std_logic	:=	'0';
		int_pmaif_g3_pma_signal_det	:	out	std_logic	:=	'0';
		int_pmaif_g3_rcvd_clk	:	out	std_logic	:=	'0';
		int_pmaif_krfec_rx_pma_data	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		int_pmaif_krfec_rx_signal_ok_in	:	out	std_logic	:=	'0';
		int_pmaif_pldif_prbs_err	:	out	std_logic	:=	'0';
		int_pmaif_pldif_prbs_err_done	:	out	std_logic	:=	'0';
		int_pmaif_pldif_rx_clkdiv	:	out	std_logic	:=	'0';
		int_pmaif_pldif_rx_clkdiv_user	:	out	std_logic	:=	'0';
		int_pmaif_pldif_rx_data	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		int_pmaif_pldif_rx_detect_valid	:	out	std_logic	:=	'0';
		int_pmaif_pldif_rx_found	:	out	std_logic	:=	'0';
		int_pmaif_pldif_rxpll_lock	:	out	std_logic	:=	'0';
		int_pmaif_pldif_signal_ok	:	out	std_logic	:=	'0';
		int_rx_dft_obsrv_clk	:	out	std_logic	:=	'0';
		pma_eye_monitor	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		pma_rx_clkslip	:	out	std_logic	:=	'0';
		pma_rxpma_rstb	:	out	std_logic	:=	'0';
		prbs_err_lt	:	out	std_logic	:=	'0';
		rx_pmaif_test_out	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		rx_prbs_ver_test	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000"
	);
end twentynm_hssi_rx_pcs_pma_interface;

architecture behavior of twentynm_hssi_rx_pcs_pma_interface	is




component	twentynm_hssi_rx_pcs_pma_interface_encrypted
	generic (
		-- Architecture parameters
		block_sel	:	string	:=	"eight_g_pcs";
		channel_operation_mode	:	string	:=	"tx_rx_pair_enabled";
		clkslip_sel	:	string	:=	"pld";
		lpbk_en	:	string	:=	"disable";
		master_clk_sel	:	string	:=	"master_rx_pma_clk";
		pldif_datawidth_mode	:	string	:=	"pldif_data_10bit";
		pma_dw_rx	:	string	:=	"pma_8b_rx";
		pma_if_dft_en	:	string	:=	"dft_dis";
		pma_if_dft_val	:	string	:=	"dft_0";
		prbs9_dwidth	:	string	:=	"prbs9_64b";
		prbs_clken	:	string	:=	"prbs_clk_dis";
		prbs_ver	:	string	:=	"prbs_off";
		prot_mode_rx	:	string	:=	"disabled_prot_mode_rx";
		reconfig_settings	:	string	:=	"{}";
		rx_dyn_polarity_inversion	:	string	:=	"rx_dyn_polinv_dis";
		rx_lpbk_en	:	string	:=	"lpbk_dis";
		rx_prbs_force_signal_ok	:	string	:=	"unforce_sig_ok";
		rx_prbs_mask	:	string	:=	"prbsmask128";
		rx_prbs_mode	:	string	:=	"teng_mode";
		rx_signalok_signaldet_sel	:	string	:=	"sel_sig_det";
		rx_static_polarity_inversion	:	string	:=	"rx_stat_polinv_dis";
		rx_uhsif_lpbk_en	:	string	:=	"uhsif_lpbk_dis";
		silicon_rev	:	string	:=	"20nm5es";
		sup_mode	:	string	:=	"user_mode"
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		int_pmaif_10g_random_err	:	in	std_logic	:=	'0';
		int_pmaif_8g_rx_clkslip	:	in	std_logic	:=	'0';
		int_pmaif_pldif_eye_monitor	:	in	std_logic_vector(5 downto 0)	:=	"000000";
		int_pmaif_pldif_pmaif_rx_pld_rst_n	:	in	std_logic	:=	'0';
		int_pmaif_pldif_polinv_rx	:	in	std_logic	:=	'0';
		int_pmaif_pldif_prbs_err_clr	:	in	std_logic	:=	'0';
		int_pmaif_pldif_rx_clkslip	:	in	std_logic	:=	'0';
		int_pmaif_pldif_rxpma_rstb	:	in	std_logic	:=	'0';
		pma_rx_clkdiv_user	:	in	std_logic	:=	'0';
		pma_rx_detect_valid	:	in	std_logic	:=	'0';
		pma_rx_found	:	in	std_logic	:=	'0';
		pma_rx_pma_clk	:	in	std_logic	:=	'0';
		pma_rx_pma_data	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		pma_rx_signal_ok	:	in	std_logic	:=	'0';
		pma_rxpll_lock	:	in	std_logic	:=	'0';
		pma_signal_det	:	in	std_logic	:=	'0';
		pma_tx_pma_clk	:	in	std_logic	:=	'0';
		refclk_dig	:	in	std_logic	:=	'0';
		scan_mode_n	:	in	std_logic	:=	'0';
		tx_pma_data_loopback	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		tx_pma_uhsif_data_loopback	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		int_pmaif_10g_rx_pma_clk	:	out	std_logic	:=	'0';
		int_pmaif_10g_rx_pma_data	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		int_pmaif_10g_signal_ok	:	out	std_logic	:=	'0';
		int_pmaif_8g_pudi	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		int_pmaif_8g_rcvd_clk_pma	:	out	std_logic	:=	'0';
		int_pmaif_8g_rx_detect_valid	:	out	std_logic	:=	'0';
		int_pmaif_8g_rx_found	:	out	std_logic	:=	'0';
		int_pmaif_8g_sigdetni	:	out	std_logic	:=	'0';
		int_pmaif_g3_pma_data_in	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		int_pmaif_g3_pma_rx_detect_valid	:	out	std_logic	:=	'0';
		int_pmaif_g3_pma_rx_found	:	out	std_logic	:=	'0';
		int_pmaif_g3_pma_signal_det	:	out	std_logic	:=	'0';
		int_pmaif_g3_rcvd_clk	:	out	std_logic	:=	'0';
		int_pmaif_krfec_rx_pma_data	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		int_pmaif_krfec_rx_signal_ok_in	:	out	std_logic	:=	'0';
		int_pmaif_pldif_prbs_err	:	out	std_logic	:=	'0';
		int_pmaif_pldif_prbs_err_done	:	out	std_logic	:=	'0';
		int_pmaif_pldif_rx_clkdiv	:	out	std_logic	:=	'0';
		int_pmaif_pldif_rx_clkdiv_user	:	out	std_logic	:=	'0';
		int_pmaif_pldif_rx_data	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		int_pmaif_pldif_rx_detect_valid	:	out	std_logic	:=	'0';
		int_pmaif_pldif_rx_found	:	out	std_logic	:=	'0';
		int_pmaif_pldif_rxpll_lock	:	out	std_logic	:=	'0';
		int_pmaif_pldif_signal_ok	:	out	std_logic	:=	'0';
		int_rx_dft_obsrv_clk	:	out	std_logic	:=	'0';
		pma_eye_monitor	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		pma_rx_clkslip	:	out	std_logic	:=	'0';
		pma_rxpma_rstb	:	out	std_logic	:=	'0';
		prbs_err_lt	:	out	std_logic	:=	'0';
		rx_pmaif_test_out	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		rx_prbs_ver_test	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000"
	);
end component;

begin



inst : twentynm_hssi_rx_pcs_pma_interface_encrypted
	generic map (
		-- Instance parameters
		block_sel	=>	block_sel,
		channel_operation_mode	=>	channel_operation_mode,
		clkslip_sel	=>	clkslip_sel,
		lpbk_en	=>	lpbk_en,
		master_clk_sel	=>	master_clk_sel,
		pldif_datawidth_mode	=>	pldif_datawidth_mode,
		pma_dw_rx	=>	pma_dw_rx,
		pma_if_dft_en	=>	pma_if_dft_en,
		pma_if_dft_val	=>	pma_if_dft_val,
		prbs9_dwidth	=>	prbs9_dwidth,
		prbs_clken	=>	prbs_clken,
		prbs_ver	=>	prbs_ver,
		prot_mode_rx	=>	prot_mode_rx,
		reconfig_settings	=>	reconfig_settings,
		rx_dyn_polarity_inversion	=>	rx_dyn_polarity_inversion,
		rx_lpbk_en	=>	rx_lpbk_en,
		rx_prbs_force_signal_ok	=>	rx_prbs_force_signal_ok,
		rx_prbs_mask	=>	rx_prbs_mask,
		rx_prbs_mode	=>	rx_prbs_mode,
		rx_signalok_signaldet_sel	=>	rx_signalok_signaldet_sel,
		rx_static_polarity_inversion	=>	rx_static_polarity_inversion,
		rx_uhsif_lpbk_en	=>	rx_uhsif_lpbk_en,
		silicon_rev	=>	silicon_rev,
		sup_mode	=>	sup_mode
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		int_pmaif_10g_random_err	=>	int_pmaif_10g_random_err,
		int_pmaif_8g_rx_clkslip	=>	int_pmaif_8g_rx_clkslip,
		int_pmaif_pldif_eye_monitor	=>	int_pmaif_pldif_eye_monitor,
		int_pmaif_pldif_pmaif_rx_pld_rst_n	=>	int_pmaif_pldif_pmaif_rx_pld_rst_n,
		int_pmaif_pldif_polinv_rx	=>	int_pmaif_pldif_polinv_rx,
		int_pmaif_pldif_prbs_err_clr	=>	int_pmaif_pldif_prbs_err_clr,
		int_pmaif_pldif_rx_clkslip	=>	int_pmaif_pldif_rx_clkslip,
		int_pmaif_pldif_rxpma_rstb	=>	int_pmaif_pldif_rxpma_rstb,
		pma_rx_clkdiv_user	=>	pma_rx_clkdiv_user,
		pma_rx_detect_valid	=>	pma_rx_detect_valid,
		pma_rx_found	=>	pma_rx_found,
		pma_rx_pma_clk	=>	pma_rx_pma_clk,
		pma_rx_pma_data	=>	pma_rx_pma_data,
		pma_rx_signal_ok	=>	pma_rx_signal_ok,
		pma_rxpll_lock	=>	pma_rxpll_lock,
		pma_signal_det	=>	pma_signal_det,
		pma_tx_pma_clk	=>	pma_tx_pma_clk,
		refclk_dig	=>	refclk_dig,
		scan_mode_n	=>	scan_mode_n,
		tx_pma_data_loopback	=>	tx_pma_data_loopback,
		tx_pma_uhsif_data_loopback	=>	tx_pma_uhsif_data_loopback,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		int_pmaif_10g_rx_pma_clk	=>	int_pmaif_10g_rx_pma_clk,
		int_pmaif_10g_rx_pma_data	=>	int_pmaif_10g_rx_pma_data,
		int_pmaif_10g_signal_ok	=>	int_pmaif_10g_signal_ok,
		int_pmaif_8g_pudi	=>	int_pmaif_8g_pudi,
		int_pmaif_8g_rcvd_clk_pma	=>	int_pmaif_8g_rcvd_clk_pma,
		int_pmaif_8g_rx_detect_valid	=>	int_pmaif_8g_rx_detect_valid,
		int_pmaif_8g_rx_found	=>	int_pmaif_8g_rx_found,
		int_pmaif_8g_sigdetni	=>	int_pmaif_8g_sigdetni,
		int_pmaif_g3_pma_data_in	=>	int_pmaif_g3_pma_data_in,
		int_pmaif_g3_pma_rx_detect_valid	=>	int_pmaif_g3_pma_rx_detect_valid,
		int_pmaif_g3_pma_rx_found	=>	int_pmaif_g3_pma_rx_found,
		int_pmaif_g3_pma_signal_det	=>	int_pmaif_g3_pma_signal_det,
		int_pmaif_g3_rcvd_clk	=>	int_pmaif_g3_rcvd_clk,
		int_pmaif_krfec_rx_pma_data	=>	int_pmaif_krfec_rx_pma_data,
		int_pmaif_krfec_rx_signal_ok_in	=>	int_pmaif_krfec_rx_signal_ok_in,
		int_pmaif_pldif_prbs_err	=>	int_pmaif_pldif_prbs_err,
		int_pmaif_pldif_prbs_err_done	=>	int_pmaif_pldif_prbs_err_done,
		int_pmaif_pldif_rx_clkdiv	=>	int_pmaif_pldif_rx_clkdiv,
		int_pmaif_pldif_rx_clkdiv_user	=>	int_pmaif_pldif_rx_clkdiv_user,
		int_pmaif_pldif_rx_data	=>	int_pmaif_pldif_rx_data,
		int_pmaif_pldif_rx_detect_valid	=>	int_pmaif_pldif_rx_detect_valid,
		int_pmaif_pldif_rx_found	=>	int_pmaif_pldif_rx_found,
		int_pmaif_pldif_rxpll_lock	=>	int_pmaif_pldif_rxpll_lock,
		int_pmaif_pldif_signal_ok	=>	int_pmaif_pldif_signal_ok,
		int_rx_dft_obsrv_clk	=>	int_rx_dft_obsrv_clk,
		pma_eye_monitor	=>	pma_eye_monitor,
		pma_rx_clkslip	=>	pma_rx_clkslip,
		pma_rxpma_rstb	=>	pma_rxpma_rstb,
		prbs_err_lt	=>	prbs_err_lt,
		rx_pmaif_test_out	=>	rx_pmaif_test_out,
		rx_prbs_ver_test	=>	rx_prbs_ver_test
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_rx_pld_pcs_interface	is
	generic (
		-- Entity parameters
		hd_10g_advanced_user_mode_rx	:	string	:=	"disable";
		hd_10g_channel_operation_mode	:	string	:=	"tx_rx_pair_enabled";
		hd_10g_ctrl_plane_bonding_rx	:	string	:=	"individual_rx";
		hd_10g_fifo_mode_rx	:	string	:=	"fifo_rx";
		hd_10g_low_latency_en_rx	:	string	:=	"enable";
		hd_10g_lpbk_en	:	string	:=	"disable";
		hd_10g_pma_dw_rx	:	string	:=	"pma_64b_rx";
		hd_10g_prot_mode_rx	:	string	:=	"disabled_prot_mode_rx";
		hd_10g_shared_fifo_width_rx	:	string	:=	"single_rx";
		hd_10g_sup_mode	:	string	:=	"user_mode";
		hd_10g_test_bus_mode	:	string	:=	"tx";
		hd_8g_channel_operation_mode	:	string	:=	"tx_rx_pair_enabled";
		hd_8g_ctrl_plane_bonding_rx	:	string	:=	"individual_rx";
		hd_8g_fifo_mode_rx	:	string	:=	"fifo_rx";
		hd_8g_hip_mode	:	string	:=	"disable";
		hd_8g_lpbk_en	:	string	:=	"disable";
		hd_8g_pma_dw_rx	:	string	:=	"pma_8b_rx";
		hd_8g_prot_mode_rx	:	string	:=	"disabled_prot_mode_rx";
		hd_8g_sup_mode	:	string	:=	"user_mode";
		hd_chnl_channel_operation_mode	:	string	:=	"tx_rx_pair_enabled";
		hd_chnl_clklow_clk_hz	:	bit_vector	:=	B"000000000000000000000000000000";
		hd_chnl_ctrl_plane_bonding_rx	:	string	:=	"individual_rx";
		hd_chnl_fref_clk_hz	:	bit_vector	:=	B"000000000000000000000000000000";
		hd_chnl_frequency_rules_en	:	string	:=	"disable";
		hd_chnl_func_mode	:	string	:=	"disable";
		hd_chnl_hclk_clk_hz	:	bit_vector	:=	B"000000000000000000000000000000";
		hd_chnl_hip_en	:	string	:=	"disable";
		hd_chnl_hrdrstctl_en	:	string	:=	"disable";
		hd_chnl_low_latency_en_rx	:	string	:=	"disable";
		hd_chnl_lpbk_en	:	string	:=	"disable";
		hd_chnl_operating_voltage	:	string	:=	"standard";
		hd_chnl_pcs_ac_pwr_rules_en	:	string	:=	"disable";
		hd_chnl_pcs_pair_ac_pwr_uw_per_mhz	:	bit_vector	:=	B"00000000000000000000";
		hd_chnl_pcs_rx_ac_pwr_uw_per_mhz	:	bit_vector	:=	B"00000000000000000000";
		hd_chnl_pcs_rx_pwr_scaling_clk	:	string	:=	"pma_rx_clk";
		hd_chnl_pld_8g_refclk_dig_nonatpg_mode_clk_hz	:	bit_vector	:=	B"000000000000000000000000000000";
		hd_chnl_pld_fifo_mode_rx	:	string	:=	"fifo_rx";
		hd_chnl_pld_pcs_refclk_dig_nonatpg_mode_clk_hz	:	bit_vector	:=	B"000000000000000000000000000000";
		hd_chnl_pld_rx_clk_hz	:	bit_vector	:=	B"000000000000000000000000000000";
		hd_chnl_pma_dw_rx	:	string	:=	"pma_8b_rx";
		hd_chnl_pma_rx_clk_hz	:	bit_vector	:=	B"000000000000000000000000000000";
		hd_chnl_prot_mode_rx	:	string	:=	"disabled_prot_mode_rx";
		hd_chnl_shared_fifo_width_rx	:	string	:=	"single_rx";
		hd_chnl_speed_grade	:	string	:=	"e2";
		hd_chnl_sup_mode	:	string	:=	"user_mode";
		hd_chnl_transparent_pcs_rx	:	string	:=	"disable";
		hd_fifo_channel_operation_mode	:	string	:=	"tx_rx_pair_enabled";
		hd_fifo_prot_mode_rx	:	string	:=	"teng_mode_rx";
		hd_fifo_shared_fifo_width_rx	:	string	:=	"single_rx";
		hd_fifo_sup_mode	:	string	:=	"user_mode";
		hd_g3_prot_mode	:	string	:=	"disabled_prot_mode";
		hd_g3_sup_mode	:	string	:=	"user_mode";
		hd_krfec_channel_operation_mode	:	string	:=	"tx_rx_pair_enabled";
		hd_krfec_low_latency_en_rx	:	string	:=	"disable";
		hd_krfec_lpbk_en	:	string	:=	"disable";
		hd_krfec_prot_mode_rx	:	string	:=	"disabled_prot_mode_rx";
		hd_krfec_sup_mode	:	string	:=	"user_mode";
		hd_krfec_test_bus_mode	:	string	:=	"tx";
		hd_pldif_hrdrstctl_en	:	string	:=	"disable";
		hd_pldif_prot_mode_rx	:	string	:=	"disabled_prot_mode_rx";
		hd_pldif_sup_mode	:	string	:=	"user_mode";
		hd_pmaif_channel_operation_mode	:	string	:=	"tx_rx_pair_enabled";
		hd_pmaif_lpbk_en	:	string	:=	"disable";
		hd_pmaif_pma_dw_rx	:	string	:=	"pma_8b_rx";
		hd_pmaif_prot_mode_rx	:	string	:=	"disabled_prot_mode_rx";
		hd_pmaif_sim_mode	:	string	:=	"disable";
		hd_pmaif_sup_mode	:	string	:=	"user_mode";
		pcs_rx_block_sel	:	string	:=	"pcs_direct";
		pcs_rx_clk_out_sel	:	string	:=	"teng_clk_out";
		pcs_rx_clk_sel	:	string	:=	"pld_rx_clk";
		pcs_rx_hip_clk_en	:	string	:=	"hip_rx_enable";
		pcs_rx_output_sel	:	string	:=	"teng_output";
		reconfig_settings	:	string	:=	"{}";
		silicon_rev	:	string	:=	"20nm5es"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		int_pldif_10g_rx_align_val	:	in	std_logic	:=	'0';
		int_pldif_10g_rx_blk_lock	:	in	std_logic	:=	'0';
		int_pldif_10g_rx_clk_out	:	in	std_logic	:=	'0';
		int_pldif_10g_rx_clk_out_pld_if	:	in	std_logic	:=	'0';
		int_pldif_10g_rx_control	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		int_pldif_10g_rx_crc32_err	:	in	std_logic	:=	'0';
		int_pldif_10g_rx_data	:	in	std_logic_vector(127 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		int_pldif_10g_rx_data_valid	:	in	std_logic	:=	'0';
		int_pldif_10g_rx_diag_status	:	in	std_logic_vector(1 downto 0)	:=	"00";
		int_pldif_10g_rx_empty	:	in	std_logic	:=	'0';
		int_pldif_10g_rx_fifo_del	:	in	std_logic	:=	'0';
		int_pldif_10g_rx_fifo_insert	:	in	std_logic	:=	'0';
		int_pldif_10g_rx_fifo_num	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		int_pldif_10g_rx_frame_lock	:	in	std_logic	:=	'0';
		int_pldif_10g_rx_hi_ber	:	in	std_logic	:=	'0';
		int_pldif_10g_rx_oflw_err	:	in	std_logic	:=	'0';
		int_pldif_10g_rx_pempty	:	in	std_logic	:=	'0';
		int_pldif_10g_rx_pfull	:	in	std_logic	:=	'0';
		int_pldif_10g_rx_rx_frame	:	in	std_logic	:=	'0';
		int_pldif_8g_a1a2_k1k2_flag	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		int_pldif_8g_empty_rmf	:	in	std_logic	:=	'0';
		int_pldif_8g_empty_rx	:	in	std_logic	:=	'0';
		int_pldif_8g_full_rmf	:	in	std_logic	:=	'0';
		int_pldif_8g_full_rx	:	in	std_logic	:=	'0';
		int_pldif_8g_phystatus	:	in	std_logic	:=	'0';
		int_pldif_8g_rx_blk_start	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		int_pldif_8g_rx_clk	:	in	std_logic	:=	'0';
		int_pldif_8g_rx_clk_out_pld_if	:	in	std_logic	:=	'0';
		int_pldif_8g_rx_data_valid	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		int_pldif_8g_rx_rstn_sync2wrfifo	:	in	std_logic	:=	'0';
		int_pldif_8g_rx_sync_hdr	:	in	std_logic_vector(1 downto 0)	:=	"00";
		int_pldif_8g_rxd	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		int_pldif_8g_rxelecidle	:	in	std_logic	:=	'0';
		int_pldif_8g_rxstatus	:	in	std_logic_vector(2 downto 0)	:=	"000";
		int_pldif_8g_rxvalid	:	in	std_logic	:=	'0';
		int_pldif_8g_signal_detect_out	:	in	std_logic	:=	'0';
		int_pldif_8g_wa_boundary	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		int_pldif_krfec_rx_block_lock	:	in	std_logic	:=	'0';
		int_pldif_krfec_rx_data_status	:	in	std_logic_vector(1 downto 0)	:=	"00";
		int_pldif_krfec_rx_frame	:	in	std_logic	:=	'0';
		int_pldif_pmaif_clkdiv_rx	:	in	std_logic	:=	'0';
		int_pldif_pmaif_clkdiv_rx_user	:	in	std_logic	:=	'0';
		int_pldif_pmaif_rx_data	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		int_pldif_pmaif_rx_prbs_done	:	in	std_logic	:=	'0';
		int_pldif_pmaif_rx_prbs_err	:	in	std_logic	:=	'0';
		int_pldif_pmaif_rxpll_lock	:	in	std_logic	:=	'0';
		int_pldif_pmaif_signal_ok	:	in	std_logic	:=	'0';
		int_pldif_usr_rst_sel	:	in	std_logic	:=	'0';
		pld_10g_krfec_rx_clr_errblk_cnt	:	in	std_logic	:=	'0';
		pld_10g_krfec_rx_pld_rst_n	:	in	std_logic	:=	'0';
		pld_10g_rx_align_clr	:	in	std_logic	:=	'0';
		pld_10g_rx_clr_ber_count	:	in	std_logic	:=	'0';
		pld_10g_rx_rd_en	:	in	std_logic	:=	'0';
		pld_8g_a1a2_size	:	in	std_logic	:=	'0';
		pld_8g_bitloc_rev_en	:	in	std_logic	:=	'0';
		pld_8g_byte_rev_en	:	in	std_logic	:=	'0';
		pld_8g_encdt	:	in	std_logic	:=	'0';
		pld_8g_g3_rx_pld_rst_n	:	in	std_logic	:=	'0';
		pld_8g_rdenable_rx	:	in	std_logic	:=	'0';
		pld_8g_rxpolarity	:	in	std_logic	:=	'0';
		pld_8g_wrdisable_rx	:	in	std_logic	:=	'0';
		pld_bitslip	:	in	std_logic	:=	'0';
		pld_partial_reconfig	:	in	std_logic	:=	'0';
		pld_pma_rxpma_rstb	:	in	std_logic	:=	'0';
		pld_pmaif_rx_pld_rst_n	:	in	std_logic	:=	'0';
		pld_pmaif_rxclkslip	:	in	std_logic	:=	'0';
		pld_polinv_rx	:	in	std_logic	:=	'0';
		pld_rx_clk	:	in	std_logic	:=	'0';
		pld_rx_prbs_err_clr	:	in	std_logic	:=	'0';
		pld_syncsm_en	:	in	std_logic	:=	'0';
		scan_mode_n	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		pld_8g_wa_boundary_txclk_fastreg	:	out	std_logic	:=	'0';
		pld_8g_wa_boundary_txclk_reg	:	out	std_logic	:=	'0';
		pld_bitslip_10g_txclk_reg	:	out	std_logic	:=	'0';
		pld_bitslip_8g_txclk_reg	:	out	std_logic	:=	'0';
		pld_bitslip_rxclk_parallel_loopback_reg	:	out	std_logic	:=	'0';
		pld_bitslip_rxclk_reg	:	out	std_logic	:=	'0';
		pld_pcs_rx_clk_out_pcsdirect_wire	:	out	std_logic	:=	'0';
		pld_pma_rx_clk_out_10g_or_pcsdirect_wire	:	out	std_logic	:=	'0';
		pld_pma_rx_clk_out_8g_wire	:	out	std_logic	:=	'0';
		pld_pmaif_rx_pld_rst_n_reg	:	out	std_logic	:=	'0';
		pld_pmaif_tx_pld_rst_n_txclk_reg	:	out	std_logic	:=	'0';
		pld_polinv_rx_reg	:	out	std_logic	:=	'0';
		pld_rx_clk_fifo	:	out	std_logic	:=	'0';
		pld_rx_control_fifo	:	out	std_logic	:=	'0';
		pld_rx_control_pcsdirect_reg	:	out	std_logic	:=	'0';
		pld_rx_data_fifo	:	out	std_logic	:=	'0';
		pld_rx_data_pcsdirect_reg	:	out	std_logic	:=	'0';
		pld_rx_prbs_done_reg	:	out	std_logic	:=	'0';
		pld_rx_prbs_done_txclk_reg	:	out	std_logic	:=	'0';
		pld_rx_prbs_err_clr_pcsdirect_txclk_reg	:	out	std_logic	:=	'0';
		pld_rx_prbs_err_clr_reg	:	out	std_logic	:=	'0';
		pld_rx_prbs_err_disprbs_reg	:	out	std_logic	:=	'0';
		pld_rx_prbs_err_pcsdirect_txclk_reg	:	out	std_logic	:=	'0';
		pld_rx_prbs_err_reg	:	out	std_logic	:=	'0';
		pma_rx_pma_clk_reg	:	out	std_logic	:=	'0';
		hip_rx_ctrl	:	out	std_logic_vector(1 downto 0)	:=	"00";
		hip_rx_data	:	out	std_logic_vector(50 downto 0)	:=	"000000000000000000000000000000000000000000000000000";
		int_pldif_10g_rx_align_clr	:	out	std_logic	:=	'0';
		int_pldif_10g_rx_bitslip	:	out	std_logic	:=	'0';
		int_pldif_10g_rx_clr_ber_count	:	out	std_logic	:=	'0';
		int_pldif_10g_rx_clr_errblk_cnt	:	out	std_logic	:=	'0';
		int_pldif_10g_rx_control_fb	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		int_pldif_10g_rx_data_fb	:	out	std_logic_vector(127 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		int_pldif_10g_rx_data_valid_fb	:	out	std_logic	:=	'0';
		int_pldif_10g_rx_pld_clk	:	out	std_logic	:=	'0';
		int_pldif_10g_rx_pld_rst_n	:	out	std_logic	:=	'0';
		int_pldif_10g_rx_prbs_err_clr	:	out	std_logic	:=	'0';
		int_pldif_10g_rx_rd_en	:	out	std_logic	:=	'0';
		int_pldif_8g_a1a2_size	:	out	std_logic	:=	'0';
		int_pldif_8g_bitloc_rev_en	:	out	std_logic	:=	'0';
		int_pldif_8g_bitslip	:	out	std_logic	:=	'0';
		int_pldif_8g_byte_rev_en	:	out	std_logic	:=	'0';
		int_pldif_8g_encdt	:	out	std_logic	:=	'0';
		int_pldif_8g_pld_rx_clk	:	out	std_logic	:=	'0';
		int_pldif_8g_rdenable_rx	:	out	std_logic	:=	'0';
		int_pldif_8g_rxpolarity	:	out	std_logic	:=	'0';
		int_pldif_8g_rxurstpcs_n	:	out	std_logic	:=	'0';
		int_pldif_8g_syncsm_en	:	out	std_logic	:=	'0';
		int_pldif_8g_wrdisable_rx	:	out	std_logic	:=	'0';
		int_pldif_g3_syncsm_en	:	out	std_logic	:=	'0';
		int_pldif_krfec_rx_clr_counters	:	out	std_logic	:=	'0';
		int_pldif_pmaif_polinv_rx	:	out	std_logic	:=	'0';
		int_pldif_pmaif_rx_clkslip	:	out	std_logic	:=	'0';
		int_pldif_pmaif_rx_pld_clk	:	out	std_logic	:=	'0';
		int_pldif_pmaif_rx_pld_rst_n	:	out	std_logic	:=	'0';
		int_pldif_pmaif_rx_prbs_err_clr	:	out	std_logic	:=	'0';
		int_pldif_pmaif_rxpma_rstb	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_blk_lock	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_diag_data_status	:	out	std_logic_vector(1 downto 0)	:=	"00";
		pld_10g_krfec_rx_frame	:	out	std_logic	:=	'0';
		pld_10g_rx_align_val	:	out	std_logic	:=	'0';
		pld_10g_rx_crc32_err	:	out	std_logic	:=	'0';
		pld_10g_rx_data_valid	:	out	std_logic	:=	'0';
		pld_10g_rx_empty	:	out	std_logic	:=	'0';
		pld_10g_rx_fifo_del	:	out	std_logic	:=	'0';
		pld_10g_rx_fifo_insert	:	out	std_logic	:=	'0';
		pld_10g_rx_fifo_num	:	out	std_logic_vector(4 downto 0)	:=	"00000";
		pld_10g_rx_frame_lock	:	out	std_logic	:=	'0';
		pld_10g_rx_hi_ber	:	out	std_logic	:=	'0';
		pld_10g_rx_oflw_err	:	out	std_logic	:=	'0';
		pld_10g_rx_pempty	:	out	std_logic	:=	'0';
		pld_10g_rx_pfull	:	out	std_logic	:=	'0';
		pld_8g_a1a2_k1k2_flag	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		pld_8g_empty_rmf	:	out	std_logic	:=	'0';
		pld_8g_empty_rx	:	out	std_logic	:=	'0';
		pld_8g_full_rmf	:	out	std_logic	:=	'0';
		pld_8g_full_rx	:	out	std_logic	:=	'0';
		pld_8g_rxelecidle	:	out	std_logic	:=	'0';
		pld_8g_signal_detect_out	:	out	std_logic	:=	'0';
		pld_8g_wa_boundary	:	out	std_logic_vector(4 downto 0)	:=	"00000";
		pld_pcs_rx_clk_out	:	out	std_logic	:=	'0';
		pld_pma_clkdiv_rx_user	:	out	std_logic	:=	'0';
		pld_pma_rx_clk_out	:	out	std_logic	:=	'0';
		pld_pma_signal_ok	:	out	std_logic	:=	'0';
		pld_rx_control	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		pld_rx_data	:	out	std_logic_vector(127 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		pld_rx_prbs_done	:	out	std_logic	:=	'0';
		pld_rx_prbs_err	:	out	std_logic	:=	'0'
	);
end twentynm_hssi_rx_pld_pcs_interface;

architecture behavior of twentynm_hssi_rx_pld_pcs_interface	is

constant hd_chnl_clklow_clk_hz_int	:	integer	:=	bin2int(hd_chnl_clklow_clk_hz);
constant hd_chnl_fref_clk_hz_int	:	integer	:=	bin2int(hd_chnl_fref_clk_hz);
constant hd_chnl_hclk_clk_hz_int	:	integer	:=	bin2int(hd_chnl_hclk_clk_hz);
constant hd_chnl_pcs_pair_ac_pwr_uw_per_mhz_int	:	integer	:=	bin2int(hd_chnl_pcs_pair_ac_pwr_uw_per_mhz);
constant hd_chnl_pcs_rx_ac_pwr_uw_per_mhz_int	:	integer	:=	bin2int(hd_chnl_pcs_rx_ac_pwr_uw_per_mhz);
constant hd_chnl_pld_8g_refclk_dig_nonatpg_mode_clk_hz_int	:	integer	:=	bin2int(hd_chnl_pld_8g_refclk_dig_nonatpg_mode_clk_hz);
constant hd_chnl_pld_pcs_refclk_dig_nonatpg_mode_clk_hz_int	:	integer	:=	bin2int(hd_chnl_pld_pcs_refclk_dig_nonatpg_mode_clk_hz);
constant hd_chnl_pld_rx_clk_hz_int	:	integer	:=	bin2int(hd_chnl_pld_rx_clk_hz);
constant hd_chnl_pma_rx_clk_hz_int	:	integer	:=	bin2int(hd_chnl_pma_rx_clk_hz);



component	twentynm_hssi_rx_pld_pcs_interface_encrypted
	generic (
		-- Architecture parameters
		hd_10g_advanced_user_mode_rx	:	string	:=	"disable";
		hd_10g_channel_operation_mode	:	string	:=	"tx_rx_pair_enabled";
		hd_10g_ctrl_plane_bonding_rx	:	string	:=	"individual_rx";
		hd_10g_fifo_mode_rx	:	string	:=	"fifo_rx";
		hd_10g_low_latency_en_rx	:	string	:=	"enable";
		hd_10g_lpbk_en	:	string	:=	"disable";
		hd_10g_pma_dw_rx	:	string	:=	"pma_64b_rx";
		hd_10g_prot_mode_rx	:	string	:=	"disabled_prot_mode_rx";
		hd_10g_shared_fifo_width_rx	:	string	:=	"single_rx";
		hd_10g_sup_mode	:	string	:=	"user_mode";
		hd_10g_test_bus_mode	:	string	:=	"tx";
		hd_8g_channel_operation_mode	:	string	:=	"tx_rx_pair_enabled";
		hd_8g_ctrl_plane_bonding_rx	:	string	:=	"individual_rx";
		hd_8g_fifo_mode_rx	:	string	:=	"fifo_rx";
		hd_8g_hip_mode	:	string	:=	"disable";
		hd_8g_lpbk_en	:	string	:=	"disable";
		hd_8g_pma_dw_rx	:	string	:=	"pma_8b_rx";
		hd_8g_prot_mode_rx	:	string	:=	"disabled_prot_mode_rx";
		hd_8g_sup_mode	:	string	:=	"user_mode";
		hd_chnl_channel_operation_mode	:	string	:=	"tx_rx_pair_enabled";
		hd_chnl_clklow_clk_hz	:	integer	:=	0;
		hd_chnl_ctrl_plane_bonding_rx	:	string	:=	"individual_rx";
		hd_chnl_fref_clk_hz	:	integer	:=	0;
		hd_chnl_frequency_rules_en	:	string	:=	"disable";
		hd_chnl_func_mode	:	string	:=	"disable";
		hd_chnl_hclk_clk_hz	:	integer	:=	0;
		hd_chnl_hip_en	:	string	:=	"disable";
		hd_chnl_hrdrstctl_en	:	string	:=	"disable";
		hd_chnl_low_latency_en_rx	:	string	:=	"disable";
		hd_chnl_lpbk_en	:	string	:=	"disable";
		hd_chnl_operating_voltage	:	string	:=	"standard";
		hd_chnl_pcs_ac_pwr_rules_en	:	string	:=	"disable";
		hd_chnl_pcs_pair_ac_pwr_uw_per_mhz	:	integer	:=	0;
		hd_chnl_pcs_rx_ac_pwr_uw_per_mhz	:	integer	:=	0;
		hd_chnl_pcs_rx_pwr_scaling_clk	:	string	:=	"pma_rx_clk";
		hd_chnl_pld_8g_refclk_dig_nonatpg_mode_clk_hz	:	integer	:=	0;
		hd_chnl_pld_fifo_mode_rx	:	string	:=	"fifo_rx";
		hd_chnl_pld_pcs_refclk_dig_nonatpg_mode_clk_hz	:	integer	:=	0;
		hd_chnl_pld_rx_clk_hz	:	integer	:=	0;
		hd_chnl_pma_dw_rx	:	string	:=	"pma_8b_rx";
		hd_chnl_pma_rx_clk_hz	:	integer	:=	0;
		hd_chnl_prot_mode_rx	:	string	:=	"disabled_prot_mode_rx";
		hd_chnl_shared_fifo_width_rx	:	string	:=	"single_rx";
		hd_chnl_speed_grade	:	string	:=	"e2";
		hd_chnl_sup_mode	:	string	:=	"user_mode";
		hd_chnl_transparent_pcs_rx	:	string	:=	"disable";
		hd_fifo_channel_operation_mode	:	string	:=	"tx_rx_pair_enabled";
		hd_fifo_prot_mode_rx	:	string	:=	"teng_mode_rx";
		hd_fifo_shared_fifo_width_rx	:	string	:=	"single_rx";
		hd_fifo_sup_mode	:	string	:=	"user_mode";
		hd_g3_prot_mode	:	string	:=	"disabled_prot_mode";
		hd_g3_sup_mode	:	string	:=	"user_mode";
		hd_krfec_channel_operation_mode	:	string	:=	"tx_rx_pair_enabled";
		hd_krfec_low_latency_en_rx	:	string	:=	"disable";
		hd_krfec_lpbk_en	:	string	:=	"disable";
		hd_krfec_prot_mode_rx	:	string	:=	"disabled_prot_mode_rx";
		hd_krfec_sup_mode	:	string	:=	"user_mode";
		hd_krfec_test_bus_mode	:	string	:=	"tx";
		hd_pldif_hrdrstctl_en	:	string	:=	"disable";
		hd_pldif_prot_mode_rx	:	string	:=	"disabled_prot_mode_rx";
		hd_pldif_sup_mode	:	string	:=	"user_mode";
		hd_pmaif_channel_operation_mode	:	string	:=	"tx_rx_pair_enabled";
		hd_pmaif_lpbk_en	:	string	:=	"disable";
		hd_pmaif_pma_dw_rx	:	string	:=	"pma_8b_rx";
		hd_pmaif_prot_mode_rx	:	string	:=	"disabled_prot_mode_rx";
		hd_pmaif_sim_mode	:	string	:=	"disable";
		hd_pmaif_sup_mode	:	string	:=	"user_mode";
		pcs_rx_block_sel	:	string	:=	"pcs_direct";
		pcs_rx_clk_out_sel	:	string	:=	"teng_clk_out";
		pcs_rx_clk_sel	:	string	:=	"pld_rx_clk";
		pcs_rx_hip_clk_en	:	string	:=	"hip_rx_enable";
		pcs_rx_output_sel	:	string	:=	"teng_output";
		reconfig_settings	:	string	:=	"{}";
		silicon_rev	:	string	:=	"20nm5es"
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		int_pldif_10g_rx_align_val	:	in	std_logic	:=	'0';
		int_pldif_10g_rx_blk_lock	:	in	std_logic	:=	'0';
		int_pldif_10g_rx_clk_out	:	in	std_logic	:=	'0';
		int_pldif_10g_rx_clk_out_pld_if	:	in	std_logic	:=	'0';
		int_pldif_10g_rx_control	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		int_pldif_10g_rx_crc32_err	:	in	std_logic	:=	'0';
		int_pldif_10g_rx_data	:	in	std_logic_vector(127 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		int_pldif_10g_rx_data_valid	:	in	std_logic	:=	'0';
		int_pldif_10g_rx_diag_status	:	in	std_logic_vector(1 downto 0)	:=	"00";
		int_pldif_10g_rx_empty	:	in	std_logic	:=	'0';
		int_pldif_10g_rx_fifo_del	:	in	std_logic	:=	'0';
		int_pldif_10g_rx_fifo_insert	:	in	std_logic	:=	'0';
		int_pldif_10g_rx_fifo_num	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		int_pldif_10g_rx_frame_lock	:	in	std_logic	:=	'0';
		int_pldif_10g_rx_hi_ber	:	in	std_logic	:=	'0';
		int_pldif_10g_rx_oflw_err	:	in	std_logic	:=	'0';
		int_pldif_10g_rx_pempty	:	in	std_logic	:=	'0';
		int_pldif_10g_rx_pfull	:	in	std_logic	:=	'0';
		int_pldif_10g_rx_rx_frame	:	in	std_logic	:=	'0';
		int_pldif_8g_a1a2_k1k2_flag	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		int_pldif_8g_empty_rmf	:	in	std_logic	:=	'0';
		int_pldif_8g_empty_rx	:	in	std_logic	:=	'0';
		int_pldif_8g_full_rmf	:	in	std_logic	:=	'0';
		int_pldif_8g_full_rx	:	in	std_logic	:=	'0';
		int_pldif_8g_phystatus	:	in	std_logic	:=	'0';
		int_pldif_8g_rx_blk_start	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		int_pldif_8g_rx_clk	:	in	std_logic	:=	'0';
		int_pldif_8g_rx_clk_out_pld_if	:	in	std_logic	:=	'0';
		int_pldif_8g_rx_data_valid	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		int_pldif_8g_rx_rstn_sync2wrfifo	:	in	std_logic	:=	'0';
		int_pldif_8g_rx_sync_hdr	:	in	std_logic_vector(1 downto 0)	:=	"00";
		int_pldif_8g_rxd	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		int_pldif_8g_rxelecidle	:	in	std_logic	:=	'0';
		int_pldif_8g_rxstatus	:	in	std_logic_vector(2 downto 0)	:=	"000";
		int_pldif_8g_rxvalid	:	in	std_logic	:=	'0';
		int_pldif_8g_signal_detect_out	:	in	std_logic	:=	'0';
		int_pldif_8g_wa_boundary	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		int_pldif_krfec_rx_block_lock	:	in	std_logic	:=	'0';
		int_pldif_krfec_rx_data_status	:	in	std_logic_vector(1 downto 0)	:=	"00";
		int_pldif_krfec_rx_frame	:	in	std_logic	:=	'0';
		int_pldif_pmaif_clkdiv_rx	:	in	std_logic	:=	'0';
		int_pldif_pmaif_clkdiv_rx_user	:	in	std_logic	:=	'0';
		int_pldif_pmaif_rx_data	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		int_pldif_pmaif_rx_prbs_done	:	in	std_logic	:=	'0';
		int_pldif_pmaif_rx_prbs_err	:	in	std_logic	:=	'0';
		int_pldif_pmaif_rxpll_lock	:	in	std_logic	:=	'0';
		int_pldif_pmaif_signal_ok	:	in	std_logic	:=	'0';
		int_pldif_usr_rst_sel	:	in	std_logic	:=	'0';
		pld_10g_krfec_rx_clr_errblk_cnt	:	in	std_logic	:=	'0';
		pld_10g_krfec_rx_pld_rst_n	:	in	std_logic	:=	'0';
		pld_10g_rx_align_clr	:	in	std_logic	:=	'0';
		pld_10g_rx_clr_ber_count	:	in	std_logic	:=	'0';
		pld_10g_rx_rd_en	:	in	std_logic	:=	'0';
		pld_8g_a1a2_size	:	in	std_logic	:=	'0';
		pld_8g_bitloc_rev_en	:	in	std_logic	:=	'0';
		pld_8g_byte_rev_en	:	in	std_logic	:=	'0';
		pld_8g_encdt	:	in	std_logic	:=	'0';
		pld_8g_g3_rx_pld_rst_n	:	in	std_logic	:=	'0';
		pld_8g_rdenable_rx	:	in	std_logic	:=	'0';
		pld_8g_rxpolarity	:	in	std_logic	:=	'0';
		pld_8g_wrdisable_rx	:	in	std_logic	:=	'0';
		pld_bitslip	:	in	std_logic	:=	'0';
		pld_partial_reconfig	:	in	std_logic	:=	'0';
		pld_pma_rxpma_rstb	:	in	std_logic	:=	'0';
		pld_pmaif_rx_pld_rst_n	:	in	std_logic	:=	'0';
		pld_pmaif_rxclkslip	:	in	std_logic	:=	'0';
		pld_polinv_rx	:	in	std_logic	:=	'0';
		pld_rx_clk	:	in	std_logic	:=	'0';
		pld_rx_prbs_err_clr	:	in	std_logic	:=	'0';
		pld_syncsm_en	:	in	std_logic	:=	'0';
		scan_mode_n	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		pld_8g_wa_boundary_txclk_fastreg	:	out	std_logic	:=	'0';
		pld_8g_wa_boundary_txclk_reg	:	out	std_logic	:=	'0';
		pld_bitslip_10g_txclk_reg	:	out	std_logic	:=	'0';
		pld_bitslip_8g_txclk_reg	:	out	std_logic	:=	'0';
		pld_bitslip_rxclk_parallel_loopback_reg	:	out	std_logic	:=	'0';
		pld_bitslip_rxclk_reg	:	out	std_logic	:=	'0';
		pld_pcs_rx_clk_out_pcsdirect_wire	:	out	std_logic	:=	'0';
		pld_pma_rx_clk_out_10g_or_pcsdirect_wire	:	out	std_logic	:=	'0';
		pld_pma_rx_clk_out_8g_wire	:	out	std_logic	:=	'0';
		pld_pmaif_rx_pld_rst_n_reg	:	out	std_logic	:=	'0';
		pld_pmaif_tx_pld_rst_n_txclk_reg	:	out	std_logic	:=	'0';
		pld_polinv_rx_reg	:	out	std_logic	:=	'0';
		pld_rx_clk_fifo	:	out	std_logic	:=	'0';
		pld_rx_control_fifo	:	out	std_logic	:=	'0';
		pld_rx_control_pcsdirect_reg	:	out	std_logic	:=	'0';
		pld_rx_data_fifo	:	out	std_logic	:=	'0';
		pld_rx_data_pcsdirect_reg	:	out	std_logic	:=	'0';
		pld_rx_prbs_done_reg	:	out	std_logic	:=	'0';
		pld_rx_prbs_done_txclk_reg	:	out	std_logic	:=	'0';
		pld_rx_prbs_err_clr_pcsdirect_txclk_reg	:	out	std_logic	:=	'0';
		pld_rx_prbs_err_clr_reg	:	out	std_logic	:=	'0';
		pld_rx_prbs_err_disprbs_reg	:	out	std_logic	:=	'0';
		pld_rx_prbs_err_pcsdirect_txclk_reg	:	out	std_logic	:=	'0';
		pld_rx_prbs_err_reg	:	out	std_logic	:=	'0';
		pma_rx_pma_clk_reg	:	out	std_logic	:=	'0';
		hip_rx_ctrl	:	out	std_logic_vector(1 downto 0)	:=	"00";
		hip_rx_data	:	out	std_logic_vector(50 downto 0)	:=	"000000000000000000000000000000000000000000000000000";
		int_pldif_10g_rx_align_clr	:	out	std_logic	:=	'0';
		int_pldif_10g_rx_bitslip	:	out	std_logic	:=	'0';
		int_pldif_10g_rx_clr_ber_count	:	out	std_logic	:=	'0';
		int_pldif_10g_rx_clr_errblk_cnt	:	out	std_logic	:=	'0';
		int_pldif_10g_rx_control_fb	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		int_pldif_10g_rx_data_fb	:	out	std_logic_vector(127 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		int_pldif_10g_rx_data_valid_fb	:	out	std_logic	:=	'0';
		int_pldif_10g_rx_pld_clk	:	out	std_logic	:=	'0';
		int_pldif_10g_rx_pld_rst_n	:	out	std_logic	:=	'0';
		int_pldif_10g_rx_prbs_err_clr	:	out	std_logic	:=	'0';
		int_pldif_10g_rx_rd_en	:	out	std_logic	:=	'0';
		int_pldif_8g_a1a2_size	:	out	std_logic	:=	'0';
		int_pldif_8g_bitloc_rev_en	:	out	std_logic	:=	'0';
		int_pldif_8g_bitslip	:	out	std_logic	:=	'0';
		int_pldif_8g_byte_rev_en	:	out	std_logic	:=	'0';
		int_pldif_8g_encdt	:	out	std_logic	:=	'0';
		int_pldif_8g_pld_rx_clk	:	out	std_logic	:=	'0';
		int_pldif_8g_rdenable_rx	:	out	std_logic	:=	'0';
		int_pldif_8g_rxpolarity	:	out	std_logic	:=	'0';
		int_pldif_8g_rxurstpcs_n	:	out	std_logic	:=	'0';
		int_pldif_8g_syncsm_en	:	out	std_logic	:=	'0';
		int_pldif_8g_wrdisable_rx	:	out	std_logic	:=	'0';
		int_pldif_g3_syncsm_en	:	out	std_logic	:=	'0';
		int_pldif_krfec_rx_clr_counters	:	out	std_logic	:=	'0';
		int_pldif_pmaif_polinv_rx	:	out	std_logic	:=	'0';
		int_pldif_pmaif_rx_clkslip	:	out	std_logic	:=	'0';
		int_pldif_pmaif_rx_pld_clk	:	out	std_logic	:=	'0';
		int_pldif_pmaif_rx_pld_rst_n	:	out	std_logic	:=	'0';
		int_pldif_pmaif_rx_prbs_err_clr	:	out	std_logic	:=	'0';
		int_pldif_pmaif_rxpma_rstb	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_blk_lock	:	out	std_logic	:=	'0';
		pld_10g_krfec_rx_diag_data_status	:	out	std_logic_vector(1 downto 0)	:=	"00";
		pld_10g_krfec_rx_frame	:	out	std_logic	:=	'0';
		pld_10g_rx_align_val	:	out	std_logic	:=	'0';
		pld_10g_rx_crc32_err	:	out	std_logic	:=	'0';
		pld_10g_rx_data_valid	:	out	std_logic	:=	'0';
		pld_10g_rx_empty	:	out	std_logic	:=	'0';
		pld_10g_rx_fifo_del	:	out	std_logic	:=	'0';
		pld_10g_rx_fifo_insert	:	out	std_logic	:=	'0';
		pld_10g_rx_fifo_num	:	out	std_logic_vector(4 downto 0)	:=	"00000";
		pld_10g_rx_frame_lock	:	out	std_logic	:=	'0';
		pld_10g_rx_hi_ber	:	out	std_logic	:=	'0';
		pld_10g_rx_oflw_err	:	out	std_logic	:=	'0';
		pld_10g_rx_pempty	:	out	std_logic	:=	'0';
		pld_10g_rx_pfull	:	out	std_logic	:=	'0';
		pld_8g_a1a2_k1k2_flag	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		pld_8g_empty_rmf	:	out	std_logic	:=	'0';
		pld_8g_empty_rx	:	out	std_logic	:=	'0';
		pld_8g_full_rmf	:	out	std_logic	:=	'0';
		pld_8g_full_rx	:	out	std_logic	:=	'0';
		pld_8g_rxelecidle	:	out	std_logic	:=	'0';
		pld_8g_signal_detect_out	:	out	std_logic	:=	'0';
		pld_8g_wa_boundary	:	out	std_logic_vector(4 downto 0)	:=	"00000";
		pld_pcs_rx_clk_out	:	out	std_logic	:=	'0';
		pld_pma_clkdiv_rx_user	:	out	std_logic	:=	'0';
		pld_pma_rx_clk_out	:	out	std_logic	:=	'0';
		pld_pma_signal_ok	:	out	std_logic	:=	'0';
		pld_rx_control	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		pld_rx_data	:	out	std_logic_vector(127 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		pld_rx_prbs_done	:	out	std_logic	:=	'0';
		pld_rx_prbs_err	:	out	std_logic	:=	'0'
	);
end component;

begin



inst : twentynm_hssi_rx_pld_pcs_interface_encrypted
	generic map (
		-- Instance parameters
		hd_10g_advanced_user_mode_rx	=>	hd_10g_advanced_user_mode_rx,
		hd_10g_channel_operation_mode	=>	hd_10g_channel_operation_mode,
		hd_10g_ctrl_plane_bonding_rx	=>	hd_10g_ctrl_plane_bonding_rx,
		hd_10g_fifo_mode_rx	=>	hd_10g_fifo_mode_rx,
		hd_10g_low_latency_en_rx	=>	hd_10g_low_latency_en_rx,
		hd_10g_lpbk_en	=>	hd_10g_lpbk_en,
		hd_10g_pma_dw_rx	=>	hd_10g_pma_dw_rx,
		hd_10g_prot_mode_rx	=>	hd_10g_prot_mode_rx,
		hd_10g_shared_fifo_width_rx	=>	hd_10g_shared_fifo_width_rx,
		hd_10g_sup_mode	=>	hd_10g_sup_mode,
		hd_10g_test_bus_mode	=>	hd_10g_test_bus_mode,
		hd_8g_channel_operation_mode	=>	hd_8g_channel_operation_mode,
		hd_8g_ctrl_plane_bonding_rx	=>	hd_8g_ctrl_plane_bonding_rx,
		hd_8g_fifo_mode_rx	=>	hd_8g_fifo_mode_rx,
		hd_8g_hip_mode	=>	hd_8g_hip_mode,
		hd_8g_lpbk_en	=>	hd_8g_lpbk_en,
		hd_8g_pma_dw_rx	=>	hd_8g_pma_dw_rx,
		hd_8g_prot_mode_rx	=>	hd_8g_prot_mode_rx,
		hd_8g_sup_mode	=>	hd_8g_sup_mode,
		hd_chnl_channel_operation_mode	=>	hd_chnl_channel_operation_mode,
		hd_chnl_clklow_clk_hz	=>	hd_chnl_clklow_clk_hz_int,
		hd_chnl_ctrl_plane_bonding_rx	=>	hd_chnl_ctrl_plane_bonding_rx,
		hd_chnl_fref_clk_hz	=>	hd_chnl_fref_clk_hz_int,
		hd_chnl_frequency_rules_en	=>	hd_chnl_frequency_rules_en,
		hd_chnl_func_mode	=>	hd_chnl_func_mode,
		hd_chnl_hclk_clk_hz	=>	hd_chnl_hclk_clk_hz_int,
		hd_chnl_hip_en	=>	hd_chnl_hip_en,
		hd_chnl_hrdrstctl_en	=>	hd_chnl_hrdrstctl_en,
		hd_chnl_low_latency_en_rx	=>	hd_chnl_low_latency_en_rx,
		hd_chnl_lpbk_en	=>	hd_chnl_lpbk_en,
		hd_chnl_operating_voltage	=>	hd_chnl_operating_voltage,
		hd_chnl_pcs_ac_pwr_rules_en	=>	hd_chnl_pcs_ac_pwr_rules_en,
		hd_chnl_pcs_pair_ac_pwr_uw_per_mhz	=>	hd_chnl_pcs_pair_ac_pwr_uw_per_mhz_int,
		hd_chnl_pcs_rx_ac_pwr_uw_per_mhz	=>	hd_chnl_pcs_rx_ac_pwr_uw_per_mhz_int,
		hd_chnl_pcs_rx_pwr_scaling_clk	=>	hd_chnl_pcs_rx_pwr_scaling_clk,
		hd_chnl_pld_8g_refclk_dig_nonatpg_mode_clk_hz	=>	hd_chnl_pld_8g_refclk_dig_nonatpg_mode_clk_hz_int,
		hd_chnl_pld_fifo_mode_rx	=>	hd_chnl_pld_fifo_mode_rx,
		hd_chnl_pld_pcs_refclk_dig_nonatpg_mode_clk_hz	=>	hd_chnl_pld_pcs_refclk_dig_nonatpg_mode_clk_hz_int,
		hd_chnl_pld_rx_clk_hz	=>	hd_chnl_pld_rx_clk_hz_int,
		hd_chnl_pma_dw_rx	=>	hd_chnl_pma_dw_rx,
		hd_chnl_pma_rx_clk_hz	=>	hd_chnl_pma_rx_clk_hz_int,
		hd_chnl_prot_mode_rx	=>	hd_chnl_prot_mode_rx,
		hd_chnl_shared_fifo_width_rx	=>	hd_chnl_shared_fifo_width_rx,
		hd_chnl_speed_grade	=>	hd_chnl_speed_grade,
		hd_chnl_sup_mode	=>	hd_chnl_sup_mode,
		hd_chnl_transparent_pcs_rx	=>	hd_chnl_transparent_pcs_rx,
		hd_fifo_channel_operation_mode	=>	hd_fifo_channel_operation_mode,
		hd_fifo_prot_mode_rx	=>	hd_fifo_prot_mode_rx,
		hd_fifo_shared_fifo_width_rx	=>	hd_fifo_shared_fifo_width_rx,
		hd_fifo_sup_mode	=>	hd_fifo_sup_mode,
		hd_g3_prot_mode	=>	hd_g3_prot_mode,
		hd_g3_sup_mode	=>	hd_g3_sup_mode,
		hd_krfec_channel_operation_mode	=>	hd_krfec_channel_operation_mode,
		hd_krfec_low_latency_en_rx	=>	hd_krfec_low_latency_en_rx,
		hd_krfec_lpbk_en	=>	hd_krfec_lpbk_en,
		hd_krfec_prot_mode_rx	=>	hd_krfec_prot_mode_rx,
		hd_krfec_sup_mode	=>	hd_krfec_sup_mode,
		hd_krfec_test_bus_mode	=>	hd_krfec_test_bus_mode,
		hd_pldif_hrdrstctl_en	=>	hd_pldif_hrdrstctl_en,
		hd_pldif_prot_mode_rx	=>	hd_pldif_prot_mode_rx,
		hd_pldif_sup_mode	=>	hd_pldif_sup_mode,
		hd_pmaif_channel_operation_mode	=>	hd_pmaif_channel_operation_mode,
		hd_pmaif_lpbk_en	=>	hd_pmaif_lpbk_en,
		hd_pmaif_pma_dw_rx	=>	hd_pmaif_pma_dw_rx,
		hd_pmaif_prot_mode_rx	=>	hd_pmaif_prot_mode_rx,
		hd_pmaif_sim_mode	=>	hd_pmaif_sim_mode,
		hd_pmaif_sup_mode	=>	hd_pmaif_sup_mode,
		pcs_rx_block_sel	=>	pcs_rx_block_sel,
		pcs_rx_clk_out_sel	=>	pcs_rx_clk_out_sel,
		pcs_rx_clk_sel	=>	pcs_rx_clk_sel,
		pcs_rx_hip_clk_en	=>	pcs_rx_hip_clk_en,
		pcs_rx_output_sel	=>	pcs_rx_output_sel,
		reconfig_settings	=>	reconfig_settings,
		silicon_rev	=>	silicon_rev
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		int_pldif_10g_rx_align_val	=>	int_pldif_10g_rx_align_val,
		int_pldif_10g_rx_blk_lock	=>	int_pldif_10g_rx_blk_lock,
		int_pldif_10g_rx_clk_out	=>	int_pldif_10g_rx_clk_out,
		int_pldif_10g_rx_clk_out_pld_if	=>	int_pldif_10g_rx_clk_out_pld_if,
		int_pldif_10g_rx_control	=>	int_pldif_10g_rx_control,
		int_pldif_10g_rx_crc32_err	=>	int_pldif_10g_rx_crc32_err,
		int_pldif_10g_rx_data	=>	int_pldif_10g_rx_data,
		int_pldif_10g_rx_data_valid	=>	int_pldif_10g_rx_data_valid,
		int_pldif_10g_rx_diag_status	=>	int_pldif_10g_rx_diag_status,
		int_pldif_10g_rx_empty	=>	int_pldif_10g_rx_empty,
		int_pldif_10g_rx_fifo_del	=>	int_pldif_10g_rx_fifo_del,
		int_pldif_10g_rx_fifo_insert	=>	int_pldif_10g_rx_fifo_insert,
		int_pldif_10g_rx_fifo_num	=>	int_pldif_10g_rx_fifo_num,
		int_pldif_10g_rx_frame_lock	=>	int_pldif_10g_rx_frame_lock,
		int_pldif_10g_rx_hi_ber	=>	int_pldif_10g_rx_hi_ber,
		int_pldif_10g_rx_oflw_err	=>	int_pldif_10g_rx_oflw_err,
		int_pldif_10g_rx_pempty	=>	int_pldif_10g_rx_pempty,
		int_pldif_10g_rx_pfull	=>	int_pldif_10g_rx_pfull,
		int_pldif_10g_rx_rx_frame	=>	int_pldif_10g_rx_rx_frame,
		int_pldif_8g_a1a2_k1k2_flag	=>	int_pldif_8g_a1a2_k1k2_flag,
		int_pldif_8g_empty_rmf	=>	int_pldif_8g_empty_rmf,
		int_pldif_8g_empty_rx	=>	int_pldif_8g_empty_rx,
		int_pldif_8g_full_rmf	=>	int_pldif_8g_full_rmf,
		int_pldif_8g_full_rx	=>	int_pldif_8g_full_rx,
		int_pldif_8g_phystatus	=>	int_pldif_8g_phystatus,
		int_pldif_8g_rx_blk_start	=>	int_pldif_8g_rx_blk_start,
		int_pldif_8g_rx_clk	=>	int_pldif_8g_rx_clk,
		int_pldif_8g_rx_clk_out_pld_if	=>	int_pldif_8g_rx_clk_out_pld_if,
		int_pldif_8g_rx_data_valid	=>	int_pldif_8g_rx_data_valid,
		int_pldif_8g_rx_rstn_sync2wrfifo	=>	int_pldif_8g_rx_rstn_sync2wrfifo,
		int_pldif_8g_rx_sync_hdr	=>	int_pldif_8g_rx_sync_hdr,
		int_pldif_8g_rxd	=>	int_pldif_8g_rxd,
		int_pldif_8g_rxelecidle	=>	int_pldif_8g_rxelecidle,
		int_pldif_8g_rxstatus	=>	int_pldif_8g_rxstatus,
		int_pldif_8g_rxvalid	=>	int_pldif_8g_rxvalid,
		int_pldif_8g_signal_detect_out	=>	int_pldif_8g_signal_detect_out,
		int_pldif_8g_wa_boundary	=>	int_pldif_8g_wa_boundary,
		int_pldif_krfec_rx_block_lock	=>	int_pldif_krfec_rx_block_lock,
		int_pldif_krfec_rx_data_status	=>	int_pldif_krfec_rx_data_status,
		int_pldif_krfec_rx_frame	=>	int_pldif_krfec_rx_frame,
		int_pldif_pmaif_clkdiv_rx	=>	int_pldif_pmaif_clkdiv_rx,
		int_pldif_pmaif_clkdiv_rx_user	=>	int_pldif_pmaif_clkdiv_rx_user,
		int_pldif_pmaif_rx_data	=>	int_pldif_pmaif_rx_data,
		int_pldif_pmaif_rx_prbs_done	=>	int_pldif_pmaif_rx_prbs_done,
		int_pldif_pmaif_rx_prbs_err	=>	int_pldif_pmaif_rx_prbs_err,
		int_pldif_pmaif_rxpll_lock	=>	int_pldif_pmaif_rxpll_lock,
		int_pldif_pmaif_signal_ok	=>	int_pldif_pmaif_signal_ok,
		int_pldif_usr_rst_sel	=>	int_pldif_usr_rst_sel,
		pld_10g_krfec_rx_clr_errblk_cnt	=>	pld_10g_krfec_rx_clr_errblk_cnt,
		pld_10g_krfec_rx_pld_rst_n	=>	pld_10g_krfec_rx_pld_rst_n,
		pld_10g_rx_align_clr	=>	pld_10g_rx_align_clr,
		pld_10g_rx_clr_ber_count	=>	pld_10g_rx_clr_ber_count,
		pld_10g_rx_rd_en	=>	pld_10g_rx_rd_en,
		pld_8g_a1a2_size	=>	pld_8g_a1a2_size,
		pld_8g_bitloc_rev_en	=>	pld_8g_bitloc_rev_en,
		pld_8g_byte_rev_en	=>	pld_8g_byte_rev_en,
		pld_8g_encdt	=>	pld_8g_encdt,
		pld_8g_g3_rx_pld_rst_n	=>	pld_8g_g3_rx_pld_rst_n,
		pld_8g_rdenable_rx	=>	pld_8g_rdenable_rx,
		pld_8g_rxpolarity	=>	pld_8g_rxpolarity,
		pld_8g_wrdisable_rx	=>	pld_8g_wrdisable_rx,
		pld_bitslip	=>	pld_bitslip,
		pld_partial_reconfig	=>	pld_partial_reconfig,
		pld_pma_rxpma_rstb	=>	pld_pma_rxpma_rstb,
		pld_pmaif_rx_pld_rst_n	=>	pld_pmaif_rx_pld_rst_n,
		pld_pmaif_rxclkslip	=>	pld_pmaif_rxclkslip,
		pld_polinv_rx	=>	pld_polinv_rx,
		pld_rx_clk	=>	pld_rx_clk,
		pld_rx_prbs_err_clr	=>	pld_rx_prbs_err_clr,
		pld_syncsm_en	=>	pld_syncsm_en,
		scan_mode_n	=>	scan_mode_n,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		pld_8g_wa_boundary_txclk_fastreg	=>	pld_8g_wa_boundary_txclk_fastreg,
		pld_8g_wa_boundary_txclk_reg	=>	pld_8g_wa_boundary_txclk_reg,
		pld_bitslip_10g_txclk_reg	=>	pld_bitslip_10g_txclk_reg,
		pld_bitslip_8g_txclk_reg	=>	pld_bitslip_8g_txclk_reg,
		pld_bitslip_rxclk_parallel_loopback_reg	=>	pld_bitslip_rxclk_parallel_loopback_reg,
		pld_bitslip_rxclk_reg	=>	pld_bitslip_rxclk_reg,
		pld_pcs_rx_clk_out_pcsdirect_wire	=>	pld_pcs_rx_clk_out_pcsdirect_wire,
		pld_pma_rx_clk_out_10g_or_pcsdirect_wire	=>	pld_pma_rx_clk_out_10g_or_pcsdirect_wire,
		pld_pma_rx_clk_out_8g_wire	=>	pld_pma_rx_clk_out_8g_wire,
		pld_pmaif_rx_pld_rst_n_reg	=>	pld_pmaif_rx_pld_rst_n_reg,
		pld_pmaif_tx_pld_rst_n_txclk_reg	=>	pld_pmaif_tx_pld_rst_n_txclk_reg,
		pld_polinv_rx_reg	=>	pld_polinv_rx_reg,
		pld_rx_clk_fifo	=>	pld_rx_clk_fifo,
		pld_rx_control_fifo	=>	pld_rx_control_fifo,
		pld_rx_control_pcsdirect_reg	=>	pld_rx_control_pcsdirect_reg,
		pld_rx_data_fifo	=>	pld_rx_data_fifo,
		pld_rx_data_pcsdirect_reg	=>	pld_rx_data_pcsdirect_reg,
		pld_rx_prbs_done_reg	=>	pld_rx_prbs_done_reg,
		pld_rx_prbs_done_txclk_reg	=>	pld_rx_prbs_done_txclk_reg,
		pld_rx_prbs_err_clr_pcsdirect_txclk_reg	=>	pld_rx_prbs_err_clr_pcsdirect_txclk_reg,
		pld_rx_prbs_err_clr_reg	=>	pld_rx_prbs_err_clr_reg,
		pld_rx_prbs_err_disprbs_reg	=>	pld_rx_prbs_err_disprbs_reg,
		pld_rx_prbs_err_pcsdirect_txclk_reg	=>	pld_rx_prbs_err_pcsdirect_txclk_reg,
		pld_rx_prbs_err_reg	=>	pld_rx_prbs_err_reg,
		pma_rx_pma_clk_reg	=>	pma_rx_pma_clk_reg,
		hip_rx_ctrl	=>	hip_rx_ctrl,
		hip_rx_data	=>	hip_rx_data,
		int_pldif_10g_rx_align_clr	=>	int_pldif_10g_rx_align_clr,
		int_pldif_10g_rx_bitslip	=>	int_pldif_10g_rx_bitslip,
		int_pldif_10g_rx_clr_ber_count	=>	int_pldif_10g_rx_clr_ber_count,
		int_pldif_10g_rx_clr_errblk_cnt	=>	int_pldif_10g_rx_clr_errblk_cnt,
		int_pldif_10g_rx_control_fb	=>	int_pldif_10g_rx_control_fb,
		int_pldif_10g_rx_data_fb	=>	int_pldif_10g_rx_data_fb,
		int_pldif_10g_rx_data_valid_fb	=>	int_pldif_10g_rx_data_valid_fb,
		int_pldif_10g_rx_pld_clk	=>	int_pldif_10g_rx_pld_clk,
		int_pldif_10g_rx_pld_rst_n	=>	int_pldif_10g_rx_pld_rst_n,
		int_pldif_10g_rx_prbs_err_clr	=>	int_pldif_10g_rx_prbs_err_clr,
		int_pldif_10g_rx_rd_en	=>	int_pldif_10g_rx_rd_en,
		int_pldif_8g_a1a2_size	=>	int_pldif_8g_a1a2_size,
		int_pldif_8g_bitloc_rev_en	=>	int_pldif_8g_bitloc_rev_en,
		int_pldif_8g_bitslip	=>	int_pldif_8g_bitslip,
		int_pldif_8g_byte_rev_en	=>	int_pldif_8g_byte_rev_en,
		int_pldif_8g_encdt	=>	int_pldif_8g_encdt,
		int_pldif_8g_pld_rx_clk	=>	int_pldif_8g_pld_rx_clk,
		int_pldif_8g_rdenable_rx	=>	int_pldif_8g_rdenable_rx,
		int_pldif_8g_rxpolarity	=>	int_pldif_8g_rxpolarity,
		int_pldif_8g_rxurstpcs_n	=>	int_pldif_8g_rxurstpcs_n,
		int_pldif_8g_syncsm_en	=>	int_pldif_8g_syncsm_en,
		int_pldif_8g_wrdisable_rx	=>	int_pldif_8g_wrdisable_rx,
		int_pldif_g3_syncsm_en	=>	int_pldif_g3_syncsm_en,
		int_pldif_krfec_rx_clr_counters	=>	int_pldif_krfec_rx_clr_counters,
		int_pldif_pmaif_polinv_rx	=>	int_pldif_pmaif_polinv_rx,
		int_pldif_pmaif_rx_clkslip	=>	int_pldif_pmaif_rx_clkslip,
		int_pldif_pmaif_rx_pld_clk	=>	int_pldif_pmaif_rx_pld_clk,
		int_pldif_pmaif_rx_pld_rst_n	=>	int_pldif_pmaif_rx_pld_rst_n,
		int_pldif_pmaif_rx_prbs_err_clr	=>	int_pldif_pmaif_rx_prbs_err_clr,
		int_pldif_pmaif_rxpma_rstb	=>	int_pldif_pmaif_rxpma_rstb,
		pld_10g_krfec_rx_blk_lock	=>	pld_10g_krfec_rx_blk_lock,
		pld_10g_krfec_rx_diag_data_status	=>	pld_10g_krfec_rx_diag_data_status,
		pld_10g_krfec_rx_frame	=>	pld_10g_krfec_rx_frame,
		pld_10g_rx_align_val	=>	pld_10g_rx_align_val,
		pld_10g_rx_crc32_err	=>	pld_10g_rx_crc32_err,
		pld_10g_rx_data_valid	=>	pld_10g_rx_data_valid,
		pld_10g_rx_empty	=>	pld_10g_rx_empty,
		pld_10g_rx_fifo_del	=>	pld_10g_rx_fifo_del,
		pld_10g_rx_fifo_insert	=>	pld_10g_rx_fifo_insert,
		pld_10g_rx_fifo_num	=>	pld_10g_rx_fifo_num,
		pld_10g_rx_frame_lock	=>	pld_10g_rx_frame_lock,
		pld_10g_rx_hi_ber	=>	pld_10g_rx_hi_ber,
		pld_10g_rx_oflw_err	=>	pld_10g_rx_oflw_err,
		pld_10g_rx_pempty	=>	pld_10g_rx_pempty,
		pld_10g_rx_pfull	=>	pld_10g_rx_pfull,
		pld_8g_a1a2_k1k2_flag	=>	pld_8g_a1a2_k1k2_flag,
		pld_8g_empty_rmf	=>	pld_8g_empty_rmf,
		pld_8g_empty_rx	=>	pld_8g_empty_rx,
		pld_8g_full_rmf	=>	pld_8g_full_rmf,
		pld_8g_full_rx	=>	pld_8g_full_rx,
		pld_8g_rxelecidle	=>	pld_8g_rxelecidle,
		pld_8g_signal_detect_out	=>	pld_8g_signal_detect_out,
		pld_8g_wa_boundary	=>	pld_8g_wa_boundary,
		pld_pcs_rx_clk_out	=>	pld_pcs_rx_clk_out,
		pld_pma_clkdiv_rx_user	=>	pld_pma_clkdiv_rx_user,
		pld_pma_rx_clk_out	=>	pld_pma_rx_clk_out,
		pld_pma_signal_ok	=>	pld_pma_signal_ok,
		pld_rx_control	=>	pld_rx_control,
		pld_rx_data	=>	pld_rx_data,
		pld_rx_prbs_done	=>	pld_rx_prbs_done,
		pld_rx_prbs_err	=>	pld_rx_prbs_err
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_tx_pcs_pma_interface	is
	generic (
		-- Entity parameters
		bypass_pma_txelecidle	:	string	:=	"false";
		channel_operation_mode	:	string	:=	"tx_rx_pair_enabled";
		lpbk_en	:	string	:=	"disable";
		master_clk_sel	:	string	:=	"master_tx_pma_clk";
		pcie_sub_prot_mode_tx	:	string	:=	"other_prot_mode";
		pldif_datawidth_mode	:	string	:=	"pldif_data_10bit";
		pma_dw_tx	:	string	:=	"pma_8b_tx";
		pma_if_dft_en	:	string	:=	"dft_dis";
		pmagate_en	:	string	:=	"pmagate_dis";
		prbs9_dwidth	:	string	:=	"prbs9_64b";
		prbs_clken	:	string	:=	"prbs_clk_dis";
		prbs_gen_pat	:	string	:=	"prbs_gen_dis";
		prot_mode_tx	:	string	:=	"disabled_prot_mode_tx";
		reconfig_settings	:	string	:=	"{}";
		silicon_rev	:	string	:=	"20nm5es";
		sq_wave_num	:	string	:=	"sq_wave_4";
		sqwgen_clken	:	string	:=	"sqwgen_clk_dis";
		sup_mode	:	string	:=	"user_mode";
		tx_dyn_polarity_inversion	:	string	:=	"tx_dyn_polinv_dis";
		tx_pma_data_sel	:	string	:=	"pld_dir";
		tx_static_polarity_inversion	:	string	:=	"tx_stat_polinv_dis";
		uhsif_cnt_step_filt_before_lock	:	string	:=	"uhsif_filt_stepsz_b4lock_4";
		uhsif_cnt_thresh_filt_after_lock_value	:	bit_vector	:=	B"1011";
		uhsif_cnt_thresh_filt_before_lock	:	string	:=	"uhsif_filt_cntthr_b4lock_16";
		uhsif_dcn_test_update_period	:	string	:=	"uhsif_dcn_test_period_4";
		uhsif_dcn_testmode_enable	:	string	:=	"uhsif_dcn_test_mode_disable";
		uhsif_dead_zone_count_thresh	:	string	:=	"uhsif_dzt_cnt_thr_4";
		uhsif_dead_zone_detection_enable	:	string	:=	"uhsif_dzt_enable";
		uhsif_dead_zone_obser_window	:	string	:=	"uhsif_dzt_obr_win_32";
		uhsif_dead_zone_skip_size	:	string	:=	"uhsif_dzt_skipsz_8";
		uhsif_delay_cell_index_sel	:	string	:=	"uhsif_index_internal";
		uhsif_delay_cell_margin	:	string	:=	"uhsif_dcn_margin_4";
		uhsif_delay_cell_static_index_value	:	bit_vector	:=	B"10000000";
		uhsif_dft_dead_zone_control	:	string	:=	"uhsif_dft_dz_det_val_0";
		uhsif_dft_up_filt_control	:	string	:=	"uhsif_dft_up_val_0";
		uhsif_enable	:	string	:=	"uhsif_disable";
		uhsif_lock_det_segsz_after_lock	:	string	:=	"uhsif_lkd_segsz_aflock_2048";
		uhsif_lock_det_segsz_before_lock	:	string	:=	"uhsif_lkd_segsz_b4lock_32";
		uhsif_lock_det_thresh_cnt_after_lock_value	:	bit_vector	:=	B"1000";
		uhsif_lock_det_thresh_cnt_before_lock_value	:	bit_vector	:=	B"1000";
		uhsif_lock_det_thresh_diff_after_lock_value	:	bit_vector	:=	B"0011";
		uhsif_lock_det_thresh_diff_before_lock_value	:	bit_vector	:=	B"0011"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		int_pmaif_10g_tx_clk_out	:	in	std_logic	:=	'0';
		int_pmaif_10g_tx_pma_data	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		int_pmaif_10g_tx_pma_data_gate_val	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		int_pmaif_8g_pudr	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		int_pmaif_8g_tx_clk_out	:	in	std_logic	:=	'0';
		int_pmaif_8g_tx_elec_idle	:	in	std_logic	:=	'0';
		int_pmaif_g3_data_sel	:	in	std_logic	:=	'0';
		int_pmaif_g3_pma_data_out	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		int_pmaif_g3_pma_tx_elec_idle	:	in	std_logic	:=	'0';
		int_pmaif_pldif_pmaif_tx_pld_rst_n	:	in	std_logic	:=	'0';
		int_pmaif_pldif_polinv_tx	:	in	std_logic	:=	'0';
		int_pmaif_pldif_tx_data	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		int_pmaif_pldif_txelecidle	:	in	std_logic	:=	'0';
		int_pmaif_pldif_txpma_rstb	:	in	std_logic	:=	'0';
		int_pmaif_pldif_uhsif_scan_chain_in	:	in	std_logic	:=	'0';
		int_pmaif_pldif_uhsif_tx_clk	:	in	std_logic	:=	'0';
		int_pmaif_pldif_uhsif_tx_data	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		pma_tx_clkdiv_user	:	in	std_logic	:=	'0';
		pma_tx_pma_clk	:	in	std_logic	:=	'0';
		refclk_dig	:	in	std_logic	:=	'0';
		refclk_dig_uhsif	:	in	std_logic	:=	'0';
		scan_mode_n	:	in	std_logic	:=	'0';
		uhsif_scan_mode_n	:	in	std_logic	:=	'0';
		uhsif_scan_shift_n	:	in	std_logic	:=	'0';
		write_en	:	in	std_logic_vector(1 downto 0)	:=	"00";
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		avmm_user_dataout	:	out	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		int_pmaif_10g_tx_pma_clk	:	out	std_logic	:=	'0';
		int_pmaif_8g_txpma_local_clk	:	out	std_logic	:=	'0';
		int_pmaif_pldif_tx_clkdiv	:	out	std_logic	:=	'0';
		int_pmaif_pldif_tx_clkdiv_user	:	out	std_logic	:=	'0';
		int_pmaif_pldif_uhsif_lock	:	out	std_logic	:=	'0';
		int_pmaif_pldif_uhsif_scan_chain_out	:	out	std_logic	:=	'0';
		int_pmaif_pldif_uhsif_tx_clk_out	:	out	std_logic	:=	'0';
		int_tx_dft_obsrv_clk	:	out	std_logic_vector(4 downto 0)	:=	"00000";
		pma_tx_elec_idle	:	out	std_logic	:=	'0';
		pma_tx_pma_data	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		pma_txpma_rstb	:	out	std_logic	:=	'0';
		tx_pma_data_loopback	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		tx_pma_uhsif_data_loopback	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		tx_prbs_gen_test	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		uhsif_test_out_1	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		uhsif_test_out_2	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		uhsif_test_out_3	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		write_en_ack	:	out	std_logic_vector(1 downto 0)	:=	"00"
	);
end twentynm_hssi_tx_pcs_pma_interface;

architecture behavior of twentynm_hssi_tx_pcs_pma_interface	is

constant uhsif_cnt_thresh_filt_after_lock_value_int	:	integer	:=	bin2int(uhsif_cnt_thresh_filt_after_lock_value);
constant uhsif_delay_cell_static_index_value_int	:	integer	:=	bin2int(uhsif_delay_cell_static_index_value);
constant uhsif_lock_det_thresh_cnt_after_lock_value_int	:	integer	:=	bin2int(uhsif_lock_det_thresh_cnt_after_lock_value);
constant uhsif_lock_det_thresh_cnt_before_lock_value_int	:	integer	:=	bin2int(uhsif_lock_det_thresh_cnt_before_lock_value);
constant uhsif_lock_det_thresh_diff_after_lock_value_int	:	integer	:=	bin2int(uhsif_lock_det_thresh_diff_after_lock_value);
constant uhsif_lock_det_thresh_diff_before_lock_value_int	:	integer	:=	bin2int(uhsif_lock_det_thresh_diff_before_lock_value);



component	twentynm_hssi_tx_pcs_pma_interface_encrypted
	generic (
		-- Architecture parameters
		bypass_pma_txelecidle	:	string	:=	"false";
		channel_operation_mode	:	string	:=	"tx_rx_pair_enabled";
		lpbk_en	:	string	:=	"disable";
		master_clk_sel	:	string	:=	"master_tx_pma_clk";
		pcie_sub_prot_mode_tx	:	string	:=	"other_prot_mode";
		pldif_datawidth_mode	:	string	:=	"pldif_data_10bit";
		pma_dw_tx	:	string	:=	"pma_8b_tx";
		pma_if_dft_en	:	string	:=	"dft_dis";
		pmagate_en	:	string	:=	"pmagate_dis";
		prbs9_dwidth	:	string	:=	"prbs9_64b";
		prbs_clken	:	string	:=	"prbs_clk_dis";
		prbs_gen_pat	:	string	:=	"prbs_gen_dis";
		prot_mode_tx	:	string	:=	"disabled_prot_mode_tx";
		reconfig_settings	:	string	:=	"{}";
		silicon_rev	:	string	:=	"20nm5es";
		sq_wave_num	:	string	:=	"sq_wave_4";
		sqwgen_clken	:	string	:=	"sqwgen_clk_dis";
		sup_mode	:	string	:=	"user_mode";
		tx_dyn_polarity_inversion	:	string	:=	"tx_dyn_polinv_dis";
		tx_pma_data_sel	:	string	:=	"pld_dir";
		tx_static_polarity_inversion	:	string	:=	"tx_stat_polinv_dis";
		uhsif_cnt_step_filt_before_lock	:	string	:=	"uhsif_filt_stepsz_b4lock_4";
		uhsif_cnt_thresh_filt_after_lock_value	:	integer	:=	11;
		uhsif_cnt_thresh_filt_before_lock	:	string	:=	"uhsif_filt_cntthr_b4lock_16";
		uhsif_dcn_test_update_period	:	string	:=	"uhsif_dcn_test_period_4";
		uhsif_dcn_testmode_enable	:	string	:=	"uhsif_dcn_test_mode_disable";
		uhsif_dead_zone_count_thresh	:	string	:=	"uhsif_dzt_cnt_thr_4";
		uhsif_dead_zone_detection_enable	:	string	:=	"uhsif_dzt_enable";
		uhsif_dead_zone_obser_window	:	string	:=	"uhsif_dzt_obr_win_32";
		uhsif_dead_zone_skip_size	:	string	:=	"uhsif_dzt_skipsz_8";
		uhsif_delay_cell_index_sel	:	string	:=	"uhsif_index_internal";
		uhsif_delay_cell_margin	:	string	:=	"uhsif_dcn_margin_4";
		uhsif_delay_cell_static_index_value	:	integer	:=	128;
		uhsif_dft_dead_zone_control	:	string	:=	"uhsif_dft_dz_det_val_0";
		uhsif_dft_up_filt_control	:	string	:=	"uhsif_dft_up_val_0";
		uhsif_enable	:	string	:=	"uhsif_disable";
		uhsif_lock_det_segsz_after_lock	:	string	:=	"uhsif_lkd_segsz_aflock_2048";
		uhsif_lock_det_segsz_before_lock	:	string	:=	"uhsif_lkd_segsz_b4lock_32";
		uhsif_lock_det_thresh_cnt_after_lock_value	:	integer	:=	8;
		uhsif_lock_det_thresh_cnt_before_lock_value	:	integer	:=	8;
		uhsif_lock_det_thresh_diff_after_lock_value	:	integer	:=	3;
		uhsif_lock_det_thresh_diff_before_lock_value	:	integer	:=	3
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		int_pmaif_10g_tx_clk_out	:	in	std_logic	:=	'0';
		int_pmaif_10g_tx_pma_data	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		int_pmaif_10g_tx_pma_data_gate_val	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		int_pmaif_8g_pudr	:	in	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		int_pmaif_8g_tx_clk_out	:	in	std_logic	:=	'0';
		int_pmaif_8g_tx_elec_idle	:	in	std_logic	:=	'0';
		int_pmaif_g3_data_sel	:	in	std_logic	:=	'0';
		int_pmaif_g3_pma_data_out	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		int_pmaif_g3_pma_tx_elec_idle	:	in	std_logic	:=	'0';
		int_pmaif_pldif_pmaif_tx_pld_rst_n	:	in	std_logic	:=	'0';
		int_pmaif_pldif_polinv_tx	:	in	std_logic	:=	'0';
		int_pmaif_pldif_tx_data	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		int_pmaif_pldif_txelecidle	:	in	std_logic	:=	'0';
		int_pmaif_pldif_txpma_rstb	:	in	std_logic	:=	'0';
		int_pmaif_pldif_uhsif_scan_chain_in	:	in	std_logic	:=	'0';
		int_pmaif_pldif_uhsif_tx_clk	:	in	std_logic	:=	'0';
		int_pmaif_pldif_uhsif_tx_data	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		pma_tx_clkdiv_user	:	in	std_logic	:=	'0';
		pma_tx_pma_clk	:	in	std_logic	:=	'0';
		refclk_dig	:	in	std_logic	:=	'0';
		refclk_dig_uhsif	:	in	std_logic	:=	'0';
		scan_mode_n	:	in	std_logic	:=	'0';
		uhsif_scan_mode_n	:	in	std_logic	:=	'0';
		uhsif_scan_shift_n	:	in	std_logic	:=	'0';
		write_en	:	in	std_logic_vector(1 downto 0)	:=	"00";
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		avmm_user_dataout	:	out	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		int_pmaif_10g_tx_pma_clk	:	out	std_logic	:=	'0';
		int_pmaif_8g_txpma_local_clk	:	out	std_logic	:=	'0';
		int_pmaif_pldif_tx_clkdiv	:	out	std_logic	:=	'0';
		int_pmaif_pldif_tx_clkdiv_user	:	out	std_logic	:=	'0';
		int_pmaif_pldif_uhsif_lock	:	out	std_logic	:=	'0';
		int_pmaif_pldif_uhsif_scan_chain_out	:	out	std_logic	:=	'0';
		int_pmaif_pldif_uhsif_tx_clk_out	:	out	std_logic	:=	'0';
		int_tx_dft_obsrv_clk	:	out	std_logic_vector(4 downto 0)	:=	"00000";
		pma_tx_elec_idle	:	out	std_logic	:=	'0';
		pma_tx_pma_data	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		pma_txpma_rstb	:	out	std_logic	:=	'0';
		tx_pma_data_loopback	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		tx_pma_uhsif_data_loopback	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		tx_prbs_gen_test	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		uhsif_test_out_1	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		uhsif_test_out_2	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		uhsif_test_out_3	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		write_en_ack	:	out	std_logic_vector(1 downto 0)	:=	"00"
	);
end component;

begin



inst : twentynm_hssi_tx_pcs_pma_interface_encrypted
	generic map (
		-- Instance parameters
		bypass_pma_txelecidle	=>	bypass_pma_txelecidle,
		channel_operation_mode	=>	channel_operation_mode,
		lpbk_en	=>	lpbk_en,
		master_clk_sel	=>	master_clk_sel,
		pcie_sub_prot_mode_tx	=>	pcie_sub_prot_mode_tx,
		pldif_datawidth_mode	=>	pldif_datawidth_mode,
		pma_dw_tx	=>	pma_dw_tx,
		pma_if_dft_en	=>	pma_if_dft_en,
		pmagate_en	=>	pmagate_en,
		prbs9_dwidth	=>	prbs9_dwidth,
		prbs_clken	=>	prbs_clken,
		prbs_gen_pat	=>	prbs_gen_pat,
		prot_mode_tx	=>	prot_mode_tx,
		reconfig_settings	=>	reconfig_settings,
		silicon_rev	=>	silicon_rev,
		sq_wave_num	=>	sq_wave_num,
		sqwgen_clken	=>	sqwgen_clken,
		sup_mode	=>	sup_mode,
		tx_dyn_polarity_inversion	=>	tx_dyn_polarity_inversion,
		tx_pma_data_sel	=>	tx_pma_data_sel,
		tx_static_polarity_inversion	=>	tx_static_polarity_inversion,
		uhsif_cnt_step_filt_before_lock	=>	uhsif_cnt_step_filt_before_lock,
		uhsif_cnt_thresh_filt_after_lock_value	=>	uhsif_cnt_thresh_filt_after_lock_value_int,
		uhsif_cnt_thresh_filt_before_lock	=>	uhsif_cnt_thresh_filt_before_lock,
		uhsif_dcn_test_update_period	=>	uhsif_dcn_test_update_period,
		uhsif_dcn_testmode_enable	=>	uhsif_dcn_testmode_enable,
		uhsif_dead_zone_count_thresh	=>	uhsif_dead_zone_count_thresh,
		uhsif_dead_zone_detection_enable	=>	uhsif_dead_zone_detection_enable,
		uhsif_dead_zone_obser_window	=>	uhsif_dead_zone_obser_window,
		uhsif_dead_zone_skip_size	=>	uhsif_dead_zone_skip_size,
		uhsif_delay_cell_index_sel	=>	uhsif_delay_cell_index_sel,
		uhsif_delay_cell_margin	=>	uhsif_delay_cell_margin,
		uhsif_delay_cell_static_index_value	=>	uhsif_delay_cell_static_index_value_int,
		uhsif_dft_dead_zone_control	=>	uhsif_dft_dead_zone_control,
		uhsif_dft_up_filt_control	=>	uhsif_dft_up_filt_control,
		uhsif_enable	=>	uhsif_enable,
		uhsif_lock_det_segsz_after_lock	=>	uhsif_lock_det_segsz_after_lock,
		uhsif_lock_det_segsz_before_lock	=>	uhsif_lock_det_segsz_before_lock,
		uhsif_lock_det_thresh_cnt_after_lock_value	=>	uhsif_lock_det_thresh_cnt_after_lock_value_int,
		uhsif_lock_det_thresh_cnt_before_lock_value	=>	uhsif_lock_det_thresh_cnt_before_lock_value_int,
		uhsif_lock_det_thresh_diff_after_lock_value	=>	uhsif_lock_det_thresh_diff_after_lock_value_int,
		uhsif_lock_det_thresh_diff_before_lock_value	=>	uhsif_lock_det_thresh_diff_before_lock_value_int
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		int_pmaif_10g_tx_clk_out	=>	int_pmaif_10g_tx_clk_out,
		int_pmaif_10g_tx_pma_data	=>	int_pmaif_10g_tx_pma_data,
		int_pmaif_10g_tx_pma_data_gate_val	=>	int_pmaif_10g_tx_pma_data_gate_val,
		int_pmaif_8g_pudr	=>	int_pmaif_8g_pudr,
		int_pmaif_8g_tx_clk_out	=>	int_pmaif_8g_tx_clk_out,
		int_pmaif_8g_tx_elec_idle	=>	int_pmaif_8g_tx_elec_idle,
		int_pmaif_g3_data_sel	=>	int_pmaif_g3_data_sel,
		int_pmaif_g3_pma_data_out	=>	int_pmaif_g3_pma_data_out,
		int_pmaif_g3_pma_tx_elec_idle	=>	int_pmaif_g3_pma_tx_elec_idle,
		int_pmaif_pldif_pmaif_tx_pld_rst_n	=>	int_pmaif_pldif_pmaif_tx_pld_rst_n,
		int_pmaif_pldif_polinv_tx	=>	int_pmaif_pldif_polinv_tx,
		int_pmaif_pldif_tx_data	=>	int_pmaif_pldif_tx_data,
		int_pmaif_pldif_txelecidle	=>	int_pmaif_pldif_txelecidle,
		int_pmaif_pldif_txpma_rstb	=>	int_pmaif_pldif_txpma_rstb,
		int_pmaif_pldif_uhsif_scan_chain_in	=>	int_pmaif_pldif_uhsif_scan_chain_in,
		int_pmaif_pldif_uhsif_tx_clk	=>	int_pmaif_pldif_uhsif_tx_clk,
		int_pmaif_pldif_uhsif_tx_data	=>	int_pmaif_pldif_uhsif_tx_data,
		pma_tx_clkdiv_user	=>	pma_tx_clkdiv_user,
		pma_tx_pma_clk	=>	pma_tx_pma_clk,
		refclk_dig	=>	refclk_dig,
		refclk_dig_uhsif	=>	refclk_dig_uhsif,
		scan_mode_n	=>	scan_mode_n,
		uhsif_scan_mode_n	=>	uhsif_scan_mode_n,
		uhsif_scan_shift_n	=>	uhsif_scan_shift_n,
		write_en	=>	write_en,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		avmm_user_dataout	=>	avmm_user_dataout,
		int_pmaif_10g_tx_pma_clk	=>	int_pmaif_10g_tx_pma_clk,
		int_pmaif_8g_txpma_local_clk	=>	int_pmaif_8g_txpma_local_clk,
		int_pmaif_pldif_tx_clkdiv	=>	int_pmaif_pldif_tx_clkdiv,
		int_pmaif_pldif_tx_clkdiv_user	=>	int_pmaif_pldif_tx_clkdiv_user,
		int_pmaif_pldif_uhsif_lock	=>	int_pmaif_pldif_uhsif_lock,
		int_pmaif_pldif_uhsif_scan_chain_out	=>	int_pmaif_pldif_uhsif_scan_chain_out,
		int_pmaif_pldif_uhsif_tx_clk_out	=>	int_pmaif_pldif_uhsif_tx_clk_out,
		int_tx_dft_obsrv_clk	=>	int_tx_dft_obsrv_clk,
		pma_tx_elec_idle	=>	pma_tx_elec_idle,
		pma_tx_pma_data	=>	pma_tx_pma_data,
		pma_txpma_rstb	=>	pma_txpma_rstb,
		tx_pma_data_loopback	=>	tx_pma_data_loopback,
		tx_pma_uhsif_data_loopback	=>	tx_pma_uhsif_data_loopback,
		tx_prbs_gen_test	=>	tx_prbs_gen_test,
		uhsif_test_out_1	=>	uhsif_test_out_1,
		uhsif_test_out_2	=>	uhsif_test_out_2,
		uhsif_test_out_3	=>	uhsif_test_out_3,
		write_en_ack	=>	write_en_ack
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;

entity	twentynm_hssi_tx_pld_pcs_interface	is
	generic (
		-- Entity parameters
		hd_10g_advanced_user_mode_tx	:	string	:=	"disable";
		hd_10g_channel_operation_mode	:	string	:=	"tx_rx_pair_enabled";
		hd_10g_ctrl_plane_bonding_tx	:	string	:=	"individual_tx";
		hd_10g_fifo_mode_tx	:	string	:=	"fifo_tx";
		hd_10g_low_latency_en_tx	:	string	:=	"enable";
		hd_10g_lpbk_en	:	string	:=	"disable";
		hd_10g_pma_dw_tx	:	string	:=	"pma_64b_tx";
		hd_10g_prot_mode_tx	:	string	:=	"disabled_prot_mode_tx";
		hd_10g_shared_fifo_width_tx	:	string	:=	"single_tx";
		hd_10g_sup_mode	:	string	:=	"user_mode";
		hd_8g_channel_operation_mode	:	string	:=	"tx_rx_pair_enabled";
		hd_8g_ctrl_plane_bonding_tx	:	string	:=	"individual_tx";
		hd_8g_fifo_mode_tx	:	string	:=	"fifo_tx";
		hd_8g_hip_mode	:	string	:=	"disable";
		hd_8g_lpbk_en	:	string	:=	"disable";
		hd_8g_pma_dw_tx	:	string	:=	"pma_8b_tx";
		hd_8g_prot_mode_tx	:	string	:=	"disabled_prot_mode_tx";
		hd_8g_sup_mode	:	string	:=	"user_mode";
		hd_chnl_channel_operation_mode	:	string	:=	"tx_rx_pair_enabled";
		hd_chnl_ctrl_plane_bonding_tx	:	string	:=	"individual_tx";
		hd_chnl_frequency_rules_en	:	string	:=	"disable";
		hd_chnl_func_mode	:	string	:=	"disable";
		hd_chnl_hclk_clk_hz	:	bit_vector	:=	B"000000000000000000000000000000";
		hd_chnl_hip_en	:	string	:=	"disable";
		hd_chnl_hrdrstctl_en	:	string	:=	"disable";
		hd_chnl_low_latency_en_tx	:	string	:=	"disable";
		hd_chnl_lpbk_en	:	string	:=	"disable";
		hd_chnl_pcs_tx_ac_pwr_uw_per_mhz	:	bit_vector	:=	B"00000000000000000000";
		hd_chnl_pcs_tx_pwr_scaling_clk	:	string	:=	"pma_tx_clk";
		hd_chnl_pld_8g_refclk_dig_nonatpg_mode_clk_hz	:	bit_vector	:=	B"000000000000000000000000000000";
		hd_chnl_pld_fifo_mode_tx	:	string	:=	"fifo_tx";
		hd_chnl_pld_pcs_refclk_dig_nonatpg_mode_clk_hz	:	bit_vector	:=	B"000000000000000000000000000000";
		hd_chnl_pld_tx_clk_hz	:	bit_vector	:=	B"000000000000000000000000000000";
		hd_chnl_pld_uhsif_tx_clk_hz	:	bit_vector	:=	B"000000000000000000000000000000";
		hd_chnl_pma_dw_tx	:	string	:=	"pma_8b_tx";
		hd_chnl_pma_tx_clk_hz	:	bit_vector	:=	B"000000000000000000000000000000";
		hd_chnl_prot_mode_tx	:	string	:=	"disabled_prot_mode_tx";
		hd_chnl_shared_fifo_width_tx	:	string	:=	"single_tx";
		hd_chnl_speed_grade	:	string	:=	"e2";
		hd_chnl_sup_mode	:	string	:=	"user_mode";
		hd_fifo_channel_operation_mode	:	string	:=	"tx_rx_pair_enabled";
		hd_fifo_prot_mode_tx	:	string	:=	"teng_mode_tx";
		hd_fifo_shared_fifo_width_tx	:	string	:=	"single_tx";
		hd_fifo_sup_mode	:	string	:=	"user_mode";
		hd_g3_prot_mode	:	string	:=	"disabled_prot_mode";
		hd_g3_sup_mode	:	string	:=	"user_mode";
		hd_krfec_channel_operation_mode	:	string	:=	"tx_rx_pair_enabled";
		hd_krfec_low_latency_en_tx	:	string	:=	"disable";
		hd_krfec_lpbk_en	:	string	:=	"disable";
		hd_krfec_prot_mode_tx	:	string	:=	"disabled_prot_mode_tx";
		hd_krfec_sup_mode	:	string	:=	"user_mode";
		hd_pldif_hrdrstctl_en	:	string	:=	"disable";
		hd_pldif_prot_mode_tx	:	string	:=	"disabled_prot_mode_tx";
		hd_pldif_sup_mode	:	string	:=	"user_mode";
		hd_pmaif_channel_operation_mode	:	string	:=	"tx_rx_pair_enabled";
		hd_pmaif_ctrl_plane_bonding	:	string	:=	"individual";
		hd_pmaif_lpbk_en	:	string	:=	"disable";
		hd_pmaif_pma_dw_tx	:	string	:=	"pma_8b_tx";
		hd_pmaif_prot_mode_tx	:	string	:=	"disabled_prot_mode_tx";
		hd_pmaif_sim_mode	:	string	:=	"disable";
		hd_pmaif_sup_mode	:	string	:=	"user_mode";
		pcs_tx_clk_out_sel	:	string	:=	"teng_clk_out";
		pcs_tx_clk_source	:	string	:=	"teng";
		pcs_tx_data_source	:	string	:=	"hip_disable";
		pcs_tx_delay1_clk_en	:	string	:=	"delay1_clk_disable";
		pcs_tx_delay1_clk_sel	:	string	:=	"pld_tx_clk";
		pcs_tx_delay1_ctrl	:	string	:=	"delay1_path0";
		pcs_tx_delay1_data_sel	:	string	:=	"one_ff_delay";
		pcs_tx_delay2_clk_en	:	string	:=	"delay2_clk_disable";
		pcs_tx_delay2_ctrl	:	string	:=	"delay2_path0";
		pcs_tx_output_sel	:	string	:=	"teng_output";
		reconfig_settings	:	string	:=	"{}";
		silicon_rev	:	string	:=	"20nm5es"
	);
	port (
		-- Entity ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		hip_tx_data	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		int_pldif_10g_tx_burst_en_exe	:	in	std_logic	:=	'0';
		int_pldif_10g_tx_clk_out	:	in	std_logic	:=	'0';
		int_pldif_10g_tx_clk_out_pld_if	:	in	std_logic	:=	'0';
		int_pldif_10g_tx_empty	:	in	std_logic	:=	'0';
		int_pldif_10g_tx_fifo_num	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		int_pldif_10g_tx_frame	:	in	std_logic	:=	'0';
		int_pldif_10g_tx_full	:	in	std_logic	:=	'0';
		int_pldif_10g_tx_pempty	:	in	std_logic	:=	'0';
		int_pldif_10g_tx_pfull	:	in	std_logic	:=	'0';
		int_pldif_10g_tx_wordslip_exe	:	in	std_logic	:=	'0';
		int_pldif_8g_empty_tx	:	in	std_logic	:=	'0';
		int_pldif_8g_full_tx	:	in	std_logic	:=	'0';
		int_pldif_8g_tx_clk_out	:	in	std_logic	:=	'0';
		int_pldif_8g_tx_clk_out_pld_if	:	in	std_logic	:=	'0';
		int_pldif_krfec_tx_alignment	:	in	std_logic	:=	'0';
		int_pldif_krfec_tx_frame	:	in	std_logic	:=	'0';
		int_pldif_pmaif_clkdiv_tx	:	in	std_logic	:=	'0';
		int_pldif_pmaif_clkdiv_tx_user	:	in	std_logic	:=	'0';
		int_pldif_pmaif_uhsif_tx_clk_out	:	in	std_logic	:=	'0';
		pld_10g_krfec_tx_pld_rst_n	:	in	std_logic	:=	'0';
		pld_10g_tx_bitslip	:	in	std_logic_vector(6 downto 0)	:=	"0000000";
		pld_10g_tx_burst_en	:	in	std_logic	:=	'0';
		pld_10g_tx_data_valid	:	in	std_logic	:=	'0';
		pld_10g_tx_diag_status	:	in	std_logic_vector(1 downto 0)	:=	"00";
		pld_10g_tx_wordslip	:	in	std_logic	:=	'0';
		pld_8g_g3_tx_pld_rst_n	:	in	std_logic	:=	'0';
		pld_8g_rddisable_tx	:	in	std_logic	:=	'0';
		pld_8g_tx_boundary_sel	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		pld_8g_wrenable_tx	:	in	std_logic	:=	'0';
		pld_partial_reconfig	:	in	std_logic	:=	'0';
		pld_pma_txpma_rstb	:	in	std_logic	:=	'0';
		pld_pmaif_tx_pld_rst_n	:	in	std_logic	:=	'0';
		pld_polinv_tx	:	in	std_logic	:=	'0';
		pld_tx_clk	:	in	std_logic	:=	'0';
		pld_tx_control	:	in	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		pld_tx_data	:	in	std_logic_vector(127 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		pld_txelecidle	:	in	std_logic	:=	'0';
		pld_uhsif_tx_clk	:	in	std_logic	:=	'0';
		scan_mode_n	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		hip_clk_out_div_by_2_wire	:	out	std_logic	:=	'0';
		hip_clk_out_wire	:	out	std_logic	:=	'0';
		pld_10g_tx_burst_en_exe_10g_fastreg	:	out	std_logic	:=	'0';
		pld_10g_tx_burst_en_exe_plddirect_reg	:	out	std_logic	:=	'0';
		pld_10g_tx_data_valid_2ff_delay1_fastreg	:	out	std_logic	:=	'0';
		pld_10g_tx_data_valid_2ff_delay3_fastreg	:	out	std_logic	:=	'0';
		pld_10g_tx_data_valid_2ff_delay4_fastreg	:	out	std_logic	:=	'0';
		pld_10g_tx_data_valid_2ff_delay4_plddirect_fastreg	:	out	std_logic	:=	'0';
		pld_10g_tx_data_valid_2ff_delay6_fastreg	:	out	std_logic	:=	'0';
		pld_10g_tx_data_valid_2ff_delay6_plddirect_fastreg	:	out	std_logic	:=	'0';
		pld_10g_tx_data_valid_fastreg	:	out	std_logic	:=	'0';
		pld_10g_tx_data_valid_plddirect_fastreg	:	out	std_logic	:=	'0';
		pld_pcs_tx_clk_out_pma_wire	:	out	std_logic	:=	'0';
		pld_pma_tx_clk_out_wire	:	out	std_logic	:=	'0';
		pld_pmaif_tx_pld_rst_n_reg	:	out	std_logic	:=	'0';
		pld_polinv_tx_10g_pcsdirect_reg	:	out	std_logic	:=	'0';
		pld_polinv_tx_8g_reg	:	out	std_logic	:=	'0';
		pld_polinv_tx_pat_reg	:	out	std_logic	:=	'0';
		pld_tx_clk_fifo	:	out	std_logic	:=	'0';
		pld_tx_control_fifo	:	out	std_logic	:=	'0';
		pld_tx_control_hi_10g_reg	:	out	std_logic	:=	'0';
		pld_tx_control_lo_10g_2ff_delay4_fastreg	:	out	std_logic	:=	'0';
		pld_tx_control_lo_10g_2ff_delay6_fastreg	:	out	std_logic	:=	'0';
		pld_tx_control_lo_10g_fastreg	:	out	std_logic	:=	'0';
		pld_tx_control_lo_8g_2ff_delay4_fastreg	:	out	std_logic	:=	'0';
		pld_tx_control_lo_8g_2ff_delay6_fastreg	:	out	std_logic	:=	'0';
		pld_tx_control_lo_8g_fastreg	:	out	std_logic	:=	'0';
		pld_tx_control_lo_plddirect_2ff_delay1_fastreg	:	out	std_logic	:=	'0';
		pld_tx_control_lo_plddirect_2ff_delay3_fastreg	:	out	std_logic	:=	'0';
		pld_tx_control_lo_plddirect_2ff_delay4_fastreg	:	out	std_logic	:=	'0';
		pld_tx_control_lo_plddirect_2ff_delay6_fastreg	:	out	std_logic	:=	'0';
		pld_tx_control_lo_plddirect_fastreg	:	out	std_logic	:=	'0';
		pld_tx_control_lo_plddirect_reg	:	out	std_logic	:=	'0';
		pld_tx_data_hi_reg	:	out	std_logic	:=	'0';
		pld_tx_data_lo_10g_2ff_delay4_fastreg	:	out	std_logic	:=	'0';
		pld_tx_data_lo_10g_2ff_delay6_fastreg	:	out	std_logic	:=	'0';
		pld_tx_data_lo_10g_fastreg	:	out	std_logic	:=	'0';
		pld_tx_data_lo_8g_2ff_delay4_fastreg	:	out	std_logic	:=	'0';
		pld_tx_data_lo_8g_2ff_delay6_fastreg	:	out	std_logic	:=	'0';
		pld_tx_data_lo_8g_fastreg	:	out	std_logic	:=	'0';
		pld_tx_data_lo_plddirect_2ff_delay1_fastreg	:	out	std_logic	:=	'0';
		pld_tx_data_lo_plddirect_2ff_delay3_fastreg	:	out	std_logic	:=	'0';
		pld_tx_data_lo_plddirect_2ff_delay4_fastreg	:	out	std_logic	:=	'0';
		pld_tx_data_lo_plddirect_2ff_delay6_fastreg	:	out	std_logic	:=	'0';
		pld_tx_data_lo_plddirect_fastreg	:	out	std_logic	:=	'0';
		pld_tx_data_lo_plddirect_reg	:	out	std_logic	:=	'0';
		pld_uhsif_reg	:	out	std_logic	:=	'0';
		pma_tx_pma_clk_reg	:	out	std_logic	:=	'0';
		hip_tx_clk	:	out	std_logic	:=	'0';
		int_pldif_10g_tx_bitslip	:	out	std_logic_vector(6 downto 0)	:=	"0000000";
		int_pldif_10g_tx_burst_en	:	out	std_logic	:=	'0';
		int_pldif_10g_tx_control	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		int_pldif_10g_tx_control_reg	:	out	std_logic_vector(8 downto 0)	:=	"000000000";
		int_pldif_10g_tx_data	:	out	std_logic_vector(127 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		int_pldif_10g_tx_data_reg	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		int_pldif_10g_tx_data_valid	:	out	std_logic	:=	'0';
		int_pldif_10g_tx_data_valid_reg	:	out	std_logic	:=	'0';
		int_pldif_10g_tx_diag_status	:	out	std_logic_vector(1 downto 0)	:=	"00";
		int_pldif_10g_tx_pld_clk	:	out	std_logic	:=	'0';
		int_pldif_10g_tx_pld_rst_n	:	out	std_logic	:=	'0';
		int_pldif_10g_tx_wordslip	:	out	std_logic	:=	'0';
		int_pldif_8g_pld_tx_clk	:	out	std_logic	:=	'0';
		int_pldif_8g_powerdown	:	out	std_logic_vector(1 downto 0)	:=	"00";
		int_pldif_8g_rddisable_tx	:	out	std_logic	:=	'0';
		int_pldif_8g_rev_loopbk	:	out	std_logic	:=	'0';
		int_pldif_8g_tx_blk_start	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		int_pldif_8g_tx_boundary_sel	:	out	std_logic_vector(4 downto 0)	:=	"00000";
		int_pldif_8g_tx_data_valid	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		int_pldif_8g_tx_sync_hdr	:	out	std_logic_vector(1 downto 0)	:=	"00";
		int_pldif_8g_txd	:	out	std_logic_vector(43 downto 0)	:=	"00000000000000000000000000000000000000000000";
		int_pldif_8g_txd_fast_reg	:	out	std_logic_vector(43 downto 0)	:=	"00000000000000000000000000000000000000000000";
		int_pldif_8g_txdeemph	:	out	std_logic	:=	'0';
		int_pldif_8g_txdetectrxloopback	:	out	std_logic	:=	'0';
		int_pldif_8g_txelecidle	:	out	std_logic	:=	'0';
		int_pldif_8g_txmargin	:	out	std_logic_vector(2 downto 0)	:=	"000";
		int_pldif_8g_txswing	:	out	std_logic	:=	'0';
		int_pldif_8g_txurstpcs_n	:	out	std_logic	:=	'0';
		int_pldif_8g_wrenable_tx	:	out	std_logic	:=	'0';
		int_pldif_pmaif_8g_txurstpcs_n	:	out	std_logic	:=	'0';
		int_pldif_pmaif_polinv_tx	:	out	std_logic	:=	'0';
		int_pldif_pmaif_tx_data	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		int_pldif_pmaif_tx_pld_clk	:	out	std_logic	:=	'0';
		int_pldif_pmaif_tx_pld_rst_n	:	out	std_logic	:=	'0';
		int_pldif_pmaif_txelecidle	:	out	std_logic	:=	'0';
		int_pldif_pmaif_txpma_rstb	:	out	std_logic	:=	'0';
		int_pldif_pmaif_uhsif_tx_clk	:	out	std_logic	:=	'0';
		int_pldif_pmaif_uhsif_tx_data	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		pld_10g_krfec_tx_frame	:	out	std_logic	:=	'0';
		pld_10g_tx_burst_en_exe	:	out	std_logic	:=	'0';
		pld_10g_tx_empty	:	out	std_logic	:=	'0';
		pld_10g_tx_fifo_num	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		pld_10g_tx_full	:	out	std_logic	:=	'0';
		pld_10g_tx_pempty	:	out	std_logic	:=	'0';
		pld_10g_tx_pfull	:	out	std_logic	:=	'0';
		pld_10g_tx_wordslip_exe	:	out	std_logic	:=	'0';
		pld_8g_empty_tx	:	out	std_logic	:=	'0';
		pld_8g_full_tx	:	out	std_logic	:=	'0';
		pld_krfec_tx_alignment	:	out	std_logic	:=	'0';
		pld_pcs_tx_clk_out	:	out	std_logic	:=	'0';
		pld_pma_clkdiv_tx_user	:	out	std_logic	:=	'0';
		pld_pma_tx_clk_out	:	out	std_logic	:=	'0';
		pld_uhsif_tx_clk_out	:	out	std_logic	:=	'0'
	);
end twentynm_hssi_tx_pld_pcs_interface;

architecture behavior of twentynm_hssi_tx_pld_pcs_interface	is

constant hd_chnl_hclk_clk_hz_int	:	integer	:=	bin2int(hd_chnl_hclk_clk_hz);
constant hd_chnl_pcs_tx_ac_pwr_uw_per_mhz_int	:	integer	:=	bin2int(hd_chnl_pcs_tx_ac_pwr_uw_per_mhz);
constant hd_chnl_pld_8g_refclk_dig_nonatpg_mode_clk_hz_int	:	integer	:=	bin2int(hd_chnl_pld_8g_refclk_dig_nonatpg_mode_clk_hz);
constant hd_chnl_pld_pcs_refclk_dig_nonatpg_mode_clk_hz_int	:	integer	:=	bin2int(hd_chnl_pld_pcs_refclk_dig_nonatpg_mode_clk_hz);
constant hd_chnl_pld_tx_clk_hz_int	:	integer	:=	bin2int(hd_chnl_pld_tx_clk_hz);
constant hd_chnl_pld_uhsif_tx_clk_hz_int	:	integer	:=	bin2int(hd_chnl_pld_uhsif_tx_clk_hz);
constant hd_chnl_pma_tx_clk_hz_int	:	integer	:=	bin2int(hd_chnl_pma_tx_clk_hz);



component	twentynm_hssi_tx_pld_pcs_interface_encrypted
	generic (
		-- Architecture parameters
		hd_10g_advanced_user_mode_tx	:	string	:=	"disable";
		hd_10g_channel_operation_mode	:	string	:=	"tx_rx_pair_enabled";
		hd_10g_ctrl_plane_bonding_tx	:	string	:=	"individual_tx";
		hd_10g_fifo_mode_tx	:	string	:=	"fifo_tx";
		hd_10g_low_latency_en_tx	:	string	:=	"enable";
		hd_10g_lpbk_en	:	string	:=	"disable";
		hd_10g_pma_dw_tx	:	string	:=	"pma_64b_tx";
		hd_10g_prot_mode_tx	:	string	:=	"disabled_prot_mode_tx";
		hd_10g_shared_fifo_width_tx	:	string	:=	"single_tx";
		hd_10g_sup_mode	:	string	:=	"user_mode";
		hd_8g_channel_operation_mode	:	string	:=	"tx_rx_pair_enabled";
		hd_8g_ctrl_plane_bonding_tx	:	string	:=	"individual_tx";
		hd_8g_fifo_mode_tx	:	string	:=	"fifo_tx";
		hd_8g_hip_mode	:	string	:=	"disable";
		hd_8g_lpbk_en	:	string	:=	"disable";
		hd_8g_pma_dw_tx	:	string	:=	"pma_8b_tx";
		hd_8g_prot_mode_tx	:	string	:=	"disabled_prot_mode_tx";
		hd_8g_sup_mode	:	string	:=	"user_mode";
		hd_chnl_channel_operation_mode	:	string	:=	"tx_rx_pair_enabled";
		hd_chnl_ctrl_plane_bonding_tx	:	string	:=	"individual_tx";
		hd_chnl_frequency_rules_en	:	string	:=	"disable";
		hd_chnl_func_mode	:	string	:=	"disable";
		hd_chnl_hclk_clk_hz	:	integer	:=	0;
		hd_chnl_hip_en	:	string	:=	"disable";
		hd_chnl_hrdrstctl_en	:	string	:=	"disable";
		hd_chnl_low_latency_en_tx	:	string	:=	"disable";
		hd_chnl_lpbk_en	:	string	:=	"disable";
		hd_chnl_pcs_tx_ac_pwr_uw_per_mhz	:	integer	:=	0;
		hd_chnl_pcs_tx_pwr_scaling_clk	:	string	:=	"pma_tx_clk";
		hd_chnl_pld_8g_refclk_dig_nonatpg_mode_clk_hz	:	integer	:=	0;
		hd_chnl_pld_fifo_mode_tx	:	string	:=	"fifo_tx";
		hd_chnl_pld_pcs_refclk_dig_nonatpg_mode_clk_hz	:	integer	:=	0;
		hd_chnl_pld_tx_clk_hz	:	integer	:=	0;
		hd_chnl_pld_uhsif_tx_clk_hz	:	integer	:=	0;
		hd_chnl_pma_dw_tx	:	string	:=	"pma_8b_tx";
		hd_chnl_pma_tx_clk_hz	:	integer	:=	0;
		hd_chnl_prot_mode_tx	:	string	:=	"disabled_prot_mode_tx";
		hd_chnl_shared_fifo_width_tx	:	string	:=	"single_tx";
		hd_chnl_speed_grade	:	string	:=	"e2";
		hd_chnl_sup_mode	:	string	:=	"user_mode";
		hd_fifo_channel_operation_mode	:	string	:=	"tx_rx_pair_enabled";
		hd_fifo_prot_mode_tx	:	string	:=	"teng_mode_tx";
		hd_fifo_shared_fifo_width_tx	:	string	:=	"single_tx";
		hd_fifo_sup_mode	:	string	:=	"user_mode";
		hd_g3_prot_mode	:	string	:=	"disabled_prot_mode";
		hd_g3_sup_mode	:	string	:=	"user_mode";
		hd_krfec_channel_operation_mode	:	string	:=	"tx_rx_pair_enabled";
		hd_krfec_low_latency_en_tx	:	string	:=	"disable";
		hd_krfec_lpbk_en	:	string	:=	"disable";
		hd_krfec_prot_mode_tx	:	string	:=	"disabled_prot_mode_tx";
		hd_krfec_sup_mode	:	string	:=	"user_mode";
		hd_pldif_hrdrstctl_en	:	string	:=	"disable";
		hd_pldif_prot_mode_tx	:	string	:=	"disabled_prot_mode_tx";
		hd_pldif_sup_mode	:	string	:=	"user_mode";
		hd_pmaif_channel_operation_mode	:	string	:=	"tx_rx_pair_enabled";
		hd_pmaif_ctrl_plane_bonding	:	string	:=	"individual";
		hd_pmaif_lpbk_en	:	string	:=	"disable";
		hd_pmaif_pma_dw_tx	:	string	:=	"pma_8b_tx";
		hd_pmaif_prot_mode_tx	:	string	:=	"disabled_prot_mode_tx";
		hd_pmaif_sim_mode	:	string	:=	"disable";
		hd_pmaif_sup_mode	:	string	:=	"user_mode";
		pcs_tx_clk_out_sel	:	string	:=	"teng_clk_out";
		pcs_tx_clk_source	:	string	:=	"teng";
		pcs_tx_data_source	:	string	:=	"hip_disable";
		pcs_tx_delay1_clk_en	:	string	:=	"delay1_clk_disable";
		pcs_tx_delay1_clk_sel	:	string	:=	"pld_tx_clk";
		pcs_tx_delay1_ctrl	:	string	:=	"delay1_path0";
		pcs_tx_delay1_data_sel	:	string	:=	"one_ff_delay";
		pcs_tx_delay2_clk_en	:	string	:=	"delay2_clk_disable";
		pcs_tx_delay2_ctrl	:	string	:=	"delay2_path0";
		pcs_tx_output_sel	:	string	:=	"teng_output";
		reconfig_settings	:	string	:=	"{}";
		silicon_rev	:	string	:=	"20nm5es"
	);
	port (
		-- Architecture ports
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:=	"000000000";
		avmmclk	:	in	std_logic	:=	'0';
		avmmread	:	in	std_logic	:=	'0';
		avmmrstn	:	in	std_logic	:=	'0';
		avmmwrite	:	in	std_logic	:=	'0';
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		hip_tx_data	:	in	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		int_pldif_10g_tx_burst_en_exe	:	in	std_logic	:=	'0';
		int_pldif_10g_tx_clk_out	:	in	std_logic	:=	'0';
		int_pldif_10g_tx_clk_out_pld_if	:	in	std_logic	:=	'0';
		int_pldif_10g_tx_empty	:	in	std_logic	:=	'0';
		int_pldif_10g_tx_fifo_num	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		int_pldif_10g_tx_frame	:	in	std_logic	:=	'0';
		int_pldif_10g_tx_full	:	in	std_logic	:=	'0';
		int_pldif_10g_tx_pempty	:	in	std_logic	:=	'0';
		int_pldif_10g_tx_pfull	:	in	std_logic	:=	'0';
		int_pldif_10g_tx_wordslip_exe	:	in	std_logic	:=	'0';
		int_pldif_8g_empty_tx	:	in	std_logic	:=	'0';
		int_pldif_8g_full_tx	:	in	std_logic	:=	'0';
		int_pldif_8g_tx_clk_out	:	in	std_logic	:=	'0';
		int_pldif_8g_tx_clk_out_pld_if	:	in	std_logic	:=	'0';
		int_pldif_krfec_tx_alignment	:	in	std_logic	:=	'0';
		int_pldif_krfec_tx_frame	:	in	std_logic	:=	'0';
		int_pldif_pmaif_clkdiv_tx	:	in	std_logic	:=	'0';
		int_pldif_pmaif_clkdiv_tx_user	:	in	std_logic	:=	'0';
		int_pldif_pmaif_uhsif_tx_clk_out	:	in	std_logic	:=	'0';
		pld_10g_krfec_tx_pld_rst_n	:	in	std_logic	:=	'0';
		pld_10g_tx_bitslip	:	in	std_logic_vector(6 downto 0)	:=	"0000000";
		pld_10g_tx_burst_en	:	in	std_logic	:=	'0';
		pld_10g_tx_data_valid	:	in	std_logic	:=	'0';
		pld_10g_tx_diag_status	:	in	std_logic_vector(1 downto 0)	:=	"00";
		pld_10g_tx_wordslip	:	in	std_logic	:=	'0';
		pld_8g_g3_tx_pld_rst_n	:	in	std_logic	:=	'0';
		pld_8g_rddisable_tx	:	in	std_logic	:=	'0';
		pld_8g_tx_boundary_sel	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		pld_8g_wrenable_tx	:	in	std_logic	:=	'0';
		pld_partial_reconfig	:	in	std_logic	:=	'0';
		pld_pma_txpma_rstb	:	in	std_logic	:=	'0';
		pld_pmaif_tx_pld_rst_n	:	in	std_logic	:=	'0';
		pld_polinv_tx	:	in	std_logic	:=	'0';
		pld_tx_clk	:	in	std_logic	:=	'0';
		pld_tx_control	:	in	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		pld_tx_data	:	in	std_logic_vector(127 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		pld_txelecidle	:	in	std_logic	:=	'0';
		pld_uhsif_tx_clk	:	in	std_logic	:=	'0';
		scan_mode_n	:	in	std_logic	:=	'0';
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		blockselect	:	out	std_logic	:=	'0';
		hip_clk_out_div_by_2_wire	:	out	std_logic	:=	'0';
		hip_clk_out_wire	:	out	std_logic	:=	'0';
		pld_10g_tx_burst_en_exe_10g_fastreg	:	out	std_logic	:=	'0';
		pld_10g_tx_burst_en_exe_plddirect_reg	:	out	std_logic	:=	'0';
		pld_10g_tx_data_valid_2ff_delay1_fastreg	:	out	std_logic	:=	'0';
		pld_10g_tx_data_valid_2ff_delay3_fastreg	:	out	std_logic	:=	'0';
		pld_10g_tx_data_valid_2ff_delay4_fastreg	:	out	std_logic	:=	'0';
		pld_10g_tx_data_valid_2ff_delay4_plddirect_fastreg	:	out	std_logic	:=	'0';
		pld_10g_tx_data_valid_2ff_delay6_fastreg	:	out	std_logic	:=	'0';
		pld_10g_tx_data_valid_2ff_delay6_plddirect_fastreg	:	out	std_logic	:=	'0';
		pld_10g_tx_data_valid_fastreg	:	out	std_logic	:=	'0';
		pld_10g_tx_data_valid_plddirect_fastreg	:	out	std_logic	:=	'0';
		pld_pcs_tx_clk_out_pma_wire	:	out	std_logic	:=	'0';
		pld_pma_tx_clk_out_wire	:	out	std_logic	:=	'0';
		pld_pmaif_tx_pld_rst_n_reg	:	out	std_logic	:=	'0';
		pld_polinv_tx_10g_pcsdirect_reg	:	out	std_logic	:=	'0';
		pld_polinv_tx_8g_reg	:	out	std_logic	:=	'0';
		pld_polinv_tx_pat_reg	:	out	std_logic	:=	'0';
		pld_tx_clk_fifo	:	out	std_logic	:=	'0';
		pld_tx_control_fifo	:	out	std_logic	:=	'0';
		pld_tx_control_hi_10g_reg	:	out	std_logic	:=	'0';
		pld_tx_control_lo_10g_2ff_delay4_fastreg	:	out	std_logic	:=	'0';
		pld_tx_control_lo_10g_2ff_delay6_fastreg	:	out	std_logic	:=	'0';
		pld_tx_control_lo_10g_fastreg	:	out	std_logic	:=	'0';
		pld_tx_control_lo_8g_2ff_delay4_fastreg	:	out	std_logic	:=	'0';
		pld_tx_control_lo_8g_2ff_delay6_fastreg	:	out	std_logic	:=	'0';
		pld_tx_control_lo_8g_fastreg	:	out	std_logic	:=	'0';
		pld_tx_control_lo_plddirect_2ff_delay1_fastreg	:	out	std_logic	:=	'0';
		pld_tx_control_lo_plddirect_2ff_delay3_fastreg	:	out	std_logic	:=	'0';
		pld_tx_control_lo_plddirect_2ff_delay4_fastreg	:	out	std_logic	:=	'0';
		pld_tx_control_lo_plddirect_2ff_delay6_fastreg	:	out	std_logic	:=	'0';
		pld_tx_control_lo_plddirect_fastreg	:	out	std_logic	:=	'0';
		pld_tx_control_lo_plddirect_reg	:	out	std_logic	:=	'0';
		pld_tx_data_hi_reg	:	out	std_logic	:=	'0';
		pld_tx_data_lo_10g_2ff_delay4_fastreg	:	out	std_logic	:=	'0';
		pld_tx_data_lo_10g_2ff_delay6_fastreg	:	out	std_logic	:=	'0';
		pld_tx_data_lo_10g_fastreg	:	out	std_logic	:=	'0';
		pld_tx_data_lo_8g_2ff_delay4_fastreg	:	out	std_logic	:=	'0';
		pld_tx_data_lo_8g_2ff_delay6_fastreg	:	out	std_logic	:=	'0';
		pld_tx_data_lo_8g_fastreg	:	out	std_logic	:=	'0';
		pld_tx_data_lo_plddirect_2ff_delay1_fastreg	:	out	std_logic	:=	'0';
		pld_tx_data_lo_plddirect_2ff_delay3_fastreg	:	out	std_logic	:=	'0';
		pld_tx_data_lo_plddirect_2ff_delay4_fastreg	:	out	std_logic	:=	'0';
		pld_tx_data_lo_plddirect_2ff_delay6_fastreg	:	out	std_logic	:=	'0';
		pld_tx_data_lo_plddirect_fastreg	:	out	std_logic	:=	'0';
		pld_tx_data_lo_plddirect_reg	:	out	std_logic	:=	'0';
		pld_uhsif_reg	:	out	std_logic	:=	'0';
		pma_tx_pma_clk_reg	:	out	std_logic	:=	'0';
		hip_tx_clk	:	out	std_logic	:=	'0';
		int_pldif_10g_tx_bitslip	:	out	std_logic_vector(6 downto 0)	:=	"0000000";
		int_pldif_10g_tx_burst_en	:	out	std_logic	:=	'0';
		int_pldif_10g_tx_control	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		int_pldif_10g_tx_control_reg	:	out	std_logic_vector(8 downto 0)	:=	"000000000";
		int_pldif_10g_tx_data	:	out	std_logic_vector(127 downto 0)	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		int_pldif_10g_tx_data_reg	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		int_pldif_10g_tx_data_valid	:	out	std_logic	:=	'0';
		int_pldif_10g_tx_data_valid_reg	:	out	std_logic	:=	'0';
		int_pldif_10g_tx_diag_status	:	out	std_logic_vector(1 downto 0)	:=	"00";
		int_pldif_10g_tx_pld_clk	:	out	std_logic	:=	'0';
		int_pldif_10g_tx_pld_rst_n	:	out	std_logic	:=	'0';
		int_pldif_10g_tx_wordslip	:	out	std_logic	:=	'0';
		int_pldif_8g_pld_tx_clk	:	out	std_logic	:=	'0';
		int_pldif_8g_powerdown	:	out	std_logic_vector(1 downto 0)	:=	"00";
		int_pldif_8g_rddisable_tx	:	out	std_logic	:=	'0';
		int_pldif_8g_rev_loopbk	:	out	std_logic	:=	'0';
		int_pldif_8g_tx_blk_start	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		int_pldif_8g_tx_boundary_sel	:	out	std_logic_vector(4 downto 0)	:=	"00000";
		int_pldif_8g_tx_data_valid	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		int_pldif_8g_tx_sync_hdr	:	out	std_logic_vector(1 downto 0)	:=	"00";
		int_pldif_8g_txd	:	out	std_logic_vector(43 downto 0)	:=	"00000000000000000000000000000000000000000000";
		int_pldif_8g_txd_fast_reg	:	out	std_logic_vector(43 downto 0)	:=	"00000000000000000000000000000000000000000000";
		int_pldif_8g_txdeemph	:	out	std_logic	:=	'0';
		int_pldif_8g_txdetectrxloopback	:	out	std_logic	:=	'0';
		int_pldif_8g_txelecidle	:	out	std_logic	:=	'0';
		int_pldif_8g_txmargin	:	out	std_logic_vector(2 downto 0)	:=	"000";
		int_pldif_8g_txswing	:	out	std_logic	:=	'0';
		int_pldif_8g_txurstpcs_n	:	out	std_logic	:=	'0';
		int_pldif_8g_wrenable_tx	:	out	std_logic	:=	'0';
		int_pldif_pmaif_8g_txurstpcs_n	:	out	std_logic	:=	'0';
		int_pldif_pmaif_polinv_tx	:	out	std_logic	:=	'0';
		int_pldif_pmaif_tx_data	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		int_pldif_pmaif_tx_pld_clk	:	out	std_logic	:=	'0';
		int_pldif_pmaif_tx_pld_rst_n	:	out	std_logic	:=	'0';
		int_pldif_pmaif_txelecidle	:	out	std_logic	:=	'0';
		int_pldif_pmaif_txpma_rstb	:	out	std_logic	:=	'0';
		int_pldif_pmaif_uhsif_tx_clk	:	out	std_logic	:=	'0';
		int_pldif_pmaif_uhsif_tx_data	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		pld_10g_krfec_tx_frame	:	out	std_logic	:=	'0';
		pld_10g_tx_burst_en_exe	:	out	std_logic	:=	'0';
		pld_10g_tx_empty	:	out	std_logic	:=	'0';
		pld_10g_tx_fifo_num	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		pld_10g_tx_full	:	out	std_logic	:=	'0';
		pld_10g_tx_pempty	:	out	std_logic	:=	'0';
		pld_10g_tx_pfull	:	out	std_logic	:=	'0';
		pld_10g_tx_wordslip_exe	:	out	std_logic	:=	'0';
		pld_8g_empty_tx	:	out	std_logic	:=	'0';
		pld_8g_full_tx	:	out	std_logic	:=	'0';
		pld_krfec_tx_alignment	:	out	std_logic	:=	'0';
		pld_pcs_tx_clk_out	:	out	std_logic	:=	'0';
		pld_pma_clkdiv_tx_user	:	out	std_logic	:=	'0';
		pld_pma_tx_clk_out	:	out	std_logic	:=	'0';
		pld_uhsif_tx_clk_out	:	out	std_logic	:=	'0'
	);
end component;

begin



inst : twentynm_hssi_tx_pld_pcs_interface_encrypted
	generic map (
		-- Instance parameters
		hd_10g_advanced_user_mode_tx	=>	hd_10g_advanced_user_mode_tx,
		hd_10g_channel_operation_mode	=>	hd_10g_channel_operation_mode,
		hd_10g_ctrl_plane_bonding_tx	=>	hd_10g_ctrl_plane_bonding_tx,
		hd_10g_fifo_mode_tx	=>	hd_10g_fifo_mode_tx,
		hd_10g_low_latency_en_tx	=>	hd_10g_low_latency_en_tx,
		hd_10g_lpbk_en	=>	hd_10g_lpbk_en,
		hd_10g_pma_dw_tx	=>	hd_10g_pma_dw_tx,
		hd_10g_prot_mode_tx	=>	hd_10g_prot_mode_tx,
		hd_10g_shared_fifo_width_tx	=>	hd_10g_shared_fifo_width_tx,
		hd_10g_sup_mode	=>	hd_10g_sup_mode,
		hd_8g_channel_operation_mode	=>	hd_8g_channel_operation_mode,
		hd_8g_ctrl_plane_bonding_tx	=>	hd_8g_ctrl_plane_bonding_tx,
		hd_8g_fifo_mode_tx	=>	hd_8g_fifo_mode_tx,
		hd_8g_hip_mode	=>	hd_8g_hip_mode,
		hd_8g_lpbk_en	=>	hd_8g_lpbk_en,
		hd_8g_pma_dw_tx	=>	hd_8g_pma_dw_tx,
		hd_8g_prot_mode_tx	=>	hd_8g_prot_mode_tx,
		hd_8g_sup_mode	=>	hd_8g_sup_mode,
		hd_chnl_channel_operation_mode	=>	hd_chnl_channel_operation_mode,
		hd_chnl_ctrl_plane_bonding_tx	=>	hd_chnl_ctrl_plane_bonding_tx,
		hd_chnl_frequency_rules_en	=>	hd_chnl_frequency_rules_en,
		hd_chnl_func_mode	=>	hd_chnl_func_mode,
		hd_chnl_hclk_clk_hz	=>	hd_chnl_hclk_clk_hz_int,
		hd_chnl_hip_en	=>	hd_chnl_hip_en,
		hd_chnl_hrdrstctl_en	=>	hd_chnl_hrdrstctl_en,
		hd_chnl_low_latency_en_tx	=>	hd_chnl_low_latency_en_tx,
		hd_chnl_lpbk_en	=>	hd_chnl_lpbk_en,
		hd_chnl_pcs_tx_ac_pwr_uw_per_mhz	=>	hd_chnl_pcs_tx_ac_pwr_uw_per_mhz_int,
		hd_chnl_pcs_tx_pwr_scaling_clk	=>	hd_chnl_pcs_tx_pwr_scaling_clk,
		hd_chnl_pld_8g_refclk_dig_nonatpg_mode_clk_hz	=>	hd_chnl_pld_8g_refclk_dig_nonatpg_mode_clk_hz_int,
		hd_chnl_pld_fifo_mode_tx	=>	hd_chnl_pld_fifo_mode_tx,
		hd_chnl_pld_pcs_refclk_dig_nonatpg_mode_clk_hz	=>	hd_chnl_pld_pcs_refclk_dig_nonatpg_mode_clk_hz_int,
		hd_chnl_pld_tx_clk_hz	=>	hd_chnl_pld_tx_clk_hz_int,
		hd_chnl_pld_uhsif_tx_clk_hz	=>	hd_chnl_pld_uhsif_tx_clk_hz_int,
		hd_chnl_pma_dw_tx	=>	hd_chnl_pma_dw_tx,
		hd_chnl_pma_tx_clk_hz	=>	hd_chnl_pma_tx_clk_hz_int,
		hd_chnl_prot_mode_tx	=>	hd_chnl_prot_mode_tx,
		hd_chnl_shared_fifo_width_tx	=>	hd_chnl_shared_fifo_width_tx,
		hd_chnl_speed_grade	=>	hd_chnl_speed_grade,
		hd_chnl_sup_mode	=>	hd_chnl_sup_mode,
		hd_fifo_channel_operation_mode	=>	hd_fifo_channel_operation_mode,
		hd_fifo_prot_mode_tx	=>	hd_fifo_prot_mode_tx,
		hd_fifo_shared_fifo_width_tx	=>	hd_fifo_shared_fifo_width_tx,
		hd_fifo_sup_mode	=>	hd_fifo_sup_mode,
		hd_g3_prot_mode	=>	hd_g3_prot_mode,
		hd_g3_sup_mode	=>	hd_g3_sup_mode,
		hd_krfec_channel_operation_mode	=>	hd_krfec_channel_operation_mode,
		hd_krfec_low_latency_en_tx	=>	hd_krfec_low_latency_en_tx,
		hd_krfec_lpbk_en	=>	hd_krfec_lpbk_en,
		hd_krfec_prot_mode_tx	=>	hd_krfec_prot_mode_tx,
		hd_krfec_sup_mode	=>	hd_krfec_sup_mode,
		hd_pldif_hrdrstctl_en	=>	hd_pldif_hrdrstctl_en,
		hd_pldif_prot_mode_tx	=>	hd_pldif_prot_mode_tx,
		hd_pldif_sup_mode	=>	hd_pldif_sup_mode,
		hd_pmaif_channel_operation_mode	=>	hd_pmaif_channel_operation_mode,
		hd_pmaif_ctrl_plane_bonding	=>	hd_pmaif_ctrl_plane_bonding,
		hd_pmaif_lpbk_en	=>	hd_pmaif_lpbk_en,
		hd_pmaif_pma_dw_tx	=>	hd_pmaif_pma_dw_tx,
		hd_pmaif_prot_mode_tx	=>	hd_pmaif_prot_mode_tx,
		hd_pmaif_sim_mode	=>	hd_pmaif_sim_mode,
		hd_pmaif_sup_mode	=>	hd_pmaif_sup_mode,
		pcs_tx_clk_out_sel	=>	pcs_tx_clk_out_sel,
		pcs_tx_clk_source	=>	pcs_tx_clk_source,
		pcs_tx_data_source	=>	pcs_tx_data_source,
		pcs_tx_delay1_clk_en	=>	pcs_tx_delay1_clk_en,
		pcs_tx_delay1_clk_sel	=>	pcs_tx_delay1_clk_sel,
		pcs_tx_delay1_ctrl	=>	pcs_tx_delay1_ctrl,
		pcs_tx_delay1_data_sel	=>	pcs_tx_delay1_data_sel,
		pcs_tx_delay2_clk_en	=>	pcs_tx_delay2_clk_en,
		pcs_tx_delay2_ctrl	=>	pcs_tx_delay2_ctrl,
		pcs_tx_output_sel	=>	pcs_tx_output_sel,
		reconfig_settings	=>	reconfig_settings,
		silicon_rev	=>	silicon_rev
	)
	port map (
		-- Instance ports
		avmmaddress	=>	avmmaddress,
		avmmclk	=>	avmmclk,
		avmmread	=>	avmmread,
		avmmrstn	=>	avmmrstn,
		avmmwrite	=>	avmmwrite,
		avmmwritedata	=>	avmmwritedata,
		hip_tx_data	=>	hip_tx_data,
		int_pldif_10g_tx_burst_en_exe	=>	int_pldif_10g_tx_burst_en_exe,
		int_pldif_10g_tx_clk_out	=>	int_pldif_10g_tx_clk_out,
		int_pldif_10g_tx_clk_out_pld_if	=>	int_pldif_10g_tx_clk_out_pld_if,
		int_pldif_10g_tx_empty	=>	int_pldif_10g_tx_empty,
		int_pldif_10g_tx_fifo_num	=>	int_pldif_10g_tx_fifo_num,
		int_pldif_10g_tx_frame	=>	int_pldif_10g_tx_frame,
		int_pldif_10g_tx_full	=>	int_pldif_10g_tx_full,
		int_pldif_10g_tx_pempty	=>	int_pldif_10g_tx_pempty,
		int_pldif_10g_tx_pfull	=>	int_pldif_10g_tx_pfull,
		int_pldif_10g_tx_wordslip_exe	=>	int_pldif_10g_tx_wordslip_exe,
		int_pldif_8g_empty_tx	=>	int_pldif_8g_empty_tx,
		int_pldif_8g_full_tx	=>	int_pldif_8g_full_tx,
		int_pldif_8g_tx_clk_out	=>	int_pldif_8g_tx_clk_out,
		int_pldif_8g_tx_clk_out_pld_if	=>	int_pldif_8g_tx_clk_out_pld_if,
		int_pldif_krfec_tx_alignment	=>	int_pldif_krfec_tx_alignment,
		int_pldif_krfec_tx_frame	=>	int_pldif_krfec_tx_frame,
		int_pldif_pmaif_clkdiv_tx	=>	int_pldif_pmaif_clkdiv_tx,
		int_pldif_pmaif_clkdiv_tx_user	=>	int_pldif_pmaif_clkdiv_tx_user,
		int_pldif_pmaif_uhsif_tx_clk_out	=>	int_pldif_pmaif_uhsif_tx_clk_out,
		pld_10g_krfec_tx_pld_rst_n	=>	pld_10g_krfec_tx_pld_rst_n,
		pld_10g_tx_bitslip	=>	pld_10g_tx_bitslip,
		pld_10g_tx_burst_en	=>	pld_10g_tx_burst_en,
		pld_10g_tx_data_valid	=>	pld_10g_tx_data_valid,
		pld_10g_tx_diag_status	=>	pld_10g_tx_diag_status,
		pld_10g_tx_wordslip	=>	pld_10g_tx_wordslip,
		pld_8g_g3_tx_pld_rst_n	=>	pld_8g_g3_tx_pld_rst_n,
		pld_8g_rddisable_tx	=>	pld_8g_rddisable_tx,
		pld_8g_tx_boundary_sel	=>	pld_8g_tx_boundary_sel,
		pld_8g_wrenable_tx	=>	pld_8g_wrenable_tx,
		pld_partial_reconfig	=>	pld_partial_reconfig,
		pld_pma_txpma_rstb	=>	pld_pma_txpma_rstb,
		pld_pmaif_tx_pld_rst_n	=>	pld_pmaif_tx_pld_rst_n,
		pld_polinv_tx	=>	pld_polinv_tx,
		pld_tx_clk	=>	pld_tx_clk,
		pld_tx_control	=>	pld_tx_control,
		pld_tx_data	=>	pld_tx_data,
		pld_txelecidle	=>	pld_txelecidle,
		pld_uhsif_tx_clk	=>	pld_uhsif_tx_clk,
		scan_mode_n	=>	scan_mode_n,
		avmmreaddata	=>	avmmreaddata,
		blockselect	=>	blockselect,
		hip_clk_out_div_by_2_wire	=>	hip_clk_out_div_by_2_wire,
		hip_clk_out_wire	=>	hip_clk_out_wire,
		pld_10g_tx_burst_en_exe_10g_fastreg	=>	pld_10g_tx_burst_en_exe_10g_fastreg,
		pld_10g_tx_burst_en_exe_plddirect_reg	=>	pld_10g_tx_burst_en_exe_plddirect_reg,
		pld_10g_tx_data_valid_2ff_delay1_fastreg	=>	pld_10g_tx_data_valid_2ff_delay1_fastreg,
		pld_10g_tx_data_valid_2ff_delay3_fastreg	=>	pld_10g_tx_data_valid_2ff_delay3_fastreg,
		pld_10g_tx_data_valid_2ff_delay4_fastreg	=>	pld_10g_tx_data_valid_2ff_delay4_fastreg,
		pld_10g_tx_data_valid_2ff_delay4_plddirect_fastreg	=>	pld_10g_tx_data_valid_2ff_delay4_plddirect_fastreg,
		pld_10g_tx_data_valid_2ff_delay6_fastreg	=>	pld_10g_tx_data_valid_2ff_delay6_fastreg,
		pld_10g_tx_data_valid_2ff_delay6_plddirect_fastreg	=>	pld_10g_tx_data_valid_2ff_delay6_plddirect_fastreg,
		pld_10g_tx_data_valid_fastreg	=>	pld_10g_tx_data_valid_fastreg,
		pld_10g_tx_data_valid_plddirect_fastreg	=>	pld_10g_tx_data_valid_plddirect_fastreg,
		pld_pcs_tx_clk_out_pma_wire	=>	pld_pcs_tx_clk_out_pma_wire,
		pld_pma_tx_clk_out_wire	=>	pld_pma_tx_clk_out_wire,
		pld_pmaif_tx_pld_rst_n_reg	=>	pld_pmaif_tx_pld_rst_n_reg,
		pld_polinv_tx_10g_pcsdirect_reg	=>	pld_polinv_tx_10g_pcsdirect_reg,
		pld_polinv_tx_8g_reg	=>	pld_polinv_tx_8g_reg,
		pld_polinv_tx_pat_reg	=>	pld_polinv_tx_pat_reg,
		pld_tx_clk_fifo	=>	pld_tx_clk_fifo,
		pld_tx_control_fifo	=>	pld_tx_control_fifo,
		pld_tx_control_hi_10g_reg	=>	pld_tx_control_hi_10g_reg,
		pld_tx_control_lo_10g_2ff_delay4_fastreg	=>	pld_tx_control_lo_10g_2ff_delay4_fastreg,
		pld_tx_control_lo_10g_2ff_delay6_fastreg	=>	pld_tx_control_lo_10g_2ff_delay6_fastreg,
		pld_tx_control_lo_10g_fastreg	=>	pld_tx_control_lo_10g_fastreg,
		pld_tx_control_lo_8g_2ff_delay4_fastreg	=>	pld_tx_control_lo_8g_2ff_delay4_fastreg,
		pld_tx_control_lo_8g_2ff_delay6_fastreg	=>	pld_tx_control_lo_8g_2ff_delay6_fastreg,
		pld_tx_control_lo_8g_fastreg	=>	pld_tx_control_lo_8g_fastreg,
		pld_tx_control_lo_plddirect_2ff_delay1_fastreg	=>	pld_tx_control_lo_plddirect_2ff_delay1_fastreg,
		pld_tx_control_lo_plddirect_2ff_delay3_fastreg	=>	pld_tx_control_lo_plddirect_2ff_delay3_fastreg,
		pld_tx_control_lo_plddirect_2ff_delay4_fastreg	=>	pld_tx_control_lo_plddirect_2ff_delay4_fastreg,
		pld_tx_control_lo_plddirect_2ff_delay6_fastreg	=>	pld_tx_control_lo_plddirect_2ff_delay6_fastreg,
		pld_tx_control_lo_plddirect_fastreg	=>	pld_tx_control_lo_plddirect_fastreg,
		pld_tx_control_lo_plddirect_reg	=>	pld_tx_control_lo_plddirect_reg,
		pld_tx_data_hi_reg	=>	pld_tx_data_hi_reg,
		pld_tx_data_lo_10g_2ff_delay4_fastreg	=>	pld_tx_data_lo_10g_2ff_delay4_fastreg,
		pld_tx_data_lo_10g_2ff_delay6_fastreg	=>	pld_tx_data_lo_10g_2ff_delay6_fastreg,
		pld_tx_data_lo_10g_fastreg	=>	pld_tx_data_lo_10g_fastreg,
		pld_tx_data_lo_8g_2ff_delay4_fastreg	=>	pld_tx_data_lo_8g_2ff_delay4_fastreg,
		pld_tx_data_lo_8g_2ff_delay6_fastreg	=>	pld_tx_data_lo_8g_2ff_delay6_fastreg,
		pld_tx_data_lo_8g_fastreg	=>	pld_tx_data_lo_8g_fastreg,
		pld_tx_data_lo_plddirect_2ff_delay1_fastreg	=>	pld_tx_data_lo_plddirect_2ff_delay1_fastreg,
		pld_tx_data_lo_plddirect_2ff_delay3_fastreg	=>	pld_tx_data_lo_plddirect_2ff_delay3_fastreg,
		pld_tx_data_lo_plddirect_2ff_delay4_fastreg	=>	pld_tx_data_lo_plddirect_2ff_delay4_fastreg,
		pld_tx_data_lo_plddirect_2ff_delay6_fastreg	=>	pld_tx_data_lo_plddirect_2ff_delay6_fastreg,
		pld_tx_data_lo_plddirect_fastreg	=>	pld_tx_data_lo_plddirect_fastreg,
		pld_tx_data_lo_plddirect_reg	=>	pld_tx_data_lo_plddirect_reg,
		pld_uhsif_reg	=>	pld_uhsif_reg,
		pma_tx_pma_clk_reg	=>	pma_tx_pma_clk_reg,
		hip_tx_clk	=>	hip_tx_clk,
		int_pldif_10g_tx_bitslip	=>	int_pldif_10g_tx_bitslip,
		int_pldif_10g_tx_burst_en	=>	int_pldif_10g_tx_burst_en,
		int_pldif_10g_tx_control	=>	int_pldif_10g_tx_control,
		int_pldif_10g_tx_control_reg	=>	int_pldif_10g_tx_control_reg,
		int_pldif_10g_tx_data	=>	int_pldif_10g_tx_data,
		int_pldif_10g_tx_data_reg	=>	int_pldif_10g_tx_data_reg,
		int_pldif_10g_tx_data_valid	=>	int_pldif_10g_tx_data_valid,
		int_pldif_10g_tx_data_valid_reg	=>	int_pldif_10g_tx_data_valid_reg,
		int_pldif_10g_tx_diag_status	=>	int_pldif_10g_tx_diag_status,
		int_pldif_10g_tx_pld_clk	=>	int_pldif_10g_tx_pld_clk,
		int_pldif_10g_tx_pld_rst_n	=>	int_pldif_10g_tx_pld_rst_n,
		int_pldif_10g_tx_wordslip	=>	int_pldif_10g_tx_wordslip,
		int_pldif_8g_pld_tx_clk	=>	int_pldif_8g_pld_tx_clk,
		int_pldif_8g_powerdown	=>	int_pldif_8g_powerdown,
		int_pldif_8g_rddisable_tx	=>	int_pldif_8g_rddisable_tx,
		int_pldif_8g_rev_loopbk	=>	int_pldif_8g_rev_loopbk,
		int_pldif_8g_tx_blk_start	=>	int_pldif_8g_tx_blk_start,
		int_pldif_8g_tx_boundary_sel	=>	int_pldif_8g_tx_boundary_sel,
		int_pldif_8g_tx_data_valid	=>	int_pldif_8g_tx_data_valid,
		int_pldif_8g_tx_sync_hdr	=>	int_pldif_8g_tx_sync_hdr,
		int_pldif_8g_txd	=>	int_pldif_8g_txd,
		int_pldif_8g_txd_fast_reg	=>	int_pldif_8g_txd_fast_reg,
		int_pldif_8g_txdeemph	=>	int_pldif_8g_txdeemph,
		int_pldif_8g_txdetectrxloopback	=>	int_pldif_8g_txdetectrxloopback,
		int_pldif_8g_txelecidle	=>	int_pldif_8g_txelecidle,
		int_pldif_8g_txmargin	=>	int_pldif_8g_txmargin,
		int_pldif_8g_txswing	=>	int_pldif_8g_txswing,
		int_pldif_8g_txurstpcs_n	=>	int_pldif_8g_txurstpcs_n,
		int_pldif_8g_wrenable_tx	=>	int_pldif_8g_wrenable_tx,
		int_pldif_pmaif_8g_txurstpcs_n	=>	int_pldif_pmaif_8g_txurstpcs_n,
		int_pldif_pmaif_polinv_tx	=>	int_pldif_pmaif_polinv_tx,
		int_pldif_pmaif_tx_data	=>	int_pldif_pmaif_tx_data,
		int_pldif_pmaif_tx_pld_clk	=>	int_pldif_pmaif_tx_pld_clk,
		int_pldif_pmaif_tx_pld_rst_n	=>	int_pldif_pmaif_tx_pld_rst_n,
		int_pldif_pmaif_txelecidle	=>	int_pldif_pmaif_txelecidle,
		int_pldif_pmaif_txpma_rstb	=>	int_pldif_pmaif_txpma_rstb,
		int_pldif_pmaif_uhsif_tx_clk	=>	int_pldif_pmaif_uhsif_tx_clk,
		int_pldif_pmaif_uhsif_tx_data	=>	int_pldif_pmaif_uhsif_tx_data,
		pld_10g_krfec_tx_frame	=>	pld_10g_krfec_tx_frame,
		pld_10g_tx_burst_en_exe	=>	pld_10g_tx_burst_en_exe,
		pld_10g_tx_empty	=>	pld_10g_tx_empty,
		pld_10g_tx_fifo_num	=>	pld_10g_tx_fifo_num,
		pld_10g_tx_full	=>	pld_10g_tx_full,
		pld_10g_tx_pempty	=>	pld_10g_tx_pempty,
		pld_10g_tx_pfull	=>	pld_10g_tx_pfull,
		pld_10g_tx_wordslip_exe	=>	pld_10g_tx_wordslip_exe,
		pld_8g_empty_tx	=>	pld_8g_empty_tx,
		pld_8g_full_tx	=>	pld_8g_full_tx,
		pld_krfec_tx_alignment	=>	pld_krfec_tx_alignment,
		pld_pcs_tx_clk_out	=>	pld_pcs_tx_clk_out,
		pld_pma_clkdiv_tx_user	=>	pld_pma_clkdiv_tx_user,
		pld_pma_tx_clk_out	=>	pld_pma_tx_clk_out,
		pld_uhsif_tx_clk_out	=>	pld_uhsif_tx_clk_out
	);

end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HSSI_COMPONENTS.all;


entity	twentynm_hssi_avmm_if	is
	generic	(
		silicon_rev	:	string	:=	"reve";
		calibration_en	:	string	:=	"enable";
		arbiter_ctrl	:	string	:=	"uc";
		cal_done	:	string	:=	"cal_done_assert";
		hip_cal_en	:	string	:=	"disable";
		cal_reserved	:	bit_vector	:=	B"00000";
		calibration_type	:	string	:=	"one_time"
	);
	port	(
		avmmclk	:	in	std_logic	:= '0';
		avmmwrite	:	in	std_logic	:= '0';
		avmmread	:	in	std_logic	:= '0';
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:= "000000000";
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:= "00000000";
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:= "00000000";
		avmmrequest	:	in	std_logic	:= '0';
		avmmbusy	:	out	std_logic	:= '0';
		hipcaldone	:	out	std_logic	:= '0';
		pldcaldone	:	out	std_logic	:= '0';
		clkchnl	:	out	std_logic	:= '0';
		rstnchnl	:	out	std_logic	:= '0';
		writedatachnl	:	out	std_logic_vector(7 downto 0)	:= "00000000";
		regaddrchnl	:	out	std_logic_vector(8 downto 0)	:= "000000000";
		writechnl	:	out	std_logic	:= '0';
		readchnl	:	out	std_logic	:= '0';
		blockselect	:	in	std_logic_vector(69 downto 0)	:= "0000000000000000000000000000000000000000000000000000000000000000000000";
		readdatachnl	:	in	std_logic_vector(559 downto 0)	:= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		avmmrstn	:	in	std_logic	:= '0';
		scanmoden	:	in	std_logic	:= '0';
		scanshiftn	:	in	std_logic	:= '0';
		avmmreservedin	:	in	std_logic	:= '0';
		avmmreservedout	:	out		std_logic	:= '0'
	);
end	twentynm_hssi_avmm_if;

architecture behavior of twentynm_hssi_avmm_if is

constant cal_reserved_int        :       integer :=      bin2int(cal_reserved);
component	twentynm_hssi_avmm_if_encrypted
	generic
	(
		silicon_rev	:	string	:=	"reve";
		calibration_en	:	string	:=	"enable";
		arbiter_ctrl	:	string	:=	"uc";
		cal_done	:	string	:=	"cal_done_assert";
		hip_cal_en	:	string	:=	"disable";
		cal_reserved	:	integer	:=	0;
		calibration_type	:	string	:=	"one_time"
	);
	port	(
		avmmclk	:	in	std_logic	:= '0';
		avmmwrite	:	in	std_logic	:= '0';
		avmmread	:	in	std_logic	:= '0';
		avmmaddress	:	in	std_logic_vector(8 downto 0)	:= "000000000";
		avmmwritedata	:	in	std_logic_vector(7 downto 0)	:= "00000000";
		avmmreaddata	:	out	std_logic_vector(7 downto 0)	:= "00000000";
		avmmrequest	:	in	std_logic	:= '0';
		avmmbusy	:	out	std_logic	:= '0';
		hipcaldone	:	out	std_logic	:= '0';
		pldcaldone	:	out	std_logic	:= '0';
		clkchnl	:	out	std_logic	:= '0';
		rstnchnl	:	out	std_logic	:= '0';
		writedatachnl	:	out	std_logic_vector(7 downto 0)	:= "00000000";
		regaddrchnl	:	out	std_logic_vector(8 downto 0)	:= "000000000";
		writechnl	:	out	std_logic	:= '0';
		readchnl	:	out	std_logic	:= '0';
		blockselect	:	in	std_logic_vector(69 downto 0)	:= "0000000000000000000000000000000000000000000000000000000000000000000000";
		readdatachnl	:	in	std_logic_vector(559 downto 0)	:= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		avmmrstn	:	in	std_logic	:= '0';
		scanmoden	:	in	std_logic	:= '0';
		scanshiftn	:	in	std_logic	:= '0';
		avmmreservedin	:	in	std_logic	:= '0';
		avmmreservedout	:	out		std_logic	:= '0'
	);
end component;

begin


inst : twentynm_hssi_avmm_if_encrypted
	generic map	(
		silicon_rev	=>	silicon_rev,
		calibration_en	=>	calibration_en,
		arbiter_ctrl	=>	arbiter_ctrl,
		cal_done	=>	cal_done,
		hip_cal_en	=>	hip_cal_en,
		cal_reserved	=>	cal_reserved_int,
		calibration_type	=>	calibration_type
	)
	port map	(
		avmmclk	=>	avmmclk,
		avmmwrite	=>	avmmwrite,
		avmmread	=>	avmmread,
		avmmaddress	=>	avmmaddress,
		avmmwritedata	=>	avmmwritedata,
		avmmreaddata	=>	avmmreaddata,
		avmmrequest	=>	avmmrequest,
		avmmbusy	=>	avmmbusy,
		hipcaldone	=>	hipcaldone,
		pldcaldone	=>	pldcaldone,
		clkchnl	=>	clkchnl,
		rstnchnl	=>	rstnchnl,
		writedatachnl	=>	writedatachnl,
		regaddrchnl	=>	regaddrchnl,
		writechnl	=>	writechnl,
		readchnl	=>	readchnl,
		blockselect	=>	blockselect,
		readdatachnl	=>	readdatachnl,
		avmmrstn	=>	avmmrstn,
		scanmoden	=>	scanmoden,
		scanshiftn	=>	scanshiftn,
		avmmreservedin	=>	avmmreservedin,
		avmmreservedout	=>	avmmreservedout
	);


end behavior;

