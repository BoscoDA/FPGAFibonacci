-- Copyright (C) 2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, the Intel Quartus Prime License Agreement, the Intel
-- MegaCore Function License Agreement, or other applicable 
-- license agreement, including, without limitation, that your
-- use is for the sole purpose of simulating designs for use 
-- exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- Quartus Prime 17.0.1 Build 598 06/07/2017

LIBRARY IEEE;
use IEEE.STD_LOGIC_1164.all;

package TWENTYNM_HIP_COMPONENTS is

-- GENERIC utility functions BEGIN
function bin2int (s : std_logic_vector) return integer;
function bin2int (s : bit_vector) return integer;
function bin2int (s : std_logic) return integer;
function bin2int (s : bit) return integer;
function int2bit (arg : boolean) return std_logic;
function str2bin (s : string) return std_logic_vector;
function str2int (s : string) return integer;
function int2bin (arg : integer; size : integer) return std_logic_vector;
function int2bin (arg : boolean; size : integer) return std_logic_vector;
function int2bit (arg : integer) return std_logic;

component	twentynm_hssi_gen3_x8_pcie_hip
	generic (
		-- Architecture parameters
		acknack_base	:	bit_vector	:=	B"0000000000000";
		acknack_set	:	string	:=	"false";
		advance_error_reporting	:	string	:=	"disable";
		app_interface_width	:	string	:=	"avst_64bit";
		arb_upfc_30us_counter	:	bit_vector	:=	B"0000";
		arb_upfc_30us_en	:	string	:=	"enable";
		aspm_config_management	:	string	:=	"true";
		aspm_patch_disable	:	string	:=	"enable_both";
		ast_width_rx	:	string	:=	"rx_64";
		ast_width_tx	:	string	:=	"tx_64";
		atomic_malformed	:	string	:=	"false";
		atomic_op_completer_32bit	:	string	:=	"false";
		atomic_op_completer_64bit	:	string	:=	"false";
		atomic_op_routing	:	string	:=	"false";
		auto_msg_drop_enable	:	string	:=	"false";
		avmm_cvp_inter_sel_csr_ctrl	:	string	:=	"disable";
		avmm_dprio_broadcast_en_csr_ctrl	:	string	:=	"disable";
		avmm_force_inter_sel_csr_ctrl	:	string	:=	"disable";
		avmm_power_iso_en_csr_ctrl	:	string	:=	"disable";
		bar0_size_mask	:	bit_vector	:=	B"1111111111111111111111111111";
		bar0_type	:	string	:=	"bar0_64bit_prefetch_mem";
		bar1_size_mask	:	bit_vector	:=	B"0000000000000000000000000000";
		bar1_type	:	string	:=	"bar1_disable";
		bar2_size_mask	:	bit_vector	:=	B"0000000000000000000000000000";
		bar2_type	:	string	:=	"bar2_disable";
		bar3_size_mask	:	bit_vector	:=	B"0000000000000000000000000000";
		bar3_type	:	string	:=	"bar3_disable";
		bar4_size_mask	:	bit_vector	:=	B"0000000000000000000000000000";
		bar4_type	:	string	:=	"bar4_disable";
		bar5_size_mask	:	bit_vector	:=	B"0000000000000000000000000000";
		bar5_type	:	string	:=	"bar5_disable";
		base_counter_sel	:	string	:=	"count_clk_62p5";
		bist_memory_settings	:	string	:=	"000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		bridge_port_ssid_support	:	string	:=	"false";
		bridge_port_vga_enable	:	string	:=	"false";
		bypass_cdc	:	string	:=	"false";
		bypass_clk_switch	:	string	:=	"false";
		bypass_tl	:	string	:=	"false";
		capab_rate_rxcfg_en	:	string	:=	"disable";
		cas_completer_128bit	:	string	:=	"false";
		cdc_clk_relation	:	string	:=	"plesiochronous";
		cdc_dummy_insert_limit	:	bit_vector	:=	B"1011";
		cfg_parchk_ena	:	string	:=	"disable";
		cfgbp_req_recov_disable	:	string	:=	"false";
		class_code	:	bit_vector	:=	B"111111110000000000000000";
		clock_pwr_management	:	string	:=	"false";
		completion_timeout	:	string	:=	"abcd";
		core_clk_divider	:	string	:=	"div_1";
		core_clk_freq_mhz	:	string	:=	"core_clk_250mhz";
		core_clk_out_sel	:	string	:=	"core_clk_out_div_1";
		core_clk_sel	:	string	:=	"pld_clk";
		core_clk_source	:	string	:=	"pll_fixed_clk";
		cseb_bar_match_checking	:	string	:=	"enable";
		cseb_config_bypass	:	string	:=	"disable";
		cseb_cpl_status_during_cvp	:	string	:=	"completer_abort";
		cseb_cpl_tag_checking	:	string	:=	"enable";
		cseb_disable_auto_crs	:	string	:=	"false";
		cseb_extend_pci	:	string	:=	"false";
		cseb_extend_pcie	:	string	:=	"false";
		cseb_min_error_checking	:	string	:=	"false";
		cseb_route_to_avl_rx_st	:	string	:=	"cseb";
		cseb_temp_busy_crs	:	string	:=	"completer_abort_tmp_busy";
		cvp_clk_reset	:	string	:=	"false";
		cvp_data_compressed	:	string	:=	"false";
		cvp_data_encrypted	:	string	:=	"false";
		cvp_enable	:	string	:=	"cvp_dis";
		cvp_mode_reset	:	string	:=	"false";
		cvp_rate_sel	:	string	:=	"full_rate";
		d0_pme	:	string	:=	"false";
		d1_pme	:	string	:=	"false";
		d1_support	:	string	:=	"false";
		d2_pme	:	string	:=	"false";
		d2_support	:	string	:=	"false";
		d3_cold_pme	:	string	:=	"false";
		d3_hot_pme	:	string	:=	"false";
		data_pack_rx	:	string	:=	"disable";
		deemphasis_enable	:	string	:=	"false";
		deskew_comma	:	string	:=	"skp_eieos_deskw";
		device_id	:	bit_vector	:=	B"1110000000000001";
		device_number	:	bit_vector	:=	B"00000";
		device_specific_init	:	string	:=	"false";
		dft_clock_obsrv_en	:	string	:=	"disable";
		dft_clock_obsrv_sel	:	string	:=	"dft_pclk";
		diffclock_nfts_count	:	bit_vector	:=	B"00000000";
		dis_cplovf	:	string	:=	"disable";
		dis_paritychk	:	string	:=	"enable";
		disable_link_x2_support	:	string	:=	"false";
		disable_snoop_packet	:	string	:=	"false";
		dl_tx_check_parity_edb	:	string	:=	"disable";
		dll_active_report_support	:	string	:=	"false";
		early_dl_up	:	string	:=	"true";
		eco_fb332688_dis	:	string	:=	"true";
		ecrc_check_capable	:	string	:=	"true";
		ecrc_gen_capable	:	string	:=	"true";
		egress_block_err_report_ena	:	string	:=	"false";
		ei_delay_powerdown_count	:	bit_vector	:=	B"00001010";
		eie_before_nfts_count	:	bit_vector	:=	B"0100";
		electromech_interlock	:	string	:=	"false";
		en_ieiupdatefc	:	string	:=	"false";
		en_lane_errchk	:	string	:=	"false";
		en_phystatus_dly	:	string	:=	"false";
		ena_ido_cpl	:	string	:=	"false";
		ena_ido_req	:	string	:=	"false";
		enable_adapter_half_rate_mode	:	string	:=	"false";
		enable_ch01_pclk_out	:	string	:=	"pclk_ch0";
		enable_ch0_pclk_out	:	string	:=	"pclk_ch01";
		enable_completion_timeout_disable	:	string	:=	"true";
		enable_directed_spd_chng	:	string	:=	"false";
		enable_function_msix_support	:	string	:=	"true";
		enable_l0s_aspm	:	string	:=	"false";
		enable_l1_aspm	:	string	:=	"false";
		enable_rx_buffer_checking	:	string	:=	"false";
		enable_rx_reordering	:	string	:=	"true";
		enable_slot_register	:	string	:=	"false";
		endpoint_l0_latency	:	bit_vector	:=	B"000";
		endpoint_l1_latency	:	bit_vector	:=	B"000";
		eql_rq_int_en_number	:	bit_vector	:=	B"000000";
		errmgt_fcpe_patch_dis	:	string	:=	"enable";
		errmgt_fep_patch_dis	:	string	:=	"enable";
		expansion_base_address_register	:	string	:=	"00000000000000000000000000000000";
		extend_tag_field	:	string	:=	"false";
		extended_format_field	:	string	:=	"true";
		extended_tag_reset	:	string	:=	"false";
		fc_init_timer	:	bit_vector	:=	B"10000000000";
		flow_control_timeout_count	:	bit_vector	:=	B"11001000";
		flow_control_update_count	:	bit_vector	:=	B"11110";
		flr_capability	:	string	:=	"true";
		force_dis_to_det	:	string	:=	"false";
		force_gen1_dis	:	string	:=	"false";
		force_tx_coeff_preset_lpbk	:	string	:=	"false";
		frame_err_patch_dis	:	string	:=	"enable";
		func_mode	:	string	:=	"disable";
		g3_bypass_equlz	:	string	:=	"false";
		g3_coeff_done_tmout	:	string	:=	"enable";
		g3_deskew_char	:	string	:=	"default_sdsos";
		g3_dis_be_frm_err	:	string	:=	"false";
		g3_dn_rx_hint_eqlz_0	:	bit_vector	:=	B"000";
		g3_dn_rx_hint_eqlz_1	:	bit_vector	:=	B"000";
		g3_dn_rx_hint_eqlz_2	:	bit_vector	:=	B"000";
		g3_dn_rx_hint_eqlz_3	:	bit_vector	:=	B"000";
		g3_dn_rx_hint_eqlz_4	:	bit_vector	:=	B"000";
		g3_dn_rx_hint_eqlz_5	:	bit_vector	:=	B"000";
		g3_dn_rx_hint_eqlz_6	:	bit_vector	:=	B"000";
		g3_dn_rx_hint_eqlz_7	:	bit_vector	:=	B"000";
		g3_dn_tx_preset_eqlz_0	:	bit_vector	:=	B"0000";
		g3_dn_tx_preset_eqlz_1	:	bit_vector	:=	B"0000";
		g3_dn_tx_preset_eqlz_2	:	bit_vector	:=	B"0000";
		g3_dn_tx_preset_eqlz_3	:	bit_vector	:=	B"0000";
		g3_dn_tx_preset_eqlz_4	:	bit_vector	:=	B"0000";
		g3_dn_tx_preset_eqlz_5	:	bit_vector	:=	B"0000";
		g3_dn_tx_preset_eqlz_6	:	bit_vector	:=	B"0000";
		g3_dn_tx_preset_eqlz_7	:	bit_vector	:=	B"0000";
		g3_force_ber_max	:	string	:=	"false";
		g3_force_ber_min	:	string	:=	"false";
		g3_lnk_trn_rx_ts	:	string	:=	"false";
		g3_ltssm_eq_dbg	:	string	:=	"false";
		g3_ltssm_rec_dbg	:	string	:=	"false";
		g3_pause_ltssm_rec_en	:	string	:=	"disable";
		g3_quiesce_guarant	:	string	:=	"false";
		g3_redo_equlz_dis	:	string	:=	"false";
		g3_redo_equlz_en	:	string	:=	"false";
		g3_up_rx_hint_eqlz_0	:	bit_vector	:=	B"000";
		g3_up_rx_hint_eqlz_1	:	bit_vector	:=	B"000";
		g3_up_rx_hint_eqlz_2	:	bit_vector	:=	B"000";
		g3_up_rx_hint_eqlz_3	:	bit_vector	:=	B"000";
		g3_up_rx_hint_eqlz_4	:	bit_vector	:=	B"000";
		g3_up_rx_hint_eqlz_5	:	bit_vector	:=	B"000";
		g3_up_rx_hint_eqlz_6	:	bit_vector	:=	B"000";
		g3_up_rx_hint_eqlz_7	:	bit_vector	:=	B"000";
		g3_up_tx_preset_eqlz_0	:	bit_vector	:=	B"0000";
		g3_up_tx_preset_eqlz_1	:	bit_vector	:=	B"0000";
		g3_up_tx_preset_eqlz_2	:	bit_vector	:=	B"0000";
		g3_up_tx_preset_eqlz_3	:	bit_vector	:=	B"0000";
		g3_up_tx_preset_eqlz_4	:	bit_vector	:=	B"0000";
		g3_up_tx_preset_eqlz_5	:	bit_vector	:=	B"0000";
		g3_up_tx_preset_eqlz_6	:	bit_vector	:=	B"0000";
		g3_up_tx_preset_eqlz_7	:	bit_vector	:=	B"0000";
		gen123_lane_rate_mode	:	string	:=	"gen1_rate";
		gen2_diffclock_nfts_count	:	bit_vector	:=	B"11111111";
		gen2_pma_pll_usage	:	string	:=	"not_applicaple";
		gen2_sameclock_nfts_count	:	bit_vector	:=	B"11111111";
		gen3_coeff_1	:	bit_vector	:=	B"000000000000000100";
		gen3_coeff_10	:	bit_vector	:=	B"000000000000000111";
		gen3_coeff_10_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_10_nxtber_less	:	bit_vector	:=	B"1111";
		gen3_coeff_10_nxtber_more	:	bit_vector	:=	B"1010";
		gen3_coeff_10_preset_hint	:	bit_vector	:=	B"011";
		gen3_coeff_10_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_10_sel	:	string	:=	"preset_10";
		gen3_coeff_11	:	bit_vector	:=	B"000000000000000111";
		gen3_coeff_11_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_11_nxtber_less	:	bit_vector	:=	B"1111";
		gen3_coeff_11_nxtber_more	:	bit_vector	:=	B"1111";
		gen3_coeff_11_preset_hint	:	bit_vector	:=	B"100";
		gen3_coeff_11_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_11_sel	:	string	:=	"preset_11";
		gen3_coeff_12	:	bit_vector	:=	B"000000000000000111";
		gen3_coeff_12_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_12_nxtber_less	:	bit_vector	:=	B"1111";
		gen3_coeff_12_nxtber_more	:	bit_vector	:=	B"1111";
		gen3_coeff_12_preset_hint	:	bit_vector	:=	B"010";
		gen3_coeff_12_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_12_sel	:	string	:=	"preset_12";
		gen3_coeff_13	:	bit_vector	:=	B"000000000000000100";
		gen3_coeff_13_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_13_nxtber_less	:	bit_vector	:=	B"1101";
		gen3_coeff_13_nxtber_more	:	bit_vector	:=	B"0001";
		gen3_coeff_13_preset_hint	:	bit_vector	:=	B"100";
		gen3_coeff_13_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_13_sel	:	string	:=	"preset_13";
		gen3_coeff_14	:	bit_vector	:=	B"000000000000000100";
		gen3_coeff_14_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_14_nxtber_less	:	bit_vector	:=	B"1111";
		gen3_coeff_14_nxtber_more	:	bit_vector	:=	B"0010";
		gen3_coeff_14_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_14_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_14_sel	:	string	:=	"preset_14";
		gen3_coeff_15	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_15_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_15_nxtber_less	:	bit_vector	:=	B"0000";
		gen3_coeff_15_nxtber_more	:	bit_vector	:=	B"0000";
		gen3_coeff_15_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_15_reqber	:	bit_vector	:=	B"00000";
		gen3_coeff_15_sel	:	string	:=	"coeff_15";
		gen3_coeff_16	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_16_ber_meas	:	bit_vector	:=	B"000000";
		gen3_coeff_16_nxtber_less	:	bit_vector	:=	B"0000";
		gen3_coeff_16_nxtber_more	:	bit_vector	:=	B"0000";
		gen3_coeff_16_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_16_reqber	:	bit_vector	:=	B"00000";
		gen3_coeff_16_sel	:	string	:=	"coeff_16";
		gen3_coeff_17	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_17_ber_meas	:	bit_vector	:=	B"000000";
		gen3_coeff_17_nxtber_less	:	bit_vector	:=	B"0000";
		gen3_coeff_17_nxtber_more	:	bit_vector	:=	B"0000";
		gen3_coeff_17_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_17_reqber	:	bit_vector	:=	B"00000";
		gen3_coeff_17_sel	:	string	:=	"coeff_17";
		gen3_coeff_18	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_18_ber_meas	:	bit_vector	:=	B"000000";
		gen3_coeff_18_nxtber_less	:	bit_vector	:=	B"0000";
		gen3_coeff_18_nxtber_more	:	bit_vector	:=	B"0000";
		gen3_coeff_18_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_18_reqber	:	bit_vector	:=	B"00000";
		gen3_coeff_18_sel	:	string	:=	"coeff_18";
		gen3_coeff_19	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_19_ber_meas	:	bit_vector	:=	B"000000";
		gen3_coeff_19_nxtber_less	:	bit_vector	:=	B"0000";
		gen3_coeff_19_nxtber_more	:	bit_vector	:=	B"0000";
		gen3_coeff_19_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_19_reqber	:	bit_vector	:=	B"00000";
		gen3_coeff_19_sel	:	string	:=	"coeff_19";
		gen3_coeff_1_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_1_nxtber_less	:	bit_vector	:=	B"1100";
		gen3_coeff_1_nxtber_more	:	bit_vector	:=	B"0110";
		gen3_coeff_1_preset_hint	:	bit_vector	:=	B"010";
		gen3_coeff_1_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_1_sel	:	string	:=	"preset_1";
		gen3_coeff_2	:	bit_vector	:=	B"000000000000000001";
		gen3_coeff_20	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_20_ber_meas	:	bit_vector	:=	B"000000";
		gen3_coeff_20_nxtber_less	:	bit_vector	:=	B"0000";
		gen3_coeff_20_nxtber_more	:	bit_vector	:=	B"0000";
		gen3_coeff_20_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_20_reqber	:	bit_vector	:=	B"00000";
		gen3_coeff_20_sel	:	string	:=	"coeff_20";
		gen3_coeff_21	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_21_ber_meas	:	bit_vector	:=	B"000000";
		gen3_coeff_21_nxtber_less	:	bit_vector	:=	B"0000";
		gen3_coeff_21_nxtber_more	:	bit_vector	:=	B"0000";
		gen3_coeff_21_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_21_reqber	:	bit_vector	:=	B"00000";
		gen3_coeff_21_sel	:	string	:=	"coeff_21";
		gen3_coeff_22	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_22_ber_meas	:	bit_vector	:=	B"000000";
		gen3_coeff_22_nxtber_less	:	bit_vector	:=	B"0000";
		gen3_coeff_22_nxtber_more	:	bit_vector	:=	B"0000";
		gen3_coeff_22_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_22_reqber	:	bit_vector	:=	B"00000";
		gen3_coeff_22_sel	:	string	:=	"coeff_22";
		gen3_coeff_23	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_23_ber_meas	:	bit_vector	:=	B"000000";
		gen3_coeff_23_nxtber_less	:	bit_vector	:=	B"0000";
		gen3_coeff_23_nxtber_more	:	bit_vector	:=	B"0000";
		gen3_coeff_23_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_23_reqber	:	bit_vector	:=	B"00000";
		gen3_coeff_23_sel	:	string	:=	"coeff_23";
		gen3_coeff_24	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_24_ber_meas	:	bit_vector	:=	B"000000";
		gen3_coeff_24_nxtber_less	:	bit_vector	:=	B"0000";
		gen3_coeff_24_nxtber_more	:	bit_vector	:=	B"0000";
		gen3_coeff_24_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_24_reqber	:	bit_vector	:=	B"00000";
		gen3_coeff_24_sel	:	string	:=	"coeff_24";
		gen3_coeff_2_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_2_nxtber_less	:	bit_vector	:=	B"0010";
		gen3_coeff_2_nxtber_more	:	bit_vector	:=	B"0100";
		gen3_coeff_2_preset_hint	:	bit_vector	:=	B"100";
		gen3_coeff_2_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_2_sel	:	string	:=	"preset_2";
		gen3_coeff_3	:	bit_vector	:=	B"000000000000000001";
		gen3_coeff_3_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_3_nxtber_less	:	bit_vector	:=	B"1111";
		gen3_coeff_3_nxtber_more	:	bit_vector	:=	B"0011";
		gen3_coeff_3_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_3_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_3_sel	:	string	:=	"preset_3";
		gen3_coeff_4	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_4_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_4_nxtber_less	:	bit_vector	:=	B"1111";
		gen3_coeff_4_nxtber_more	:	bit_vector	:=	B"0100";
		gen3_coeff_4_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_4_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_4_sel	:	string	:=	"preset_4";
		gen3_coeff_5	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_5_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_5_nxtber_less	:	bit_vector	:=	B"1111";
		gen3_coeff_5_nxtber_more	:	bit_vector	:=	B"0101";
		gen3_coeff_5_preset_hint	:	bit_vector	:=	B"100";
		gen3_coeff_5_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_5_sel	:	string	:=	"preset_5";
		gen3_coeff_6	:	bit_vector	:=	B"000000000000000111";
		gen3_coeff_6_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_6_nxtber_less	:	bit_vector	:=	B"1111";
		gen3_coeff_6_nxtber_more	:	bit_vector	:=	B"1111";
		gen3_coeff_6_preset_hint	:	bit_vector	:=	B"100";
		gen3_coeff_6_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_6_sel	:	string	:=	"preset_6";
		gen3_coeff_7	:	bit_vector	:=	B"000000000000000001";
		gen3_coeff_7_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_7_nxtber_less	:	bit_vector	:=	B"0001";
		gen3_coeff_7_nxtber_more	:	bit_vector	:=	B"0111";
		gen3_coeff_7_preset_hint	:	bit_vector	:=	B"010";
		gen3_coeff_7_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_7_sel	:	string	:=	"preset_7";
		gen3_coeff_8	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_8_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_8_nxtber_less	:	bit_vector	:=	B"0100";
		gen3_coeff_8_nxtber_more	:	bit_vector	:=	B"1000";
		gen3_coeff_8_preset_hint	:	bit_vector	:=	B"010";
		gen3_coeff_8_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_8_sel	:	string	:=	"preset_8";
		gen3_coeff_9	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_9_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_9_nxtber_less	:	bit_vector	:=	B"1011";
		gen3_coeff_9_nxtber_more	:	bit_vector	:=	B"1001";
		gen3_coeff_9_preset_hint	:	bit_vector	:=	B"011";
		gen3_coeff_9_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_9_sel	:	string	:=	"preset_9";
		gen3_coeff_delay_count	:	bit_vector	:=	B"1111101";
		gen3_coeff_errchk	:	string	:=	"enable";
		gen3_dcbal_en	:	string	:=	"true";
		gen3_diffclock_nfts_count	:	bit_vector	:=	B"10000000";
		gen3_force_local_coeff	:	string	:=	"false";
		gen3_full_swing	:	bit_vector	:=	B"111111";
		gen3_half_swing	:	string	:=	"false";
		gen3_low_freq	:	bit_vector	:=	B"000001";
		gen3_paritychk	:	string	:=	"enable";
		gen3_pl_framing_err_dis	:	string	:=	"enable";
		gen3_preset_coeff_1	:	bit_vector	:=	B"000000110101001010";
		gen3_preset_coeff_10	:	bit_vector	:=	B"001011110100000000";
		gen3_preset_coeff_11	:	bit_vector	:=	B"011110100001000000";
		gen3_preset_coeff_2	:	bit_vector	:=	B"000000110100001011";
		gen3_preset_coeff_3	:	bit_vector	:=	B"000000110010001101";
		gen3_preset_coeff_4	:	bit_vector	:=	B"000000110111001000";
		gen3_preset_coeff_5	:	bit_vector	:=	B"000000111111000000";
		gen3_preset_coeff_6	:	bit_vector	:=	B"000110111001000000";
		gen3_preset_coeff_7	:	bit_vector	:=	B"001000110111000000";
		gen3_preset_coeff_8	:	bit_vector	:=	B"000110101100001101";
		gen3_preset_coeff_9	:	bit_vector	:=	B"001000101111001000";
		gen3_reset_eieos_cnt_bit	:	string	:=	"false";
		gen3_rxfreqlock_counter	:	bit_vector	:=	B"00000000000000000000";
		gen3_sameclock_nfts_count	:	bit_vector	:=	B"10000000";
		gen3_scrdscr_bypass	:	string	:=	"false";
		gen3_skip_ph2_ph3	:	string	:=	"false";
		hard_reset_bypass	:	string	:=	"false";
		hard_rst_sig_chnl_en	:	string	:=	"disable_hrc_sig";
		hard_rst_tx_pll_rst_chnl_en	:	string	:=	"disable_hrc_txpll_rst";
		hip_ac_pwr_clk_freq_in_hz	:	bit_vector	:=	B"000000000000000000000000000000";
		hip_ac_pwr_uw_per_mhz	:	bit_vector	:=	B"000000000000000000000000000000";
		hip_base_address	:	bit_vector	:=	B"0000000000";
		hip_clock_dis	:	string	:=	"enable_hip_clk";
		hip_hard_reset	:	string	:=	"enable";
		hip_pcs_sig_chnl_en	:	string	:=	"disable_hip_pcs_sig";
		hot_plug_support	:	bit_vector	:=	B"0000000";
		hrc_chnl_txpll_master_cgb_rst_select	:	string	:=	"disable_master_cgb_sel";
		hrdrstctrl_en	:	string	:=	"hrdrstctrl_dis";
		iei_enable_settings	:	string	:=	"gen3gen2_infei_infsd_gen1_infei_sd";
		indicator	:	bit_vector	:=	B"111";
		intel_id_access	:	string	:=	"false";
		interrupt_pin	:	string	:=	"inta";
		io_window_addr_width	:	string	:=	"window_32_bit";
		jtag_id	:	string	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		ko_compl_data	:	bit_vector	:=	B"000000000000";
		ko_compl_header	:	bit_vector	:=	B"000000000000";
		l01_entry_latency	:	bit_vector	:=	B"11111";
		l0_exit_latency_diffclock	:	bit_vector	:=	B"110";
		l0_exit_latency_sameclock	:	bit_vector	:=	B"110";
		l0s_adj_rply_timer_dis	:	string	:=	"enable";
		l1_exit_latency_diffclock	:	bit_vector	:=	B"000";
		l1_exit_latency_sameclock	:	bit_vector	:=	B"000";
		l2_async_logic	:	string	:=	"enable";
		lane_mask	:	string	:=	"ln_mask_x4";
		lane_rate	:	string	:=	"gen1";
		link_width	:	string	:=	"x1";
		lmi_hold_off_cfg_timer_en	:	string	:=	"disable";
		low_priority_vc	:	string	:=	"single_vc_low_pr";
		ltr_mechanism	:	string	:=	"false";
		ltssm_1ms_timeout	:	string	:=	"disable";
		ltssm_freqlocked_check	:	string	:=	"disable";
		malformed_tlp_truncate_en	:	string	:=	"disable";
		max_link_width	:	string	:=	"x4_link_width";
		max_payload_size	:	string	:=	"payload_512";
		maximum_current	:	bit_vector	:=	B"000";
		millisecond_cycle_count	:	bit_vector	:=	B"00000000000000000000";
		msi_64bit_addressing_capable	:	string	:=	"true";
		msi_masking_capable	:	string	:=	"false";
		msi_multi_message_capable	:	string	:=	"count_4";
		msi_support	:	string	:=	"true";
		msix_pba_bir	:	bit_vector	:=	B"000";
		msix_pba_offset	:	bit_vector	:=	B"00000000000000000000000000000";
		msix_table_bir	:	bit_vector	:=	B"000";
		msix_table_offset	:	bit_vector	:=	B"00000000000000000000000000000";
		msix_table_size	:	bit_vector	:=	B"00000000000";
		national_inst_thru_enhance	:	string	:=	"true";
		no_command_completed	:	string	:=	"true";
		no_soft_reset	:	string	:=	"false";
		not_use_k_gbl_bits	:	string	:=	"not_used_k_gbl";
		operating_voltage	:	string	:=	"standard";
		pcie_base_spec	:	string	:=	"pcie_2p1";
		pcie_mode	:	string	:=	"shared_mode";
		pcie_spec_1p0_compliance	:	string	:=	"spec_1p1";
		pcie_spec_version	:	string	:=	"v2";
		pclk_out_sel	:	string	:=	"pclk";
		pld_in_use_reg	:	string	:=	"false";
		pm_latency_patch_dis	:	string	:=	"enable";
		pm_txdl_patch_dis	:	string	:=	"enable";
		pme_clock	:	string	:=	"false";
		port_link_number	:	bit_vector	:=	B"00000001";
		port_type	:	string	:=	"native_ep";
		powerdown_mode	:	string	:=	"powerup";
		prefetchable_mem_window_addr_width	:	string	:=	"prefetch_32";
		r2c_mask_easy	:	string	:=	"false";
		r2c_mask_enable	:	string	:=	"false";
		rec_frqlk_mon_en	:	string	:=	"disable";
		register_pipe_signals	:	string	:=	"true";
		retry_buffer_last_active_address	:	bit_vector	:=	B"1111111111";
		retry_buffer_memory_settings	:	string	:=	"000000000000000000000000000000000000";
		retry_ecc_corr_mask_dis	:	string	:=	"enable";
		revision_id	:	bit_vector	:=	B"00000001";
		role_based_error_reporting	:	string	:=	"false";
		rp_bug_fix_pri_sec_stat_reg	:	bit_vector	:=	B"1111111";
		rpltim_base	:	bit_vector	:=	B"00000000000000";
		rpltim_set	:	string	:=	"false";
		rstctl_ltssm_dis	:	string	:=	"false";
		rstctrl_1ms_count_fref_clk	:	bit_vector	:=	B"00001111010000100100";
		rstctrl_1us_count_fref_clk	:	bit_vector	:=	B"00000000000000111111";
		rstctrl_altpe3_crst_n_inv	:	string	:=	"false";
		rstctrl_altpe3_rst_n_inv	:	string	:=	"false";
		rstctrl_altpe3_srst_n_inv	:	string	:=	"false";
		rstctrl_chnl_cal_done_select	:	string	:=	"not_active_chnl_cal_done";
		rstctrl_debug_en	:	string	:=	"false";
		rstctrl_force_inactive_rst	:	string	:=	"false";
		rstctrl_fref_clk_select	:	string	:=	"ch0_sel";
		rstctrl_hard_block_enable	:	string	:=	"hard_rst_ctl";
		rstctrl_hip_ep	:	string	:=	"hip_ep";
		rstctrl_mask_tx_pll_lock_select	:	string	:=	"not_active_mask_tx_pll_lock";
		rstctrl_perst_enable	:	string	:=	"level";
		rstctrl_perstn_select	:	string	:=	"perstn_pin";
		rstctrl_pld_clr	:	string	:=	"false";
		rstctrl_pll_cal_done_select	:	string	:=	"not_active_pll_cal_done";
		rstctrl_rx_pcs_rst_n_inv	:	string	:=	"false";
		rstctrl_rx_pcs_rst_n_select	:	string	:=	"not_active_rx_pcs_rst";
		rstctrl_rx_pll_freq_lock_select	:	string	:=	"not_active_rx_pll_f_lock";
		rstctrl_rx_pll_lock_select	:	string	:=	"not_active_rx_pll_lock";
		rstctrl_rx_pma_rstb_inv	:	string	:=	"false";
		rstctrl_rx_pma_rstb_select	:	string	:=	"not_active_rx_pma_rstb";
		rstctrl_timer_a	:	bit_vector	:=	B"00001010";
		rstctrl_timer_a_type	:	string	:=	"a_timer_milli_secs";
		rstctrl_timer_b	:	bit_vector	:=	B"00001010";
		rstctrl_timer_b_type	:	string	:=	"b_timer_milli_secs";
		rstctrl_timer_c	:	bit_vector	:=	B"00001010";
		rstctrl_timer_c_type	:	string	:=	"c_timer_milli_secs";
		rstctrl_timer_d	:	bit_vector	:=	B"00010100";
		rstctrl_timer_d_type	:	string	:=	"d_timer_milli_secs";
		rstctrl_timer_e	:	bit_vector	:=	B"00000001";
		rstctrl_timer_e_type	:	string	:=	"e_timer_milli_secs";
		rstctrl_timer_f	:	bit_vector	:=	B"00001010";
		rstctrl_timer_f_type	:	string	:=	"f_timer_milli_secs";
		rstctrl_timer_g	:	bit_vector	:=	B"00001010";
		rstctrl_timer_g_type	:	string	:=	"g_timer_milli_secs";
		rstctrl_timer_h	:	bit_vector	:=	B"00000100";
		rstctrl_timer_h_type	:	string	:=	"h_timer_milli_secs";
		rstctrl_timer_i	:	bit_vector	:=	B"00010100";
		rstctrl_timer_i_type	:	string	:=	"i_timer_milli_secs";
		rstctrl_timer_j	:	bit_vector	:=	B"00010100";
		rstctrl_timer_j_type	:	string	:=	"j_timer_milli_secs";
		rstctrl_tx_lcff_pll_lock_select	:	string	:=	"not_active_lcff_pll_lock";
		rstctrl_tx_lcff_pll_rstb_select	:	string	:=	"not_active_lcff_pll_rstb";
		rstctrl_tx_pcs_rst_n_inv	:	string	:=	"false";
		rstctrl_tx_pcs_rst_n_select	:	string	:=	"not_active_tx_pcs_rst";
		rstctrl_tx_pma_rstb_inv	:	string	:=	"false";
		rstctrl_tx_pma_syncp_inv	:	string	:=	"false";
		rstctrl_tx_pma_syncp_select	:	string	:=	"not_active_tx_pma_syncp";
		rx_ast_parity	:	string	:=	"disable";
		rx_buffer_credit_alloc	:	string	:=	"balance";
		rx_buffer_fc_protect	:	bit_vector	:=	B"00000000000001000100";
		rx_buffer_protect	:	bit_vector	:=	B"00001000100";
		rx_cdc_almost_empty	:	bit_vector	:=	B"0011";
		rx_cdc_almost_full	:	bit_vector	:=	B"1100";
		rx_cred_ctl_param	:	string	:=	"disable";
		rx_ei_l0s	:	string	:=	"disable";
		rx_l0s_count_idl	:	bit_vector	:=	B"00000000";
		rx_ptr0_nonposted_dpram_max	:	bit_vector	:=	B"00000000000";
		rx_ptr0_nonposted_dpram_min	:	bit_vector	:=	B"00000000000";
		rx_ptr0_posted_dpram_max	:	bit_vector	:=	B"00000000000";
		rx_ptr0_posted_dpram_min	:	bit_vector	:=	B"00000000000";
		rx_runt_patch_dis	:	string	:=	"enable";
		rx_sop_ctrl	:	string	:=	"rx_sop_boundary_64";
		rx_trunc_patch_dis	:	string	:=	"enable";
		rx_use_prst	:	string	:=	"false";
		rx_use_prst_ep	:	string	:=	"true";
		rxbuf_ecc_corr_mask_dis	:	string	:=	"enable";
		rxdl_bad_sop_eop_filter_dis	:	string	:=	"rxdlbug1_enable_both";
		rxdl_bad_tlp_patch_dis	:	string	:=	"rxdlbug2_enable_both";
		rxdl_lcrc_patch_dis	:	string	:=	"rxdlbug3_enable_both";
		sameclock_nfts_count	:	bit_vector	:=	B"00000000";
		sel_enable_pcs_rx_fifo_err	:	string	:=	"disable_sel";
		silicon_rev	:	string	:=	"20nm5es";
		sim_mode	:	string	:=	"disable";
		simple_ro_fifo_control_en	:	string	:=	"disable";
		single_rx_detect	:	string	:=	"detect_all_lanes";
		skp_os_gen3_count	:	bit_vector	:=	B"00000000000";
		skp_os_schedule_count	:	bit_vector	:=	B"00000000000";
		slot_number	:	bit_vector	:=	B"0000000000000";
		slot_power_limit	:	bit_vector	:=	B"00000000";
		slot_power_scale	:	bit_vector	:=	B"00";
		slotclk_cfg	:	string	:=	"static_slotclkcfgon";
		ssid	:	bit_vector	:=	B"0000000000000000";
		ssvid	:	bit_vector	:=	B"0000000000000000";
		subsystem_device_id	:	bit_vector	:=	B"1110000000000001";
		subsystem_vendor_id	:	bit_vector	:=	B"0001000101110010";
		sup_mode	:	string	:=	"user_mode";
		surprise_down_error_support	:	string	:=	"false";
		tl_cfg_div	:	string	:=	"cfg_clk_div_7";
		tl_tx_check_parity_msg	:	string	:=	"disable";
		tph_completer	:	string	:=	"false";
		tx_ast_parity	:	string	:=	"disable";
		tx_cdc_almost_empty	:	bit_vector	:=	B"0101";
		tx_cdc_almost_full	:	bit_vector	:=	B"1100";
		tx_sop_ctrl	:	string	:=	"boundary_64";
		tx_swing	:	bit_vector	:=	B"00000000";
		txdl_fair_arbiter_counter	:	bit_vector	:=	B"0000";
		txdl_fair_arbiter_en	:	string	:=	"enable";
		txrate_adv	:	string	:=	"capability";
		uc_calibration_en	:	string	:=	"uc_calibration_dis";
		use_aer	:	string	:=	"false";
		use_crc_forwarding	:	string	:=	"false";
		user_id	:	bit_vector	:=	B"0000000000000000";
		vc0_clk_enable	:	string	:=	"true";
		vc0_rx_buffer_memory_settings	:	string	:=	"000000000000000000000000000000000000";
		vc0_rx_flow_ctrl_compl_data	:	bit_vector	:=	B"000111000000";
		vc0_rx_flow_ctrl_compl_header	:	bit_vector	:=	B"01110000";
		vc0_rx_flow_ctrl_nonposted_data	:	bit_vector	:=	B"00000000";
		vc0_rx_flow_ctrl_nonposted_header	:	bit_vector	:=	B"00110110";
		vc0_rx_flow_ctrl_posted_data	:	bit_vector	:=	B"000101101000";
		vc0_rx_flow_ctrl_posted_header	:	bit_vector	:=	B"00110010";
		vc1_clk_enable	:	string	:=	"false";
		vc_arbitration	:	string	:=	"single_vc_arb";
		vc_enable	:	string	:=	"single_vc";
		vendor_id	:	bit_vector	:=	B"0001000101110010";
		vsec_cap	:	bit_vector	:=	B"0000";
		vsec_id	:	bit_vector	:=	B"0001000101110010";
		wrong_device_id	:	string	:=	"disable"
	);
	port (
		-- Architecture ports
		aer_msi_num	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		app_int_err	:	in	std_logic_vector(1 downto 0)	:=	"00";
		app_inta_sts	:	in	std_logic	:=	'0';
		app_msi_num	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		app_msi_req	:	in	std_logic	:=	'0';
		app_msi_tc	:	in	std_logic_vector(2 downto 0)	:=	"000";
		atpg_los_en_n	:	in	std_logic	:=	'0';
		avmm_address	:	in	std_logic_vector(9 downto 0)	:=	"0000000000";
		avmm_byte_en	:	in	std_logic_vector(1 downto 0)	:=	"00";
		avmm_clk	:	in	std_logic	:=	'0';
		avmm_read	:	in	std_logic	:=	'0';
		avmm_rst_n	:	in	std_logic	:=	'0';
		avmm_write	:	in	std_logic	:=	'0';
		avmm_writedata	:	in	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		bist_scanen	:	in	std_logic	:=	'0';
		bist_scanin	:	in	std_logic	:=	'0';
		bisten_rcv_n	:	in	std_logic	:=	'0';
		bisten_rpl_n	:	in	std_logic	:=	'0';
		bistmode_n	:	in	std_logic	:=	'0';
		cfg_link2csr_pld	:	in	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		cfg_prmbus_pld	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		chnl_cal_done0	:	in	std_logic	:=	'0';
		chnl_cal_done1	:	in	std_logic	:=	'0';
		chnl_cal_done2	:	in	std_logic	:=	'0';
		chnl_cal_done3	:	in	std_logic	:=	'0';
		chnl_cal_done4	:	in	std_logic	:=	'0';
		chnl_cal_done5	:	in	std_logic	:=	'0';
		chnl_cal_done6	:	in	std_logic	:=	'0';
		chnl_cal_done7	:	in	std_logic	:=	'0';
		core_clk_in	:	in	std_logic	:=	'0';
		core_crst	:	in	std_logic	:=	'0';
		core_por	:	in	std_logic	:=	'0';
		core_rst	:	in	std_logic	:=	'0';
		core_srst	:	in	std_logic	:=	'0';
		cpl_err	:	in	std_logic_vector(6 downto 0)	:=	"0000000";
		cpl_pending	:	in	std_logic	:=	'0';
		cseb_rddata	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		cseb_rddata_parity	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		cseb_rdresponse	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		cseb_waitrequest	:	in	std_logic	:=	'0';
		cseb_wrresp_valid	:	in	std_logic	:=	'0';
		cseb_wrresponse	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		csr_cbdin	:	in	std_logic	:=	'0';
		csr_clk	:	in	std_logic	:=	'0';
		csr_din	:	in	std_logic	:=	'0';
		csr_en	:	in	std_logic	:=	'0';
		csr_enscan	:	in	std_logic	:=	'0';
		csr_entest	:	in	std_logic	:=	'0';
		csr_in	:	in	std_logic	:=	'0';
		csr_load_csr	:	in	std_logic	:=	'0';
		csr_pipe_in	:	in	std_logic	:=	'0';
		csr_seg	:	in	std_logic	:=	'0';
		csr_tcsrin	:	in	std_logic	:=	'0';
		csr_tverify	:	in	std_logic	:=	'0';
		cvp_config_done	:	in	std_logic	:=	'0';
		cvp_config_error	:	in	std_logic	:=	'0';
		cvp_config_ready	:	in	std_logic	:=	'0';
		cvp_en	:	in	std_logic	:=	'0';
		egress_blk_err	:	in	std_logic	:=	'0';
		entest	:	in	std_logic	:=	'0';
		flr_reset	:	in	std_logic	:=	'0';
		force_tx_eidle	:	in	std_logic	:=	'0';
		fref_clk0	:	in	std_logic	:=	'0';
		fref_clk1	:	in	std_logic	:=	'0';
		fref_clk2	:	in	std_logic	:=	'0';
		fref_clk3	:	in	std_logic	:=	'0';
		fref_clk4	:	in	std_logic	:=	'0';
		fref_clk5	:	in	std_logic	:=	'0';
		fref_clk6	:	in	std_logic	:=	'0';
		fref_clk7	:	in	std_logic	:=	'0';
		frzlogic	:	in	std_logic	:=	'0';
		frzreg	:	in	std_logic	:=	'0';
		hold_ltssm_rec	:	in	std_logic	:=	'0';
		hpg_ctrler	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		iocsrrdy_dly	:	in	std_logic	:=	'0';
		lmi_addr	:	in	std_logic_vector(11 downto 0)	:=	"000000000000";
		lmi_din	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		lmi_rden	:	in	std_logic	:=	'0';
		lmi_wren	:	in	std_logic	:=	'0';
		m10k_select	:	in	std_logic_vector(2 downto 0)	:=	"000";
		mask_tx_pll_lock0	:	in	std_logic	:=	'0';
		mask_tx_pll_lock1	:	in	std_logic	:=	'0';
		mask_tx_pll_lock2	:	in	std_logic	:=	'0';
		mask_tx_pll_lock3	:	in	std_logic	:=	'0';
		mask_tx_pll_lock4	:	in	std_logic	:=	'0';
		mask_tx_pll_lock5	:	in	std_logic	:=	'0';
		mask_tx_pll_lock6	:	in	std_logic	:=	'0';
		mask_tx_pll_lock7	:	in	std_logic	:=	'0';
		mem_hip_test_enable	:	in	std_logic	:=	'0';
		mem_regscanen_n	:	in	std_logic	:=	'0';
		mem_rscin_rcv_bot	:	in	std_logic	:=	'0';
		mem_rscin_rcv_top	:	in	std_logic	:=	'0';
		mem_rscin_rtry	:	in	std_logic	:=	'0';
		nfrzdrv	:	in	std_logic	:=	'0';
		npor	:	in	std_logic	:=	'0';
		pclk_central	:	in	std_logic	:=	'0';
		pclk_ch0	:	in	std_logic	:=	'0';
		pclk_ch1	:	in	std_logic	:=	'0';
		pex_msi_num	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		phy_rst	:	in	std_logic	:=	'0';
		phy_srst	:	in	std_logic	:=	'0';
		phystatus0	:	in	std_logic	:=	'0';
		phystatus1	:	in	std_logic	:=	'0';
		phystatus2	:	in	std_logic	:=	'0';
		phystatus3	:	in	std_logic	:=	'0';
		phystatus4	:	in	std_logic	:=	'0';
		phystatus5	:	in	std_logic	:=	'0';
		phystatus6	:	in	std_logic	:=	'0';
		phystatus7	:	in	std_logic	:=	'0';
		pin_perst_n	:	in	std_logic	:=	'0';
		pld_clk	:	in	std_logic	:=	'0';
		pld_clrhip_n	:	in	std_logic	:=	'0';
		pld_clrpcship_n	:	in	std_logic	:=	'0';
		pld_clrpmapcship_n	:	in	std_logic	:=	'0';
		pld_core_ready	:	in	std_logic	:=	'0';
		pld_gp_status	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		pld_perst_n	:	in	std_logic	:=	'0';
		pll_cal_done0	:	in	std_logic	:=	'0';
		pll_cal_done1	:	in	std_logic	:=	'0';
		pll_cal_done2	:	in	std_logic	:=	'0';
		pll_cal_done3	:	in	std_logic	:=	'0';
		pll_cal_done4	:	in	std_logic	:=	'0';
		pll_cal_done5	:	in	std_logic	:=	'0';
		pll_cal_done6	:	in	std_logic	:=	'0';
		pll_cal_done7	:	in	std_logic	:=	'0';
		pll_fixed_clk_central	:	in	std_logic	:=	'0';
		pll_fixed_clk_ch0	:	in	std_logic	:=	'0';
		pll_fixed_clk_ch1	:	in	std_logic	:=	'0';
		plniotri	:	in	std_logic	:=	'0';
		pm_auxpwr	:	in	std_logic	:=	'0';
		pm_data	:	in	std_logic_vector(9 downto 0)	:=	"0000000000";
		pm_event	:	in	std_logic	:=	'0';
		pm_exit_d0_ack	:	in	std_logic	:=	'0';
		pme_to_cr	:	in	std_logic	:=	'0';
		reserved_clk_in	:	in	std_logic	:=	'0';
		reserved_in	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		rx_cred_ctl	:	in	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		rx_pll_freq_lock0	:	in	std_logic	:=	'0';
		rx_pll_freq_lock1	:	in	std_logic	:=	'0';
		rx_pll_freq_lock2	:	in	std_logic	:=	'0';
		rx_pll_freq_lock3	:	in	std_logic	:=	'0';
		rx_pll_freq_lock4	:	in	std_logic	:=	'0';
		rx_pll_freq_lock5	:	in	std_logic	:=	'0';
		rx_pll_freq_lock6	:	in	std_logic	:=	'0';
		rx_pll_freq_lock7	:	in	std_logic	:=	'0';
		rx_pll_phase_lock0	:	in	std_logic	:=	'0';
		rx_pll_phase_lock1	:	in	std_logic	:=	'0';
		rx_pll_phase_lock2	:	in	std_logic	:=	'0';
		rx_pll_phase_lock3	:	in	std_logic	:=	'0';
		rx_pll_phase_lock4	:	in	std_logic	:=	'0';
		rx_pll_phase_lock5	:	in	std_logic	:=	'0';
		rx_pll_phase_lock6	:	in	std_logic	:=	'0';
		rx_pll_phase_lock7	:	in	std_logic	:=	'0';
		rx_st_mask	:	in	std_logic	:=	'0';
		rx_st_ready	:	in	std_logic	:=	'0';
		rxblkst0	:	in	std_logic	:=	'0';
		rxblkst1	:	in	std_logic	:=	'0';
		rxblkst2	:	in	std_logic	:=	'0';
		rxblkst3	:	in	std_logic	:=	'0';
		rxblkst4	:	in	std_logic	:=	'0';
		rxblkst5	:	in	std_logic	:=	'0';
		rxblkst6	:	in	std_logic	:=	'0';
		rxblkst7	:	in	std_logic	:=	'0';
		rxdata0	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata1	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata2	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata3	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata4	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata5	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata6	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata7	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdatak0	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak1	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak2	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak3	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak4	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak5	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak6	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak7	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdataskip0	:	in	std_logic	:=	'0';
		rxdataskip1	:	in	std_logic	:=	'0';
		rxdataskip2	:	in	std_logic	:=	'0';
		rxdataskip3	:	in	std_logic	:=	'0';
		rxdataskip4	:	in	std_logic	:=	'0';
		rxdataskip5	:	in	std_logic	:=	'0';
		rxdataskip6	:	in	std_logic	:=	'0';
		rxdataskip7	:	in	std_logic	:=	'0';
		rxelecidle0	:	in	std_logic	:=	'0';
		rxelecidle1	:	in	std_logic	:=	'0';
		rxelecidle2	:	in	std_logic	:=	'0';
		rxelecidle3	:	in	std_logic	:=	'0';
		rxelecidle4	:	in	std_logic	:=	'0';
		rxelecidle5	:	in	std_logic	:=	'0';
		rxelecidle6	:	in	std_logic	:=	'0';
		rxelecidle7	:	in	std_logic	:=	'0';
		rxfreqlocked0	:	in	std_logic	:=	'0';
		rxfreqlocked1	:	in	std_logic	:=	'0';
		rxfreqlocked2	:	in	std_logic	:=	'0';
		rxfreqlocked3	:	in	std_logic	:=	'0';
		rxfreqlocked4	:	in	std_logic	:=	'0';
		rxfreqlocked5	:	in	std_logic	:=	'0';
		rxfreqlocked6	:	in	std_logic	:=	'0';
		rxfreqlocked7	:	in	std_logic	:=	'0';
		rxstatus0	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus1	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus2	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus3	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus4	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus5	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus6	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus7	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxsynchd0	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd1	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd2	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd3	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd4	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd5	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd6	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd7	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxvalid0	:	in	std_logic	:=	'0';
		rxvalid1	:	in	std_logic	:=	'0';
		rxvalid2	:	in	std_logic	:=	'0';
		rxvalid3	:	in	std_logic	:=	'0';
		rxvalid4	:	in	std_logic	:=	'0';
		rxvalid5	:	in	std_logic	:=	'0';
		rxvalid6	:	in	std_logic	:=	'0';
		rxvalid7	:	in	std_logic	:=	'0';
		scan_mode_n	:	in	std_logic	:=	'0';
		scan_shift_n	:	in	std_logic	:=	'0';
		sw_ctmod	:	in	std_logic_vector(1 downto 0)	:=	"00";
		swdn_in	:	in	std_logic_vector(2 downto 0)	:=	"000";
		swup_in	:	in	std_logic_vector(6 downto 0)	:=	"0000000";
		test_in_1_hip	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		test_in_hip	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		test_pl_dbg_eqin	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		tx_cred_cons_select	:	in	std_logic	:=	'0';
		tx_cred_fc_sel	:	in	std_logic_vector(1 downto 0)	:=	"00";
		tx_lcff_pll_lock0	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock1	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock2	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock3	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock4	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock5	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock6	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock7	:	in	std_logic	:=	'0';
		tx_st_data	:	in	std_logic_vector(255 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		tx_st_empty	:	in	std_logic_vector(1 downto 0)	:=	"00";
		tx_st_eop	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		tx_st_err	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		tx_st_parity	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		tx_st_sop	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		tx_st_valid	:	in	std_logic	:=	'0';
		user_mode	:	in	std_logic	:=	'0';
		sta_hd_altpe3_hip_core_top_hd_altpe3_hip_core_u_clkmux_core_clk_cnt_reg_0_0_Q	:	out	std_logic	:=	'0';
		sta_hd_altpe3_hip_core_top_hd_altpe3_hip_core_u_clkmux_core_clk_cnt_reg_1_0_Q	:	out	std_logic	:=	'0';
		sta_hd_altpe3_hip_core_top_hd_altpe3_hip_core_u_clkmux_core_clk_cnt_reg_2_0_Q	:	out	std_logic	:=	'0';
		app_inta_ack	:	out	std_logic	:=	'0';
		app_msi_ack	:	out	std_logic	:=	'0';
		avmm_readdata	:	out	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		cfg_par_err	:	out	std_logic	:=	'0';
		core_clk_out	:	out	std_logic	:=	'0';
		cseb_addr	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		cseb_addr_parity	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		cseb_be	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		cseb_is_shadow	:	out	std_logic	:=	'0';
		cseb_rden	:	out	std_logic	:=	'0';
		cseb_wrdata	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		cseb_wrdata_parity	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		cseb_wren	:	out	std_logic	:=	'0';
		cseb_wrresp_req	:	out	std_logic	:=	'0';
		csr_dout	:	out	std_logic	:=	'0';
		csr_out	:	out	std_logic	:=	'0';
		csr_pipe_out	:	out	std_logic	:=	'0';
		current_coeff0	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff1	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff2	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff3	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff4	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff5	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff6	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff7	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_rxpreset0	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset1	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset2	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset3	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset4	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset5	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset6	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset7	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_speed	:	out	std_logic_vector(1 downto 0)	:=	"00";
		cvp_clk	:	out	std_logic	:=	'0';
		cvp_config	:	out	std_logic	:=	'0';
		cvp_data	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		cvp_full_config	:	out	std_logic	:=	'0';
		cvp_start_xfer	:	out	std_logic	:=	'0';
		dl_up	:	out	std_logic	:=	'0';
		dlup_exit	:	out	std_logic	:=	'0';
		eidle_infer_sel0	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel1	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel2	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel3	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel4	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel5	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel6	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel7	:	out	std_logic_vector(2 downto 0)	:=	"000";
		ev_128ns	:	out	std_logic	:=	'0';
		ev_1us	:	out	std_logic	:=	'0';
		flr_sts	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n0	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n1	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n2	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n3	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n4	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n5	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n6	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n7	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n0	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n1	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n2	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n3	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n4	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n5	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n6	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n7	:	out	std_logic	:=	'0';
		hotrst_exit	:	out	std_logic	:=	'0';
		int_status	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		k_hip_pcs_chnl_en	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		k_hrc_chnl_en	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		k_hrc_chnl_txpll_master_cgb_rst_en	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		k_hrc_chnl_txpll_rst_en	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		l2_exit	:	out	std_logic	:=	'0';
		lane_act	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		lmi_ack	:	out	std_logic	:=	'0';
		lmi_dout	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		ltssm_state	:	out	std_logic_vector(4 downto 0)	:=	"00000";
		mem_rscout_rcv_bot	:	out	std_logic	:=	'0';
		mem_rscout_rcv_top	:	out	std_logic	:=	'0';
		mem_rscout_rtry	:	out	std_logic	:=	'0';
		pld_clk_in_use	:	out	std_logic	:=	'0';
		pld_gp_ctrl	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		pm_exit_d0_req	:	out	std_logic	:=	'0';
		pme_to_sr	:	out	std_logic	:=	'0';
		powerdown0	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown1	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown2	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown3	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown4	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown5	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown6	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown7	:	out	std_logic_vector(1 downto 0)	:=	"00";
		r2c_unc_ecc	:	out	std_logic	:=	'0';
		rate0	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate1	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate2	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate3	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate4	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate5	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate6	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate7	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate_ctrl	:	out	std_logic_vector(1 downto 0)	:=	"00";
		reserved_clk_out	:	out	std_logic	:=	'0';
		reserved_out	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		reset_status	:	out	std_logic	:=	'0';
		retry_corr_ecc	:	out	std_logic	:=	'0';
		retry_unc_ecc	:	out	std_logic	:=	'0';
		rx_corr_ecc	:	out	std_logic	:=	'0';
		rx_cred_status	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		rx_par_err	:	out	std_logic	:=	'0';
		rx_pcs_rst_n0	:	out	std_logic	:=	'0';
		rx_pcs_rst_n1	:	out	std_logic	:=	'0';
		rx_pcs_rst_n2	:	out	std_logic	:=	'0';
		rx_pcs_rst_n3	:	out	std_logic	:=	'0';
		rx_pcs_rst_n4	:	out	std_logic	:=	'0';
		rx_pcs_rst_n5	:	out	std_logic	:=	'0';
		rx_pcs_rst_n6	:	out	std_logic	:=	'0';
		rx_pcs_rst_n7	:	out	std_logic	:=	'0';
		rx_pma_rstb0	:	out	std_logic	:=	'0';
		rx_pma_rstb1	:	out	std_logic	:=	'0';
		rx_pma_rstb2	:	out	std_logic	:=	'0';
		rx_pma_rstb3	:	out	std_logic	:=	'0';
		rx_pma_rstb4	:	out	std_logic	:=	'0';
		rx_pma_rstb5	:	out	std_logic	:=	'0';
		rx_pma_rstb6	:	out	std_logic	:=	'0';
		rx_pma_rstb7	:	out	std_logic	:=	'0';
		rx_st_bardec1	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		rx_st_bardec2	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		rx_st_be	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rx_st_data	:	out	std_logic_vector(255 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		rx_st_empty	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rx_st_eop	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		rx_st_err	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		rx_st_parity	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rx_st_sop	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		rx_st_valid	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		rxfc_cplbuf_ovf	:	out	std_logic	:=	'0';
		rxfc_cplovf_tag	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		rxpolarity0	:	out	std_logic	:=	'0';
		rxpolarity1	:	out	std_logic	:=	'0';
		rxpolarity2	:	out	std_logic	:=	'0';
		rxpolarity3	:	out	std_logic	:=	'0';
		rxpolarity4	:	out	std_logic	:=	'0';
		rxpolarity5	:	out	std_logic	:=	'0';
		rxpolarity6	:	out	std_logic	:=	'0';
		rxpolarity7	:	out	std_logic	:=	'0';
		serr_out	:	out	std_logic	:=	'0';
		swdn_out	:	out	std_logic_vector(6 downto 0)	:=	"0000000";
		swup_out	:	out	std_logic_vector(2 downto 0)	:=	"000";
		test_fref_clk	:	out	std_logic	:=	'0';
		test_out_1_hip	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		test_out_hip	:	out	std_logic_vector(255 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		tl_cfg_add	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		tl_cfg_ctl	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		tl_cfg_sts	:	out	std_logic_vector(52 downto 0)	:=	"00000000000000000000000000000000000000000000000000000";
		tl_cfg_sts_wr	:	out	std_logic	:=	'0';
		tx_cred_data_fc	:	out	std_logic_vector(11 downto 0)	:=	"000000000000";
		tx_cred_fc_hip_cons	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		tx_cred_fc_infinite	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		tx_cred_hdr_fc	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		tx_deemph0	:	out	std_logic	:=	'0';
		tx_deemph1	:	out	std_logic	:=	'0';
		tx_deemph2	:	out	std_logic	:=	'0';
		tx_deemph3	:	out	std_logic	:=	'0';
		tx_deemph4	:	out	std_logic	:=	'0';
		tx_deemph5	:	out	std_logic	:=	'0';
		tx_deemph6	:	out	std_logic	:=	'0';
		tx_deemph7	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb0	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb1	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb2	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb3	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb4	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb5	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb6	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb7	:	out	std_logic	:=	'0';
		tx_margin0	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin1	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin2	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin3	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin4	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin5	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin6	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin7	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_par_err	:	out	std_logic_vector(1 downto 0)	:=	"00";
		tx_pcs_rst_n0	:	out	std_logic	:=	'0';
		tx_pcs_rst_n1	:	out	std_logic	:=	'0';
		tx_pcs_rst_n2	:	out	std_logic	:=	'0';
		tx_pcs_rst_n3	:	out	std_logic	:=	'0';
		tx_pcs_rst_n4	:	out	std_logic	:=	'0';
		tx_pcs_rst_n5	:	out	std_logic	:=	'0';
		tx_pcs_rst_n6	:	out	std_logic	:=	'0';
		tx_pcs_rst_n7	:	out	std_logic	:=	'0';
		tx_pma_syncp0	:	out	std_logic	:=	'0';
		tx_pma_syncp1	:	out	std_logic	:=	'0';
		tx_pma_syncp2	:	out	std_logic	:=	'0';
		tx_pma_syncp3	:	out	std_logic	:=	'0';
		tx_pma_syncp4	:	out	std_logic	:=	'0';
		tx_pma_syncp5	:	out	std_logic	:=	'0';
		tx_pma_syncp6	:	out	std_logic	:=	'0';
		tx_pma_syncp7	:	out	std_logic	:=	'0';
		tx_st_ready	:	out	std_logic	:=	'0';
		txblkst0	:	out	std_logic	:=	'0';
		txblkst1	:	out	std_logic	:=	'0';
		txblkst2	:	out	std_logic	:=	'0';
		txblkst3	:	out	std_logic	:=	'0';
		txblkst4	:	out	std_logic	:=	'0';
		txblkst5	:	out	std_logic	:=	'0';
		txblkst6	:	out	std_logic	:=	'0';
		txblkst7	:	out	std_logic	:=	'0';
		txcompl0	:	out	std_logic	:=	'0';
		txcompl1	:	out	std_logic	:=	'0';
		txcompl2	:	out	std_logic	:=	'0';
		txcompl3	:	out	std_logic	:=	'0';
		txcompl4	:	out	std_logic	:=	'0';
		txcompl5	:	out	std_logic	:=	'0';
		txcompl6	:	out	std_logic	:=	'0';
		txcompl7	:	out	std_logic	:=	'0';
		txdata0	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata1	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata2	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata3	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata4	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata5	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata6	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata7	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdatak0	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak1	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak2	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak3	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak4	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak5	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak6	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak7	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdataskip0	:	out	std_logic	:=	'0';
		txdataskip1	:	out	std_logic	:=	'0';
		txdataskip2	:	out	std_logic	:=	'0';
		txdataskip3	:	out	std_logic	:=	'0';
		txdataskip4	:	out	std_logic	:=	'0';
		txdataskip5	:	out	std_logic	:=	'0';
		txdataskip6	:	out	std_logic	:=	'0';
		txdataskip7	:	out	std_logic	:=	'0';
		txdetectrx0	:	out	std_logic	:=	'0';
		txdetectrx1	:	out	std_logic	:=	'0';
		txdetectrx2	:	out	std_logic	:=	'0';
		txdetectrx3	:	out	std_logic	:=	'0';
		txdetectrx4	:	out	std_logic	:=	'0';
		txdetectrx5	:	out	std_logic	:=	'0';
		txdetectrx6	:	out	std_logic	:=	'0';
		txdetectrx7	:	out	std_logic	:=	'0';
		txelecidle0	:	out	std_logic	:=	'0';
		txelecidle1	:	out	std_logic	:=	'0';
		txelecidle2	:	out	std_logic	:=	'0';
		txelecidle3	:	out	std_logic	:=	'0';
		txelecidle4	:	out	std_logic	:=	'0';
		txelecidle5	:	out	std_logic	:=	'0';
		txelecidle6	:	out	std_logic	:=	'0';
		txelecidle7	:	out	std_logic	:=	'0';
		txst_prot_err	:	out	std_logic	:=	'0';
		txswing0	:	out	std_logic	:=	'0';
		txswing1	:	out	std_logic	:=	'0';
		txswing2	:	out	std_logic	:=	'0';
		txswing3	:	out	std_logic	:=	'0';
		txswing4	:	out	std_logic	:=	'0';
		txswing5	:	out	std_logic	:=	'0';
		txswing6	:	out	std_logic	:=	'0';
		txswing7	:	out	std_logic	:=	'0';
		txsynchd0	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd1	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd2	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd3	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd4	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd5	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd6	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd7	:	out	std_logic_vector(1 downto 0)	:=	"00";
		wake_oen	:	out	std_logic	:=	'0'
	);
end component;

end twentynm_hip_components;

package body TWENTYNM_HIP_COMPONENTS is

function bin2int (s : std_logic_vector) return integer is

      constant temp      : std_logic_vector(s'high-s'low DOWNTO 0) := s;      
      variable result      : integer := 0;
   begin
      for i in temp'range loop
         if (temp(i) = '1') then
            result := result + (2**i);
         end if;
      end loop;
      return(result);
   end bin2int;

function bin2int (s : bit_vector) return integer is

      constant temp      : bit_vector(s'high-s'low DOWNTO 0) := s;      
      variable result      : integer := 0;
   begin
      for i in temp'range loop
         if (temp(i) = '1') then
            result := result + (2**i);
         end if;
      end loop;
      return(result);
   end bin2int;
                  
function bin2int (s : std_logic) return integer is
      constant temp      : std_logic := s;      
      variable result      : integer := 0;
   begin
         if (temp = '1') then
            result := 1;
         else
         	result := 0;
     	 end if;
      return(result);
	end bin2int;
                  
function bin2int (s : bit) return integer is
      constant temp      : bit := s;      
      variable result      : integer := 0;
   begin
         if (temp = '1') then
            result := 1;
         else
         	result := 0;
     	 end if;
      return(result);
	end bin2int;
	
function str2bin (s : string) return std_logic_vector is
variable len : integer := s'length;
variable result : std_logic_vector(39 DOWNTO 0) := (OTHERS => '0');
variable i : integer;
begin
    for i in 1 to len loop
        case s(i) is
            when '0' => result(len - i) := '0';
            when '1' => result(len - i) := '1';
            when others =>
                ASSERT FALSE
                REPORT "Illegal Character "&  s(i) & "in string parameter! "
                SEVERITY ERROR;
        end case;
    end loop;
    return result;
end;

function str2int (s : string) return integer is
variable len : integer := s'length;
variable newdigit : integer := 0;
variable sign : integer := 1;
variable digit : integer := 0;
begin
    for i in 1 to len loop
        case s(i) is
            when '-' =>
                if i = 1 then
                    sign := -1;
                else
                    ASSERT FALSE
                    REPORT "Illegal Character "&  s(i) & "i n string parameter! " SEVERITY ERROR;
                end if;
            when '0' =>
                digit := 0;
            when '1' =>
                digit := 1;
            when '2' =>
                digit := 2;
            when '3' =>
                digit := 3;
            when '4' =>
                digit := 4;
            when '5' =>
                digit := 5;
            when '6' =>
                digit := 6;
            when '7' =>
                digit := 7;
            when '8' =>
                digit := 8;
            when '9' =>
                digit := 9;
            when others =>
                ASSERT FALSE
                REPORT "Illegal Character "&  s(i) & "in string parameter! "
                SEVERITY ERROR;
        end case;
        newdigit := newdigit * 10 + digit;
    end loop;

    return (sign*newdigit);
end;

function int2bin (arg : integer; size : integer) return std_logic_vector is
    variable int_val : integer := arg;
    variable result : std_logic_vector(size-1 downto 0);
    begin
        for i in 0 to result'left loop
            if ((int_val mod 2) = 0) then
                result(i) := '0';
            else
                result(i) := '1';
            end if;
            int_val := int_val/2;
        end loop;
        return result;
    end int2bin;
    
function int2bin (arg : boolean; size : integer) return std_logic_vector is
    variable result : std_logic_vector(size-1 downto 0);
    begin
		if(arg)then
			result := (OTHERS => '1');
		else
			result := (OTHERS => '0');
		end if;
        return result;
    end int2bin;

function int2bit (arg : integer) return std_logic is
    variable int_val : integer := arg;
    variable result : std_logic;
    begin
        
            if (int_val  = 0) then
                result := '0';
            else
                result := '1';
            end if;
            
        return result;
end int2bit;

function int2bit (arg : boolean) return std_logic is
    variable int_val : boolean := arg;
    variable result : std_logic;
    begin
        
            if (int_val ) then
                result := '1';
            else
                result := '0';
            end if;
            
        return result;
end int2bit;

end TWENTYNM_HIP_COMPONENTS;
