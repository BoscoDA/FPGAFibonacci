// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std.1
// ALTERA_TIMESTAMP:Thu Jun  8 04:05:47 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Nm5N+8CcHma9koQ7HsVsY0x/aeZShHwpcUc+AyRqajwfdyh67jp10IQIq+1YShid
JAOAf8Lcem3kOcyb/3oCGGrA4tiAFgQtZwoPJgCkRQ2EOerFxXPf2NhF/bLonMyO
3ulKw5n4vCHiHmIRQJlPOYII18Hm8W73C0fU7CybChc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1429888)
wHv1UhRqJv30JkoTirx17s8zOXywNayp8PcsWKbQeOqXAB9uEls/cY2isRwkcbh4
nv1wlSc6D1LAGRkR8Z3cHjwN95+QsFLxKlSnbmFolY2QIoHXxfRkxXULH/fcHmhD
B4b22+6ztMHkAtH0Hr65U2lKzfHIpU2UGAadSineKFwr67o2aHZobnphnZEFiVTC
y+vvr/JmvMN9qi2ZqTSkNs42PouCs5sXaFbXYN20NX9CBqtH60V7HmbHcUoG2qxx
tvVcL+4bFB3QRiA/hdRfrElDSREyNGqDbDR+UiLotrXlQE37CQT7DMYQXT2dy/iX
Z46pIWNQhZTsu348/ABo9bJA0ikkPnegIFAfLtqV+C4yc457N2+y/qCpjWpHGGib
tZHZl8RbrQWbyYfk6+oTO2vFpQayD82dkYk2usXFpHXGBfusHd3qwnH/8BSya4qM
Qz2jmd5mF9fJXf93/TuizjdRUaGcFqFLJ5obdnejZ96hWPZAqvj8fReOR64L8N/d
cJUbSPq1PooDeUg6+7DOHPLCfBxoDZLHsfM1lh4YXDSaB/XgM59v0hFqoCD0iiNu
JRbL1kEJtnZFeqfskU69xA8oLzf8+QqppBZ2zU5Ot8I19vD4V37yyvZN4TkF+uit
nhd9Cd9fuxux9IwTPMA+A+oSy3VdF+gQMZcA66xbNgL+WcV/F7aP8oA7bJknGrWB
yYqPeV7uyTAqfmm29cqjCyUbjAUlQ9oAG2ad9rzVmBP7iSAVDSdgCi3bCcq2BSL6
MhokoS9gWrhRgIci4qeG/KtlhL2uXajy+FGtA00c0uvU3y7Z5Fd6b3pFQjYoPjX2
nJpobzMExoBvx8mrCKhaz8Sef9HNZH7Zuz2sn6WEJvi8EGqr+0q8HFH4x6n4To56
xeyMvxLzcjnEpu7x9BU8Q2M+MFaVtrMQDYMTf6yc0bCkNAB15hgSSRpDfAp6St2e
XaxrHAm5aIuOUPZdkfSWHBHmCYBEG3N8ci+grNax5ETQ3srQAA94ZyMPtFRWcK3M
bYXtlRg9kIPx+wBRSCPN8r9HfRbAeKFnK6qz6byxPzvMLfTbIkN1Wc0ihrqKBV+G
tZ9NEHLMg6PVwtkTyQPyGgRJaePpi8zYD2jCdoJIqoOwVvrDySPszDVGFTAJ+qTO
JZbLRcGX4cliW9gcvSskX45F/P48Dz0nd3LadR/NwNI97hBtVvxabrLvdq+uB9jq
eq9xn5cdaT+yGgKtjjvcm9ykrs6ZYfCyo0PpXkGzn8VGBs9GAyvzw0PdCEA81y5V
k+mNXAkIqVKxEEStv+pkRD7Ci9JPpI6VGnoDx4PeuPQqDQMAIVvzwclGt9oXYiWL
4RJ9DSr1sEbhC7EFnFM4PfZ9g059M7rj1VXs+jpf8XGa11FlX+nAWxrgDPo2nwyO
mNNF1PVBBKUN+9ycnJHhLUhshqINX+RsRHoyl3ZKd/71lhMNEJJ9+a4Wkeh26R9U
+hmNZhWx04O+D5cgmY9hTIDJn/wsCkRcTOid3aN3sHCYQkv8hznYFhGx8tJJ+fAx
vdBf3xynZYCaSOdvo2GlcpL+pnHeDsQX8lcwZNWJNcP199uCvRc3oG7VY4uBGQsg
DC3u1erLxGaDbltyci6phqqlxQA/WYsL3XVQMvIXvKcOQ8Jsd/LzKbIytev5zcLk
7BCiNqS3QGoTYcuXwRCkTSW1WYjVauYRc3vm4i4rfiKjCNKroVnKQz5x0zmv9sEN
yVwhIOekLWfAUCrcSfcL/mrKcKIoXG7B3Yk+FXla9bEBVfyYdou6yqyQ2i34xksL
aMteb2jg4xxrB7uXVWMmoTzWFlJN/ClxYERAbQCabG69PAlV1mbToX/6w4ZJuD+h
gmdt5kOBSILuaYRY2SzVjfzalW+ugPkxNwINd+7+Xsdt+QM/eg7W9lrT/gDHhMtX
Ww6vdom/u0hfJyxHR2ukWlmZXk2ofU4p3noJImEu3tCHZwyWxS+IgP1x1x0h/9GP
YLLlT9NaELnI2nfjYleHA36CuMv2ATMmKYKsK0y9xSGVxdaKoXDUuSQFURX7C5jo
4r+C6WD52Eds8YLs/n3sYIYm5CuKNxryDHWPvwKzzDUq50DqRsvlpMtoWezIxIMR
MWU6wovk1sgSedWoO9nW0CJ4z4mPW9lZw48p3Fcg9Io/aI2ehAPSHKzcdtzlL4W9
WbPAhuyofz2TKskWs/7uhEqMWETqLDgDxqXCNLSKIR6FsQGTIboehxnxh7puKre5
olibpabYUDc7jveIfAc/6UzTZEx1mYMZkKddLmqhB1/fLhRhbEhmyL1ziVZZHqkN
BfvveE6Uk4pHeghdsOGYpAD6qeHJlLUmPkpT2rBunSrjLJO4TKbhSYQoHoj9FYuu
SQHjTrk4DlfojuLgf0er7tGSh9BzE9JXysiQ98/k46//FFsSGQGGI6Os8y1H9v5v
kNWv6dEHreNWSRdF8UsUwisWHzeU/qGfGfErjrASCb1ySohCfCN5oaYaNXMFvCUD
3yeT6Sy9Hmab4QgWJM8FgSnt2nDMrJ9lNAMKdsKD6A8ez1fJqHXXpagFjekAJ0sV
lxZ9jWQbeKsNiiWmr0SxnY1vrgOM6v3J98Ylhig7cs+Ifyu6HuAk1BgOF+7geiZi
G1c7sEoe17arUeC6dN7IR0q0w5O1mnu0WTk9EdWFLNNKCLRl+L20dpFwHkQTqDFh
CLapA4kYut+Zjf82X4y9zdNcjG2yVwJS7ua2W9DZ8rIS36XoiAahbagLwODwZnNt
uyVmY7Vi5RRozLYMQtHYkiEJcwhkUZxNM/N9NhUgPxlA8uQ0YQbo2f8T4BtdHU+E
im5LmYBXJNBo7ii2Q0u8wSjl3AvEysSFOZagzTiIDmbHRbOCzvdjcHHzmXmhr68Y
y0nlHkwoiImdeEGO1y9DHWYdU3azpFUvQJGjn7bkwC4XehDa6GS6kKOkf+E2xH6m
TIcesrnvLp0MJel5Xgw7P+DuPGXyuv4WqF8pw5u9EVGtAhuxGmrbk7CdHm5x6Daz
ZETfRC3zc8maumGMEbLuTGh8uOFyX00YspbYg6JLvJ6EmbhfYx3YsKzJyTtfzDmR
EOFKq/PjVZCwis/86znsX+k9+05mlOCan1ZeMsnQnNOoBEmnvabRbzH32lfNSU+T
GrZgY01R72Z3F+sueTvSAbWj7rLQgxYMQHe7CJK1mzokuyYB5xZSOAYipsGooEGt
WvzLzm7DNglQ5u6O/izWQtMz67L6G77wDB2/+VPGZbHJ3CwPVcn9BKKPY3SqgTWs
qJTqcZ0EouhBSI2AuU6TcBYg8xPZKc/CGmnSBtmSD617Ip0JbbGQAUo1aIcQyb/7
kayapvroKIon6PBg7RyJKf4lb2n9jIMuR31AuzdUnTsFvaNgne+5MglFAgV7Xo6Q
sNaXwLnyLdx5+ezC1KbWJEBjiUhERJ42WCuIg4yRAkTsxgduV+b3sAMINQLTfsG+
AXEYhzMQHvboztRIklSg681Uoit6TynMkz4CWGcqyBAKoHE/io0i53K82022aDpb
w5cv25VzOgyhgtxHUwjMBZ3B7LX8GTBML3o2CYyRB3o9FSv4PYNUyv0x2e7s06Cy
kPRKOKa4ea0vdJhrjl38JE0OBz0uHeArtMUwkF5vtuAWcuEUlnOHj6r3y5PYL61K
JMc0BEoLe2o3T3lyNQwivSmIT98gelFxoCoLppCtxE+UHZ3ktXZsWlosg66VblSh
5Y96xItLXVGC6uDwB/aFmT3UhDbfGN/M+FTT+gx1ygcu4S5F82IEXYZa4R6NYB+E
aeFGlpL/5ffYDFNJQhPx8hJ3HV2lt8+cY6aehl3g/G+hAGfseS223bs28IXv7sbK
Ez8UpuhQOWwcNPnHalq8/XIgkms4xfv/qXfl/HkJpt0tfZhFTrlNIpJmbCDmthgP
m7bvRj1kBzbrquu4PF/QPkNQSTGdRuK/Ag91d2MhdtQ+y2jkdbSNkhwuqb2w7phR
WswrpjJpndgepVqc9jvcEi2Iifo6oCOCpjHl5iNazT8M8ge+zSArYNXQ8GNeSLMW
AR+e6HiE9Fh+KuRc1LXnn2p6pH6yEdLV6h27jBYijYXrmNeIMOn6rcVmBF//F9y4
eJ7lpmmiMxjmARs8n4afWVR+biiXQZkJVoTAkKu0pVEMHYotacuBsNZUm/8SUbiG
9EGQ9X6btenl7ti1z5hH6o9DHm4pEWuabuNWtRixRe7y8nk7WfJmAxyu8keo4kiD
aQFP6uK8xMFEL8BvTi3srp7p8xvlQHPbksluKB7V5ICeafnNndLf6aTyy3aU7UaW
USj1QYYTpwyEmprUEdlICAh9eK7XojRD4FvIUk6kgBuvb5+syTGcTh3rd01ZVwui
4IMRvuLPFZxCw32dTeSDYsKQerM9d9IIrWBJHAMO/6oPuQN3Q5XcpwLcuVl7GpUn
Jiyt/llrDLbTkveQ9SBO+7PojqiXzajGkImVhEnmbKfJcMoz8sqRaRg6vqa2dzQN
zEQziorxUDmT/axo7+bIccS7yIO3b8pNcWssNsLB/OLUlsd/uSSWk6nhja9ICUjW
dlNoAxzRS0DM/sZa7rpdq8Zy3Qcs7xTve38iKVD00D/0HFeLzpEsijqi8XPCgZeu
4WOLhEIii1PZR4bF+aikaFDMuKiAtBUvH28lgDz8XYlyEy+1rurZ5PatYTVU3MXQ
3J6mFBxca4dHHspfIRxLWRkb6oVeCWjT7q/1D+jIYdB3sPwSiCFxMZWRX/GtVRRG
mREtNN350A1Cu+oItVItoYPZI0Ueq8mmWiPcBqxVk6//N+g5A/bVdSk+OXiDt0L1
Wv74/R9C8IKB1BN9abvsJhEBs1VcP5VPFROrXrfpgmhVuavp6gH7HGM/nDVdVQCf
p41QFXoMfv+sJI8tZdR2rMSz9kN1qcTWeMu9UX65NAKlFiCb2cQEnsxtnyNZe5YN
6/wYSTaZe6Hqm7j4IFYx71EKZMRhlkN2qCHzRhr7PL1wVJKUC7tthPQpTKokcdyz
vCL0QOawMX9qbVn+NyPuUGWAiUKRGkcyiNGmDNsL4Rk7ft27EXdBawVyAHwBJRQY
Eo5b8EUalaWTGgOT+AjwNmxLW22irALTGqjo7EmmmY72bATucI0o8LoMjUC3ZMBi
2i64+lL163aF5xh0CCupA1qXQc/6GBKPtOtU91XfhXRmBKKvj+8Y4FjnnA6WV18t
JtttoInK12SrCO9fQdHuLI8UInMQpPRTFEq+uKszLmOpk/cixMTVj+QU9xT8OMFY
o2du0syc7j4r0SiBCzhEBdupu2cKerzK8Lz3cmCvxUV587b/NewD5QUwRWD8KJDf
lXtc3imVbnIGr3REWOlwh370nHf6dNNGX4Q0KhEe9OUMRHffIsqU3kDzCldOslUv
DdahDCyjzeiqkJyzkui33vCh8fgyhtypWmIQE3JrVpMdE4qHu8oRU9roVVr1DDnB
tZ1egG8bSAvvxnfvKv67shKfFlsb23yg/sdXNZmq02h1xuiF0TQaqSInTioV+Vor
7BClGIMkmGQV6jVPQYHNZueHYy8rJ7LOTaDWAX1V+fE2Zv0TUVpKrVSF9JFM1jEh
+rqGeP0OWDmtFx1er5ldvIpXKBW57/By1HPC/2xcEmrxPyhy5A+o7T3NuKV2BTkY
keywlkbLJb8t8PxxlQwMu4kgfMZLHiO79L5p7bMW8xMaW5Vy20jmeuzSRScR/42y
YuvB5jaoDDPkTYBhcbZ9FEK1sJeXbC61ksTBzApQPsSeO475qFRNEEaj2RZ+fRh6
HCpsOlN4PdYrEjf/d6+msPlPe3Q/NAGe1fI/WeU51bg1nBFtXDFdFrudnWkoqXyd
LUqj2PHmQXzanmpk5/l/fbRBgJKmxwTA+85PRjE793U90+ePLhdU/YVE0bRB5Oix
gHxj93F26X9OXT0TL25rorloD+/on77Lvgscq4d91Mp2b8fAtGsrlHTPXGc6EE87
e2fYtXb94Tuc/pw1xyg1hJCj4oq74qv4kIHt51PWjeu6+9zlwpPNdBlIMGQnqH3q
2ykTZdiT6TiPW0a7pQhNyvVKFkMl1oe2dT0umpAIXBHjmkgRspSuYZgY8opJbGKI
BVbQpcqDcAyWY5jFrMjh6DoGBq4yvGvd1xHuJ12aj5jjUyygrP/vdObivSXCHxu5
2iJkZapQ22SV9Rg2uEcOuByC+HE4IoEVH5sh/SOI3UWlrI6dQGsVxseL0HfkZDLk
4z5A291gTL8JPGhMPV62UzUnu0YVrGJ61H/9WP3kWloqhxXEuEGX+r8/jQyMXhqW
n005tRVl2XwHdpA7y44CM8YsaTk5sfxE4n57YAsZEOKRRSIRDZmjwEaocIR/qj0+
FSfTTCwFlAISJGC+1yanDNgMAtCPwwJWZYI/K/xHWzxkk3VqNuv6kFShtYc4RgS6
9JTSbXZ6Ek+0MQQAkWbcxfXedZsq724UVN4/OFrve5Ck8AV6KMuhMI7g9QBvQclv
6P0xPav7+3gflVCZ62MkA74D4xoTB4l+MkyCRr4PPuJGe8SbVmjIxSlXZojnkQEc
ohcGntvS6yPa4gYD7ojdBJB/MK9Exp/ZRXoARtg20qAWYiwDpzO9LWdK6ypn1mRO
oMN4yim714+dAIozM26t3fsKgWHt9xyq0Iw8aEaiYOr2J6T7vU8ncU74QbcEk8Lh
EUpnZQVu9LnleeS5wls1c39qvyOHCDuLhaNrHFQsBfV5bSFRCyyLEPA+hdCwadd4
yuW/rLVVzt8Z6h6BwqYqTiKdLDkM6aklwvWpRJmsOAktDxKkotPA+SG/lY86chOh
6u4saCpbP8ldYWoQdqbnawmwqj3mk1TA8S11T/Mk5rlID2adiPxPmEmOuLYLEUWW
oMbpIhNtReyxEQiwSH4gC6xIk4x1A8tPf04dpk4d8lDAR7GafVPYKP5sUcVMyzh5
JlWGDMlclysoXvTLzTtc2NatmDspXYzDzijyqVoYJIbmpzwKONjE9rosfFtk2hSM
OLHNH8+i/n3EO0mJb+s9VcOZJvT3h2GZQ00u5IZyfT1jYWPDCqU+YLR5Ae5wq9TA
X/TdncLD/C+tVcKT/bZxbznl8W64p0qzGT4c5ngwPCXi6xu2NIxekOV8E1ydI+mW
+/X91JyQUtTNJCIhC3dyRouhZTgg4RTmrYIZpkp1V6Pc3JUVPLJH42+47tembpbk
XGFehVYTiGeZc/MCBFTIRVamgjt1Syuq182O3deqq/fG5oWdIkqDuxyg+Um7sfRk
2C9IWqRCMhFXAr4++i5Z3J2Vmc1EY78djWpETq1dUC78fhVrbVvkymcxIoaNdokl
ixnp23BfUx5VPWXoWy1f25QbFDmdieqIlgW5atzU3bS5zyMgPgdL4+P/yNfxPncC
GGtS+CNDwJwt/0JIjUHTC3oYwuZMhRxca/Nydp/T4k23OfKS4HBkgRfD07OhAPi9
d9poBXKgHI7oDfQV3WAQxu9JPd8WVjSmtG/GmhaucU0u8fGblADWKnnx9zEn333X
zmMaUIA5opiB+ewSWWcOyifgAhsndYhcv80SbwUmGgBYZi4Ki4OlWjwjcihv+Hk8
a0PcSR/XGs5eD/OvkdrKcF0rOQuALBVoHr84PdUY9JWCuQ+4iRT5qfKdE3e8z+fB
5R/MotvRMhriKvAf6OJ0LUUPxs30eqi6M7ArUj+pG8eQYsT6hE5P6O0vfAcKhsgh
Gw6lGVlmWzvpjvG/ymIRXoodatPbxKB30zIoVTlxHcEkUDaFT3GzOna4USh3zv3y
gcDdzLvYsqsqagEg+dboaegOUnB1LsdWwvCS49U5ZSRPub1usi/EtsJYvshMEz7F
xaPbPVSdL3RgKrVpic3+YOgiS/kCOqGV+V/S53DwwYcclu2I5MGK+uisaxJav0IB
JD4zPIZNx4RX7FSQ6TkXnQCZ1iFCA+dkoKqa+EtwtZ9GTeAt8mMjhXblEMafwr9+
gbCRzo9bPv6JXr+4oJq7JmBILSrzhnvQJSTPW0m+OcnUDlxycQyF69YmMPsVVLyl
eJITZ0Ws+eig+KSE/EFLXrbE4rwiXzE1LjjIUNL1egW+mzxrxbRpBW1knRD3U6Wh
S4jIL/yMlpjV5w7M1AcKPaBtvPp0d05xuNka4I8UsLiJw6BCRexw62196AgjD7eo
SCelLKpDOzleNqU6vJLQXI5vq3ZDEQ14unfxn9XdWvHap+SFCxuiky8MDl1cLbcG
mqtVPjWKZ8qYoaZvrKnYxC4RpCqzuBmyXL5mOL8LgFeK+QcrTWHSpzVXL4ufExsg
gAoMGDzVxVTOXCtyTqjoGkWkSTGQ5YlVPyHbYNdLV17MmoSMsBp0Y2TH6RzjZtOz
pyjIs+8DQXoPJt9PFJug84seRPhUaY5W/MCLSay8RGO8k8lLsatroW/Pnido/bck
BhNaXj1D/IkLJGDhtxSiAnOEpLx0u13UXfFi4mHoumQLXWloVmUA+U3WBmhTiogL
OFePGwyQZi2eHRroYNTIxMsNSGjr+6TwteL1/NJ9zOaccxc9q626q/rxl1kf3yRH
/zCkmlIbMBEpvheqnd6dqFq6vyDKg9QihhtvkqxxN87u9Yl+hPCjq1ck72px3+d0
KSACqFcCrWeDHS+EMLwAGN9w8GSRtJvYJqspzLg2OPFY4nJRQ8DdUoJlYGq7Vb/Z
OjNEIJjTGVPuIwKeUGrh6ROA+Rzg/WWx7BitX/m0KAjG7+aFugQAzQYfOsZ9sc/H
f4zIxJhzHQfdtpbvQ+wg7HE6a8IZuJY7WqFt4FBj3hakKs189toANj4WIoPw7shq
N6pCMxRLifQBn2OVQjAI3KWqJxlCcr8gZ1JQZGzFhr1DMVa1QHs7sv61BQJ/p6iw
fBWPRQtvmOyVgHfRbK/Mlmn4Q31IjbULW/Hl2gSHDH1tK9yS3/XtA2khuD1AA8bI
oiLqrJyf5Abasn/Nk++IelRtiHUtUOBjVJ4+PfT9Q5yHf9A+zL+H40T2E1w73Tck
M8DFz3U2aRVh0bYXUZtfYkGypvYX196g5M8TS9RUHpaRBCFz3bqiXoeie8BsAz32
XzrWP8Y0yhaEeMxs4q375B49FDwqmP8ORzbDKuTrBDg4PsAAXPAxxG0utcQkhvYN
NsIG2XTGSOkuvZonZtZ/NGhilln6Dd2Ume17PczNvO1Ot7kkkiHlZycqhki9xdkg
uyZeoDi77cLKWJxmTEk2gpOWXffbV7REbc2K5grhJoyPg5K2j4n2j5RnjE9xHbxI
rYMlyI3yBZrzLITV12AcuJ3Y9Deg7DaapAV1OWZF8qCn+NRVXrvLOIt/4epUNM3Q
uLsm9PWz+RaGBmxPpVaKxQLKkTTY1fO3k3P7jnIByi4A2V/Ip8MRJLbfxTv4r21K
K2fe9Wj/0rUz6bq9bRNSpujC6BIiurOp6Ah5h35HMnY+BG+oXlXK2gkzfh7EuxV3
7E8A0jVAWAci6yuxb+0nHr3uUb5iIIGnuIHFEJZz1MV+mbg+RIV3bGA/1U9ia6/z
8At7o7DPnJie4/xU9XwbxOmWIkTcVb9f0PXqoS795eT6WuBXwIn6ZSxL22aSiNDv
L7R6nSisuYLB5Jb5WK4WFS8gAQO/tBlRbn1kGWj8ftcHwdeGuTERXw9TDnOUpkjK
usBZEDvzWUDRKXw5og+B4+Dfq5kYgI5RzLNEONpNlKm9nkXa7uQTbVnz9VYqiV7C
l5IimomQTMLZh23/5jrnDyKyYEyCAJPS388/I78PMSismlZ5qhbKfHqlDtwud+XJ
0BB40zapSRm9eXymxRIH5Y8JjD9uiGIPR4ogo5T09b7wk2G8rUClcB8P0T4A4TwX
EVfvCwbJNh5d0i3wfD9OU9Fnti1Y6jP+7VlLi2X0UdQauwHHuyqrI+YpMto7jYJ2
5JKh9nAE4zdYwkBolcOmtTAhAxrmCuz1tHxMcEYOJ3UunhUc4uZXPXz/PEv+eqw+
bX2M+BC//G0tbd5TrKLLuGyvT+YvYfg2emfqvN9yiHQlGd5T5KDyAnsR8AjbNgyU
iE2hJIOVpAbdX9ZWzncorIPH/hSMY5OcamZ0kd3DRresy5jWz2DeC2tUK13o9zRj
Hphiw1NNjWmIfBe8irMMs2tR7ulVaLOSs195mK0OQLwrqdfKsxrBDdTdkjXI4L2m
qnJDlwBYYal0mx7zQBp+1FTXSCKGWPzbPB1GVbC4BRx6/+6G/GqYNKVBicvMOrJn
9khJ8n0cv+WgMHWsLuT3Q95BGM1orekGvmOFaQUB3l2hPc1AvQLqlOI5PJfKv6qx
2tDk6HGvKBJAkuQ3BSXXIR+pnBKCM1lMvFrSUuHGDljuSnhfm+nU3Vc3S7tdOY3z
Hz4ymAFuZBZfkcy+EkZBnNRkUEaYa2l2lDhYl2nZ8lq+DmOKspIOomSpCQxpbjZo
Pm8tZK4LQMlnN35hSr4hvhOCDIJX8IgaPPABDbx+CGTcjNmRI+9m0nsS3YL6C7Lt
z2Hl1/g1KmvTw/75njLaYZdjcI7qfOTbMxhLbCWMUjGwwKZF3LpAO02Zyedv/T8w
ademj5xZsw812Kb6ySB2uNcf1bmYLPIRz62Y273t6E22/ajHI6NP13NmI5xwBZT0
gRRzegyDa967h8GSgRuQ8FT32ZxRlo4Uzdv865hjcBqAwgPFDZB7hSIGvLLDjszV
p5dvMaq1/sWPXMxiOW+FkowComfwwrqoiXgiRTU6MX4XgPZFO1tmxGaO8Zyh0DR+
znDFYn9oPPHQiy517vgXeZ8QPDT6MwqP30S8jFq8pq8JytubqfzwecgyBLamupHn
9bd+2ISpow7P+L0ks9s3sY6TTEYIGg3JqFioDNAPaHaM3aZIElkd7V2uXrH+P3wQ
cHWpR1PC0uuCkOKoFiMMUDa1nZLyV97iXOWPPaySqhv8Edu3wqoXEofk9ypsV3MX
3ely06bfG4LqwHogdwyMrcPRA/nUazkkPBLtiazqUaBltfWYbIwpq+fg2hI41q+w
j9wyZkT175Nt7UPkHFtpW0ekbPLu1Sp4s1eGbfIduIx1iDG6G9ajLdGxUrp6Us8v
pXxyytpX32DtUCJhVsK/zzVI2L1oVOxc85iTHAdNzB9BNwTaMa8byjLlzpJvzB0B
SzoGlXOX3N3DOJYg+4SY3kDQea89VIpfymCxbBfNyCVYzVYTK7yE0P2kzkUGDKJe
mWGLarSzd2EBMyo9WJ8MzvOkyY/Q+FQZGgX2Ksmv4XdikxK2/8BaaXZF6Jww5zAv
qjKWDU2tnKbI33eaRHOyxE6IUSTUYcj9El82VloIPB279C1des104Kv2WrLNlsCk
LJzh1z8iO8DqxOVTDW+R9B/EXI0CkSNyUGIJWT68IQy9wWxOCkIQqFks2UYpCIR5
E7puQFbYUmXNStNpordM74f5V+NjDKqSu3SjjAKMMhAyfXTXbe80eG28NvzQJA2H
oKtH8rR0C1KA/+V6SSdgGH3Gy2QLGgaSwWIoqGhW+r6VvUFSK69wSch0qj6g//3Z
FajSEVSS9xwa+EQh0DABaYQq5sNzT/36DXE3ClNvkrsodAx6FSSaVLqGKzO1ULmJ
jkKynO2EJwhm7jaR2pKvH3awJ4PmJrnsohGs+PCXXXa/VW77VdPOAxoXiGg/CDCJ
KgSihy4FraXk7QtXfX/6FxJfFgzGous1mNDkjD+g/mBKy1MSof+H2iKDJJoUaq9s
XQiyM8cSFy4M8i+bq6jPfhlWPYfXl2znxGJuCxh420eI3Gtzx7DkmVmcbDSNVjAO
l3O2S+vsthX7zhKBi7YTHYS62EQI5i8/TPNGKsxGhBMCb+GCZSVZYlrCp28bkxle
B+0Q8ssKo6JnvSo4onFFlRqxE9oxLkevJ7OmvhVu/9G5q6XRqR3QSEsCraAYERqz
CXyAz/wxZNeGXaiQ6m3fsavtXrQ6s53vbJhZJGj60rQ+GrDYbXFuziu61EdPNd7x
HLZk+sC3nlfC51O6vo9NOOaw2HAU04N/Kouv09luIEk2BZVZbtkmt3oAn9oNh5yY
S0BetFTaBUk9SQ4rtynQumulWUX4CShcl+LI0+EiLOX7b6EtnyRTt97wDKfiWu8p
7F7nfB1MAx6H+qzrw7FC388W0frhd1HNzZFboFnmu965k75dlhmIB6nLwgDgUHLL
wZhD5YUZGFPjhNYbvbhvQ17bvlEopYWtdh6weVD4CA5cUCFu7DrCUt28CSVQ+tG0
HFZ6t2UL+tJR15/Bovzm2Zs6WxIcLD58oRjD8ob5guqvEyiyKmPq75bsWL4zvOSF
mfij6nqJu1M30S9BfckjePaDZZRaYtdEfyld6CVEjf2zHttYIyZsFRkIiUt7lHLN
mKlnWeOF5EHcKfjQdbq6ylfnjLSQHI2BPfw4HiUXULLrBePvfAyiWmfHkJbe3R26
UDTwnqFKCW1Nf4azS1ZU3Bxnbhvhsw6gN5ORTi3h2neC1F3fSbwibV/nzZ/hYI26
BQ9ACzknPwGPijr+bTEC8eBYOhfk8L9BvpHHeLcDiPrdJaiYLfk7sSg4eUf62SfK
nuG4XMvX/wQpAn2LbhpI1Z+KDG2hwkRqq59g6VrmjdoX7Ka0mtAaJtSgi/DQwdo9
S7gaLCOsc5X31SLQMlvD4ybdbqQcmbSJ/Y3sacAmWwlsGzxB/qzqAIPm+NKLO1DC
DtjLEiulG9a8tpdhxOHw/Rm7aw06Eu9Flrbw0XbWTDATX9nrvFoqD4R7X6DE+NLh
Wnj+jeOyUDZLsC1Xf82Cv3Mu9vUYK5pyLZ/c5WfiBQuEUzRp+n8XHOcQ7DRrRI53
1hzIEOfPxpe5lo6p1FVyX+d0mj2n6Nlzg4WcGfdzBYtNdaWHBuqU9MYePiEWSnNV
vthdjuELG3FxR8Wt2HqNUkZCimABGebdiL/eckyCTILImKPDDP4hggqoJpVLmVBS
QxWVChS6S2bGWD0dNg9vyMu7+NZ0zN4dpuQgWH4mPX/AmLnpT7kvx0/LtOXg8Bcc
tn+s09iEYkfj3+PuKcIi3NBGBZ/nlL4V0Bn7+z+nSwRSCzw6IXJiShnC9ilD2VYv
OiQ4vHBcKUvGqzZBWno2A13Y/OxCwb48ir0ZlItmLvY5DNVpo/LIbbcRyy9MHIbX
McfyJCRRD0nukmdM8H7ZMvKRWBSQxO6lP/eGB/a/ZEdx6R0CZ1yMU6pmrbUep/fD
XuBrj77C71yo5aOFYBl+kD2iqCse/Gj3NN+YWBxQOzQR4tQJ4F/ACVYi6cfd95Xv
ATq5KCaXdrVDKL11GlvfBxjDRpHzXDDdqZgtbg1CzFihGJYPAnnYxk74hSvRRbmg
MZ3l54b4NvbssBuJEJuo8EEfhahzrzqA0bnumEl579BZxMLwQVIn1tZe6X0APFVH
qmGA5p1B6jjWTQ6TTCctLd4qPZ9T4vIhjkBCZCr9g9uohkgbbtng2a1TogX5h9J1
Bc3KDAS9fE6cFqTa/HI7QLx4bjF43Yc7WRR6SHZkVIRsml06wSKWdBu3lquQs5Pk
+hZDnB1DOt0TVWX3ztHcYmUk3Q/3sTkJ2V6oYr1nE0v+eaPMnTwzHl92EmJV8A8L
SsWxHz26hVudVLM5hqJ4qcaW4ypG2PaiXXjUSnsJYo222Hi33mKGxElBX6iNSECi
AoB0K/X5rtTpaYfVzlZdtNQ0ufrz5CSy9+qH/33OuyfTnAdchtsksi5oxz1cJdiM
VoGzJonA+cD2pA4BjOgycepTzDuZPBxmr3Itc7kepms1o++VfUIY0LvTKZqe9sc6
2saV3nD0U6BS5a9b2AxyFBigQfhtN/Upd0Gtvk3IiDeeR7wD9E+/+zYgDv7xDHBs
nIRsi/xSxUfvMrJ70S0MdokfCtpmI5v5JSPusWbRA2zif2xc/SMTKWUoQRO5CNm3
BZ4PxkM5Zqc6Abv/FyksX3InCNiO86THgodDeCajJya27OWeXXbgOuBBQdyB9h36
ienMJYnmg5OArYRRmJ1jRgm396G4UKIpNLmq7DL2v5teudXWlbQXkAhMlD+QMQ6U
g+0fOBmA74X1AkcOQFGsDOqqtozR2J1wy2INMoBvIhFHIpFKLIN56/NavircNBKV
URCNLBWPjrC3Fu/MNUMzjpS8XcZMuYFdlpRAB4CAn6Eh0yqcFSuiaIqx2pqaOnlR
XMe0HoCJ6fyVfyqteRjFMh1tM5emQzAeE9pu5uzJVmepXSWBpIUwvgP1zkaXaZ0n
W0f259bmE9ongwMSIQlcSF98xm7cS2Pf3nJ6+UP9wnpujp8PADdWeqtXwJzG+xoa
HiYsaZG9iXIdLn1ZwIWMiniY00oOM9AOi5r9leIOkb9OuMMuzfQEEmAJq7jpoP2r
HfpauWfYoz0yAn6WkyV8bxtpOPaP7KU8gNT4mhbgrwImrvJMrhMzxYOfSh5IDP4d
w+bIIMDuM4HROZUheZAkCgcBemcfPCBY2xmvAO/CTw32sKsZbFO3AI/JfrD60AD2
eBGrRdrOLREnusvPVgYm413ZO5MF4v/WnsWCUrzQeItcQ3JyCdGi1iDDr4TElL3u
TEFk1MsvSs8fpHsAhi+an+VO2jUl/hvff2rMKxq47DjsFR9/InN2Itld16vBYebn
qRcTYgriqZTz42v0o5/LamhI64za/QshSVpBPwzTxUd1p5tsDmRr20eZMoDWK2oO
MxblRbV1KFsZeRhn9g/HuA8llNkjeDJDhSnOg9BW6d1bbP6sPYU4rUAeuHmDszwt
HBHfq/sD2IFNRkuZyqlUWGVu+uZnFAFCsygOsy5af+pbIaQWHdzKJ/h7wNSCduSJ
F8OqlU5gImdfyH5m+IAj+JOlvsmSmpqb+K6G9JIop70jEATyCwPR0sZqsAHG+apn
DrNuqKuN4xmqoBjYIHHAod/axR8xzr81ZYWislrOnYT7ZRkE6KxtGJBcpYmBvEOn
EBY+a6JbJUUrbNr+rxZRVEK/5BWusBp5YRWme91bub1GAihqGTsYWCxRikrF6t87
7L9SSSQ5Ee4AEALgRQpoGCPfUFQkfmpFLiBzUAVDR6UuM12jEAyOCfkd0d2Isw80
xLN9JV6R4DLtoPm0Wsj2NwK1TzORnfDwqQMCVlVLupRhC2tXn8CVZrcwHzvEic8l
iMk3nDJ4r+gAQ/HC/iMJh0UH4LpAlxDjKROIo2ScerETtB51LahL/J5Wra1m3o3w
y8Xi9yQ+OW3zUmPKxOwNob3QeI4KkXkn9M9dIHdhc/u8klyLE3RO7hDPX3S7kDZQ
eNddWmiXDhVWKFtKQDxxjVu4Cxt1kXL041G5XCmWY27Vj0VX3ZZ0L+b4FVhVdAcx
qDngTAGQF5zwPtdxcLDk6ic72zx4n+2SypdK0zKII9gyPQ2pmxC/79P3AbXpY283
vEwtU8+AtaRUGW3sQWAiJ4M2LAmS50ypaH2d0wL6VBLUsrJzbFvfc3mlfTaVjZIb
Ei0ekodFunvmohxCHi7+ZbQKP7TQmltIv+zENAr4DTJ/qNmQGmOL/ziEYnbzcFcK
Sn+QV4T/RqwTwnxr2SNbdLuCPLGXgIFItCHP/IIA2edEtWzZ8mfmgYaKk3PS/AVk
dKOrOY6RLD3WMv2XSL3+J+0413T4O4+yd4EoIwaUtrN35n2Pnfk5VzkAoStPAp3i
k4uxxO1eFuDRz3UfhayC2ftpUQb92gqHbN8WIP8aQdQMY8eBoatK4wKf3pIXVZ5U
CtAP3RmEbttjb45KJ7dwKxvb0VRvPF+oQC97jALfoT5AVfunviTIiYwaRidooso+
pJdz9/HlfrTF0lw7MYaaYQ7AjiJ2TD38Vl/0EZGehHrvkRGIpUpCkeAGVSOi5Bn8
d/oG6Lp17bo6jWNvv5dgiK67nWGMj8s2lZ5oWsCrpV1v+0uoJnTGV8WKh+YlmccZ
Z68JlXkSfaoJgdaBkzqrtySa2FOSXce79G5mPufVBuopslEMJszud7KYDv10L/gT
UVSG+cVvQR8k5MoOxUTgK/8dtSRk6STq6YuFDKxT+RNcr4LC3op4VgmZK8NCtKbg
x1nl6Br4Qe9rMZ4je4+Iv+yQ50iFXIR4+rL0JF3uKnCTKBMsgmRFBM0xmlUC4c32
4CLAyOs4z52YqmRKThyGmTVsf4fJ6I9qfN2/G708SJg83o35lv9qH1V3Zx4Kzjb8
H5ltME9NFdLF/6VvAhyYuEL82fEFdPCKYCD9vpEdejXZKdC6me4zu2HRqUqWWTOP
FjOEqKohY30f8bVXuqXUdXPLJs7RS6LsA61ip92biG5yNC9q1mHGh3lUxJGi/3uS
HWvSIP7lIiuBGvR3IkuIb9rcYM+Ye/ev7UPBUZodpKTNVw5S4rqkxWDGo6obzemd
55vlSjWokz1eaEoJ5BSJ69zSdo2UOaBdAEGJt5xpCEGXVcPlDFBTfN3/VTLelq/g
N5ziiKXcVIkPyODdcT05miRqUtc3mguYHhIYlk2GRAMMXbka3RodlG1IHqXM6XvF
nGTzkIrSaZhgxfgxQg4B1rEVhA6/gpMGF/4ZVwg9jFZYNwPU3ChrfFWoOk051Bfz
mrUR9WZp6lR79dj8OSD4lbSn5WnYd0xo1ycrBn+wJIgE01P4Sma8hei3/UDyW7QA
R6A2KglzJrjFBV0ZlNo8PNDgCOO0ozmjPfxmPTsCku8/0zHzEh2fbcTtv5wyjmMU
texKfOpACw67GHuNToB6sOiJIPLLAqG4kZhOptOiwDVDAyHOVA7JfGsj7I4jEjsP
SLfMcy3b/n49AkQsOWLUQ1KAKa3fLi2kymccSGVkUcFLl7NHJcINtiGmsEDFNcF5
5itWnCGwCM2oB+ruJ42jvR4WMc7FCTp2Z/++eEDAjcpRUbu1aK8qPfv6nPAh67td
jQWiBwtWfGbHlki2bk1KkLwd0l8oP+E93ISM43hY35cRDxeGFaQQzAFS31Ed+MJD
8pmuszM0p9r2c941Mp10s6lxrtsZTla+AGysTZKkAOdfcI6Lvl7EYPQvemk2MlQn
b2miO09qQOiM19pSXGq3vBPdo//pWvfvzFE6XmqTq/AKJfxejWc6BNrZgfpw1G8l
Iik64XvH3QhSyaDDcFLXPsLFPIdjgUOeMBBswONI+yaMWbGNUwVj5OGjomhqCZSk
Uu1+xzplsL87Xt/oczF0gKgn7MtAHUiePaDxPHY8stPek4J5rj9RQ+/876GDAF5h
z/HXPsgmhOlY6Iorx/TMkCXul0l46XSJZJzkc4ysvZQWffganCSiwaZArxPLwpg4
LOdWrEDnnAThA3ybX6ousnajm5e8yAyQbmbvfCHzel9BWllLjpx+lfvyH5YFVcLv
Ke7HDc5kqDMGucmtAk7tVM1Qq4g2u0+qfdX9QCK7xTfSQcTgF8jdi0t3Kj/yfVR2
jdXwnkU3IhzPBFVkxo5QrpJEfKj2BES+lLwyr5MWO+wML5jsKUHML2t+LQPnrHKo
MLeo+bQa17ZIxg29rZ9yKPiLSZUlC1NyyPPccrwkJ2fFF4Rpqfrltxp1lKplTnkH
Rgit2uee66l4nvitdUB75vUjA4QAsNdTaXzSIlPFDsAL0rpNRDpxUTsvjicHsrzz
rXPnxb3HnRgwxpi2wOtGOKNRzdRV06ZsP3k9FdZqor4MJHHZdo0fiifk8cHWck4l
Q0GHjP8Oc7TZkqRt36T6ayNGzjiNs1Lxr/79roVy8y/HZ7qfx3XkbMym6EwaBiLX
lqHJVWzlOorPVeCbuYkVyzJuKgeNNLtMZjhBQTcGjW1dCGpDWn9HE5mn5sB+jAxr
/lrY1W1iICTEQxwpSE8Svk3LYZ0tG9TEVsTYhCUpg5hauhiDxwjdsCCqkUpcLLo9
AK4DQv76iaqlnzON7J4S95zSTSnJTqzW3CRUOmc8LJRclFQvbQGBdkskRLAWlTwO
4NrZWUHL3rb4MusGIveIWXkob9fr/7YJ5M++m37WIclF7VESWbayoHsg7K2AJdnV
AIh3n5WwmotvoRSIBjv5Z3iP9ptxKRoWYXwuF+wCfcotgBoypKT1uV2Xu4bgK7Zi
NKjjUy/f4lIgwZQTg80GGvigq0wVN11awUSklhrO0qvHXUZiEOsYeickR7iL0Z4Z
iLeUghOg4gERvDwl1Tk30YDhr3wobVtBatGutdxjyfckp+zQ/JLjhqzIOkJh7dvM
QRrmAgcPicctgxH1qEXXV7rOtIVcu77rPYIYazWviZL3IiTTSUNFxbDBsdp8DtF+
ElobNcwkip8Xct9TyK7ZTS9ZKFnMsNUlmWFYw0KN0/7su9tg1J/0jDR8qR2Xkniv
zfOr6M7Qpy75DOMtr3QCcAf3GLA91gHiV8wGIhEV1Bf4CIB1oJX1c64QUHN8PeT+
7olRH7t7PqwiBgNRuEMljs2RvC0LFMgK0dFjJjs25y3bYBFGb/FnwKfdVBkkgTRo
uyd8xA+oelUBJ6Ce+IpGPKWEEgwlm7FfBpR5zlmg+1BCpJa9L3yAK3ARsbyUgJx+
1TplTMQezrwnMHs8G8+FNP38eJO90sEThU/bkGNRMfsHtr1DZgtqWrADT6iongCY
fYEGLmaQFmtqfh8kBwx6pUYx89eAi+4nyTiWigwVn5jtEPdZ1VWqRaGVQD23E5bi
RnnJb0EbX2HVb7dFw5J+XVySWN5Y3C/q3K8EYqLfUBVPGTt9IJrFUo81ONR0SnMo
ibGkw3ymgDZv/R/+z+5jnUJ1yHUhUm55O1kzuNiRcN5AlWeO7nsmOhYvV+0lEZFe
SYnITJLVW07w/e1kky9OT+OrkBqfn3AQx9dSmrHg7RRFSyXfhbnXC3Ac+hlojfqy
FfLC4t3DDQHKm3/vVaVVlaapSC0EDNnvotUdfltQj5Ygh3m77LtLmQk0/V6DWGML
kMLgsjlgPq3M6p2wWR5ER+tLZBAsrrTBDctrbqYAO3N9q1OOTCv7I3YtORKVWkY6
Q96dcCDqExAxX1XSEHmrSF4OAVPiQFodArqwI3rnL9GI2Ag/SRCQmZiKinYcvrXA
qcZbjN04o/GVOYCGlD31G22KS789mywGMSgzX6Xb2GgoE6J5GWrOUqvrMZcyjCzD
LAd7qC+q4qx1lquTjyd67CmT0wPrv8SXDAmnhb+wINfTQmnnln2fNd9ESwaOf+s9
MVkU8z5xPzBUeSsl4n2hyGGvoSmDWrTvYQPawfoAZ60S2PS5VIkGV0AbysEnp55m
gQEXlOuN8d2GArHyuQ4IGs9WQZP5FTiG74ZUeyrOgkLGsd27t9cz/Ek5uiKjg8w4
A9MGlfb+W3dGdWXcQt+COXl0ekckWtdiBaaTdUOBlRGz1/Wm0ngnXIKsEmQXAum3
Bp+Lo3zg+cnw2OgayrL7mPwq54So04Yu5o85ioQVBPx3ebbRHJkcOVVgosvpi5sV
7OIEenBxLl9jWZj+LYFUpNmay1J2f9QKSCAb/VCxklew4007hkIj32slGD1eEhaI
hnVFrzeRXxYE/q7q9GckEO733Z/AY88TOPK8do8IUcSu5OrgzV58FePtYpoXVjL6
UdwDUxa0GO8eDLWuksDD5PUxzSpIMUwBuSbh4FSd0uvjJ1YBvb1xv4VLD2haOime
ChuzwsOpD3L4hR//Q2ZX63g0f8AZ9+bsxpyFBzrKjTzFxobCa3GJc63ifn0Pvys9
pTlK1NkBGYzC8XNkoPLuDxWtp3cQIW5MxlYteujjHg7t2pqwDg/T2Oj2ww0BcNS5
KzGfceqLIGsTWmTBWd6jyGJc3VLd5mtFZrF/R6j3uHopp7neyN2V6d0B0/WmoU09
sMQDRqY/kR6tJfEYoura3ktgxhaZGlY9OOu7m0HWvqW8N2QqqYmhWNt5isF9vupW
hnTk4wFUYQZ4YrF+qSku1fwt1ctwcG24aWzE5Z7PeFL2013GosgwnpCCYa5JAuAr
LMsGD2GJ2xEVTizDlka+3HBlHtYM8JJ/GnTtkdQl1YKl3GnxFYRwzac4JYYo13fd
L1aEpdbf3nQZ23tGVbsxiqG1smU5GWuiqwBqe2bacnzLKnCCy/tahniBHxd+M5SS
WHRGoQ6kHxnC4jUVOJLi+/X8jMmFQ9qxF179uopeta3DBf5CAmEqjUfp4TnI9poM
NpFyl2e/pJoSf4P2ieq+lz0mnCbuBFZTjPKYdgOd0edMl3+VAND8v1bt5aM0/5Oi
scj2URDnuyY7sMj7gK9bRb2wiZRTskdfFuf0YA7V4FIHElP8ttI1C+5mn0d4NRuO
NEwTnA1vsa8mhA0vo3bBOlvF5I/nrBrs8FY2GtDGH3cB5UFh0/VU0DrKvASUW8/D
E43pqM2s21VuDT4tEbcEJhdtfKYtCqe335VbfCu72Uz/Q4k7TBFiMRl7fT78bSP2
m0crCUNrEu84qm2YpRAX+bHt2Hp1kj/9h6X7/07QX78I/SgYUAV7FcfXuyAvLH/l
avEhMvE6UFubaSmz8KBie6jbWyViF27Gyx/7zlQPTTch6OJoU/LoBa7IvSqA6peK
oq3e2KcamHpKoeHfM/x6Zsx0yItkr41UiRf5AJDmqZVCQQkS+siq+iThbbNWKq+J
nrZXXMkhCYsw0lAzodAtdTqxQgWtzgeqntxeUdzg7/c+di2NkNHeyeXKHNbRWaGB
qz4IErkAz0eYit2bFP+2D0fU/cGl10YWx60qnEV92HzlIWKg2CfwGb94pk0H/SNV
YJf1L2vmAJXokqrSBBby2z9QHECb5Fw/siJOl5MpVwzfgvjBVI7gSmboWA9qJWdl
klID8h53VAfwIX+7QWXW27GrUHmeY98lCLU3UWEFHS61mbbCVO5YYefVq5ui8BCa
YqKqZzXAqGsrgV2noJ6rKRuSJN1iP7iqapYiQpI6L1PJciesDOT4dEgIkCp+o5Xz
5324PlYFMmg8HRE5uFjDxfWNlisjfzTQO73DkSBKdZqaxouxfIjDynt1N+fMl/IZ
IkgxGT7E71f0bUvY0zDj3qT7AmK6nW/UIDeRMnna3iMgpRxjaWoaOHH5qzE01Wm1
MM1Gi294daQ6fu15vOWJM4GUmJ1WbLfEMEo4deVvsRddOJLsvNk37zWnJCk/gShE
7fN0FstZrxjz4ehgxgmbs7WRPMLcbUAFHVg62C8Com86RY1UQnscWvQjx4Btf3Jw
lGnFGRQFt0XPSWiBbbdXOfwpqcVe/aFuF/hzHucRxjBD0+wKn6CKoTQ9dQ7wlkh3
HpR/byFe//jVrWMtzLWiaWhgkKur5ARasnWOQ/HkmkWVpVFjQ1CZlLTKFnV24+zN
ZyyKv6s+Y+9u9KtMYhIGMQmyC6oCDqTUG9zDdZUn6slDBdm32PmIVaTFUAUqnm4r
CEgQ7xhH0uh2lgveVq5JEg/i/CgQGRPLjn97wORhdYZLhiI/OOgB5Agjq8fuKbiP
rYtQRLXbTcBpykfByJtJ5aQfTgfsfdcCwaKkvWY0GaHzNPtZ0PYsHRgvxv8XPNiH
MH7mKPHTPziHwestOxU3yg6u5pzm6QaVAUx3sOHDo8RoIvSLHUOrPddRArvre9DA
C9vfKsc7ZK9Gt2OoKBLe9FPlMq/aPtkHsaz1ccR6qnds0oHAyc8bPilztojAeRyc
r+CgZ2YeT3NNYR/bq+ljmh4iAakK1F77XzYVWUCsKgBcEzjFs3zYl/1vMQJf9DNJ
tOKWARZW0J3yB33oMRMUdXYGn1DVbML2EXsfESu3/D7VtqLXQLZPUXxgMmmzXqVj
NYV7BtyGMrKduWjVj5YQ6OEeHyNClEr95d7NQdRk4z9FXqhVn9Ky79+1eM7BX47g
2egylRvTD8sBUWSNCKmwqGF1feJJsIOBpoorPKk9P0o6fa4KoQnb6Kg+v6LnEkOt
QT+SZakTp+468o3c9LAuddLPYzZvkP6sRKke+bYc81jGgiQHqsCEqR74u7xoJpob
uwMG2o4zXGE7Rs/rnru2p3nuxZdmu7Nxgyb8HjXh2ideI9eF+867WYpwHkos0X5s
TGsSJCC8phZ2gU66ucJcYf7I1Zp597vkAsW65bqH/TixpSxLsYtdHpsbwNIhoR+y
ZtP+7THwntrtCGRFO6gP1Vn4j7dC/86X3JU6F8jcxWdmlLw5bNaT+mHEipM91Huc
eRQKmnJbb2gqZKXn5hI6gb5DJ8ylWMRlDH45Jr6eYhgjH+H97fLu2NX98kPjghvC
Z1XrpSkycM6ZVEL1dgjEmCSioDlL8VL40NyTvNfcifh6ZcWAqATXVMVupFQHk5H4
e0GghtVSd6dCYvxLk/u+w0rciVH2Q5VKYz46AQ7+SFjM1/SNWTAND5sI8aKzLIDJ
I1n8qyWs76dJuTArKLdECj0ATlMYYwh51xrHfGcB54f9sVDqj0IcsDIxzk5aVC56
YEJI7/61d5NplowJkmDUDFotSMGCUuiaogF++PTMujjkbM1onLTbMx8PLjGxLfb2
y+xB4q9W8RaYSMOBu70Gh01eEdM/g9FVt6BbebLkidmp/4ST4xzKNPvb3Q8irNrd
tSlJUoIhXX3Vn8WX8E4sUM8DgG37rr9B8eWKafdCs7rpUeFi89kwICRS4DctXRkO
pk4GOjLY4m2Qh3Ej/GzwIh7vF6gjthbW87Ncwhb95DCkAfoEohhQnwhUO8y2P9CV
pai8WrQEZVQs0fp65hjUQ+DJ+SeJ0zckwQJ9VE7tKdr4uSOTULyIblUAGVBPzFmq
C2ipOUkY5lJx+GPS+wkjRvQWLYLgX2SFqe39VarRH2YTqVlv6V3GMYYrWsiLnJIw
KQIgxcV3v6LpsmHlFKh1Zy2oAdkL1lUXt7q5s7ljpxkhwh1KSsNqvoclDVAuJ3tN
YCV4fIMQdSNR53nMaV8VN51/hqO3hJ4HRIz+3qeDlfMxuHe9dEjtxZG8qTwT98T8
HSJVPtK2Wjvif2nD49hza4dp0TTE7NM+XoS+7lEac1Yb2Ac7lYAN88vwj7vFjHNn
20Ua0PMDFruHmQvga/owZPJzzbzxa1sog3PbYLUoxNmWA+QHlZsSwMrNXQENEhMf
n0vxIvXERaIcHuhejgXkV/XL9UyGbBOzigM7GGbYOCQMtpY8/dVOSjhDHNsX5wsv
qAwo2mWMN/bzGvRZlUuV/RS+ZUfYjRkDXXHwYzZtvaoC++2595nIGfN6oJAoy7eM
QTx01IZwes0FRkxJlEorQrsoj1nqJPR9SM6hw+X76sCyg8CNMxQ1EagnCqR7VVWN
Lysyomk2sidAP9Q1OXA2LAL4xsOJj693GVckKjQ7oOG3rlY1Kz29ZWGMJhvu1Rgi
KWxapNvSb8X+LFEoITr7Lsjgf/doxrbETILgsYeBAzooGQW9nfUv+Gzg75hQK4Pn
8P4qveCwlRNVM1F3ZwhkggMD57gCGOp7k9rmng9fU4djTGTXWq5voCNWdMw+Hh27
Tq63H2e7hwn3kgDL53R1IyHVJ0uUhPW8JsgjjAR3QWgrg+0UhbSaxkcLQKowhnqq
D4Pk5EFh0o69y+3jtreCyRJQ+bbeXhcAq7ocwnIf2JXVvxyEmgGDx0kyuLmLhigj
y5BkXsfdV28UWOfYax9sKgVuIhcr0NYGCVT0cnr8EX+QWLAyJyosYsPQd7S8ZL7Q
fMi6sOm9AyhjjnaEJUqZaR5m0dws+KjSFILgbZsGs2QDsN1lhS6vPOYyEMRcXWwE
VRtU4IFiySg4UjdrTYRnFJ/ANCxqZ6Z449xRVjrOvEjhtsGv6Wm2FOXu9ACzFImq
cmBOn/hNNx33wIg0NHFXsL7XRuE5u7t/lIqpDX6Z7v0oZf3C/O9dwDhmLg1txX6f
ohUmxcYpl5vetGM5e1rTorcaP2rc5h1TNSRKMa7DjBi8LFZyedBHbxL6tIS6BoyP
AOK2MgSJjkAR5Rdsmb/Rm9voXnprycF4n2RR6BGie/EFiwPErr4CefgB/G3KgGY2
Rff67l4dWB+25Y7ECqezWWRJJpD8creddsRvdsBiOwfyc7I/+wM4gC3ObrvfDkwp
volKLbQJVQuEcouxJOa+1M3DH1EU2l6eQWw9OD3/hmZKL+KqFv3u4yUbHjJPxpGA
+8dg1koDicnScBdMiCgNdkIoE+BLwrtmwkGGwepCJKiWjAJlERQMLu/O6NQBcf6i
ygrwrygu6URnK1Ua6YcDugw+zXm4AKV4PmCjKoDD0nl9UhO77mWde9o9BpHB7wEe
ChIpV6iat4F+IIhEZ1mLoz6BO++U3SQsFp85X+sS5bqHUfmWvrkU2iMhHls2p6EP
3vmv1L6ynxq5Ypuw7BVCpjQ60a0DetEsVTpwuo/F9mToCHkWPT8hHslrlN7LJbR8
u1cJZPVC+eDZgXdzvguaNtYWFUcCIYXgi4svwdOirBpp68QiE9L71gnQJ9R/h3lc
4FlsFvdNo+utTm5EMsxMGdiqBn7IHad+JHiCkgmJ8b5V/ENmipuFN5D3jl7cUvgr
AuyX0KsZ1sWeSHtWHkyqowRo+5lr0SPT0U7ZSlafC4S2GVHsQyiwWWtKxtaRkKUQ
IKzE3rpMhCRJlP2Ghi6TtCIxT/hdVy5Y9wrQpo5M3+yy4Y2A7Vzf2qs2+m/pdoAI
3m7fE8xQjhwB/umLmfe5izq3ACe3uGv5mxCAJbXhb5MwZrYc6Ege14xoz3+iUr0N
I+VFvyzpjXPOy5v6v8fNUNx2SiXIuZw7LFgLIyHu6wldEqV7gBawkJleoGko9tAi
bmjeHgiM0tWLqbJUvOr41Z9HglPvxKdL/zK295LHSJ5zINaVSWzPJPlwJIZkQnLI
g4DAj1yMRr68e1OnzZJx/As0YHgrqcGTAiBVG8BOFFtCl9P1i1WZp376lGh4K94h
qoF3TZzZyNmspFhNEiwpmAyF6LxH6AK+sVCAKwnZw6o2YlsH5M+YBITpge9PWepx
ehjbfX0A+soeEUuTH/ZXeW19Fnb5k3YQsor5NQAJ/a646iO1l4uZFkuMsnKpQdJk
WLul57vKx8lzvCum1wBtzyRZ5PGBPjrWaOg+mcLw1OVyoTjn4PKyJOV4Ac0n5Mg5
93ePsjgKMLryXNP/hKe1z8MKCDtODfpMhHqXqgFPZu6fdO586XfG3TGxk86rOGhr
BZpo2sMHJzRVvDS8gYaFIVMBtNX/D783ES/Zkp1LduLEFLASrRZizu0r7xNJRZOl
amQOywUwPAoJ0Zn/87m6nwEokJXopnHFoVlRcjNEU749+oe2qsiHXXN4dcZtrtWZ
vatcxMNj4hVyqmpYlBnls+XiSXA/iNTsYF9UB6/kL+MwxlKyos9xB6qHMmS7GdKd
/Mmt+xWZldWws/Uai60MMuCGz8Hfppz9zYcbhBJa9sRwaSn06NnZ/rIWbsCDOnzO
sML6qRbItvfcCzYGwrc0DuruE4NfjKRvuOxORzqbQDuhESxBjzS9iNvlwGyzk0f1
wYyK49dEJdb67IDnouMSkklZKXNsKhxZaHanSguMrCK+prWFRilMjZD7uAlVWoln
LTQQFwlC0u3IChMqfrsT8Z0tNCnPhWhbzfy0jBBVAskTFc4i867XiEt2gGvuyQUS
/JYSOIjADJ0wIWGwfP6XZBNCNNfW3EThBiQJHfanVa8oc43wDc9sSp/Nw3aB2gNj
aDhFLh3BKB8zwlN+VhL7n0K2nT0jJ1vj2L23xT6NbLuxXGhpq2/11h+XJWkuV3Vn
sF6ovirVHW7OEfc5r/wVv0QaOMUCJE3m515Ay6lOtGHmYwLO71/E6fOJtHajdIcd
2Vz+YV+mHYlvkInJmJ4IeBBD30aDSi1t2cbs4XCry6XZMdDOq0UqUGTkg/rCj8g9
SnZ4BzBpSDaU0pboBsazB8Urn7mE46S/xpNWsiFDsLZTYzy/qKi4c+9mBLXXKIM0
NzWUWeqZhsQEe1NFMQu9FBOC4H6d6D4+X+dBZzeHUlDjzmUfwLlviQhhymh7SbeW
5okKdyMe9qXT7+ZS4kdSnPl2de7xLVJdbszVvsLfIny1LAx4nZfgTNivV23DTUl4
irmlr0Y3TWEaVXH6iZ69mmiF7xl9dUpYh1MeNm0fc8BG5wbUXtmTQZIy3nj1dEMK
+PZ5ypb38bTY9SLRaOi2aTuhucI9Y+0P/tKL0qrHM4eeobVuVHZwkQFXuYc2/nEC
g7flwtL/rNjIEpQcISo6jwEWNn6ezcDXhkrH2WwGSfwoTdAxh5JawC3pf5W9QIO/
7EebP8f3CbcHbEpVw/VySuZ4EerncEjllVY01Pb7GeB/oBKMdQ+WaQON86bwWTg5
Oy/CJsZBzwM68c95KNVhIEaa/4X8+tzN2jQRrdZgPv/qvp2FyYh2HxYodlP4tfqq
EEJqy8odz+rkEdKa2Q6oElYFW/MPGXqQjngVGDZhC1RoakiEi/0ITG86/XHauT45
IOVFecWuJ5dTn4JeH56JLkdgKYKdudfFu1YVWXoeeDb2n0iNJOkxOA6W6zXBFn9c
LivhyexGaN8RWBYBcc8cwnmlz0mSVR31pw6MmDhyMsRnw7hsdHgen6wMcib0tXQW
eNfYyREbL1dPtafva9reFTyO0MDdk1BGLEPeH5EqJbTaTf1kPETDZxWoEbEzCdr0
inNRMunVBvHLNJHTY01dtjDHz7+1H/QfmgnASNtk0bp6RbMAONl1uaecrRHPtpR8
UZvPH5Dvj2TVmf6dGFPf+9aK6NvndE/hIa1palDoRaa8hhw76mWiiDK9xwbmML7i
HKq1xBM72uk5AUaObRIMi8O6C+wFabj8QBl9at6qLWmnXu4T7evI7TzzYxuvLMDp
vFo+N4Fupg6YCA//a2VsW3ZsvcCxtOoIa81DKa/tbyoQGLWpX+QbITqPCYUWqkrL
geBpaQNy7G+aAZg2wlM6PVNxlIGpDZG0FCjnhz9hckU3wsSeL1uvPTnOj0eozOrq
c6PzWe03vlY3wHQAqenk8jFMNWCw+HEfUOdNiICg2nl/l7etoEIedTXWmZ6bKG6G
aY64LHcRzw86MYRYyFEt7WNJr1dF0U5GyiRjnY90M1BizVqcnCl0lv93PpTjdjUK
8XNyH/3/xTr5EQwOLA3v6TCHAg75EusIo2pB2ImydzpA7AoI9VmHIsxeMipEqdZl
yq//DKAkKocK32BCt1SYWeqVvsHlZixUdwr1rB4XgwlV+I9nKx0b31rtM3pgdTsC
TmWThdQgfvpYFBKytYysThWHvmjxLAYch5PcRsbdwOCZ8gnSnHq84PNqAPRHThid
NVOvZeEqriL8t9z99XaMD9I1COagE1uhSSl6pM4RvgM72IHihneW1/wXerUTZm65
cH3lLxRVf3Ealm5Nt4stckx+vxBTemL/qaIlfpRGmxbVSITBAQNefDBPb33Qkgq9
TC/O+AQg02t0iQ8/tGhopRJGXtRaMqOmmp1O7KYIGuIL8t4+pgcErJ4jgBht+exN
McJ69BGyc8to0bKwV1VxI9j2/v+8oTs73dShcc2H0RF2lJS4yWN/+e0ZBnIevhxI
w4GuGzy9IbDor6I2jbEn4ul85UA8iCygDVX0Jh1fhGU2tFE8nN0Acgw+nxngyp+9
R299e4VEYtu9v9amfBSB3Pm9wT/lFNuA0R/VYoqNMxw0MPu2kK2tmrJ7dC5AdwXm
1l0gju62HoO4PG1DRjMZFD3DL5bIRgrvxZ/TYvHrvl9Enu2FU/GjNGHjBQ0S7qUP
6H1bIdg+XdWqJzhxoeUldW94KLBoUxIdjXxY9AhF99flcQLMxmi+Q3ODu6lNEi2Y
CtDaFJfl5KwWKS2nknf5NRt6Uw0RcpNMdmZalQ0NyOaWpJYkl/mWPLDi46jS0/EU
F6sI0Gp5K3rHLXy+qHT8CQb3Wf5naQ340kRV9bvk8/+ROkYV3ccpdqOkleeJzZbW
b6hYkY3LguE+9Nl97PdfPyoucCGY6Q8b2n9PflpDUjLk4QBhTfBS0vxCHgjnfoGY
Wa6WK9y/+RW5DQk/IeNZDmKTCXhDbrh/G6piaTzwrdWWElQB9ZagMWyctYdc8bWT
fyshdAYZKwr8J40G8y/tIACVF6C+/uKN0veb6EH8uOgITNokelqOhsYXfsVAsj06
QCIOjN7YAGUWVL3DQ8xcIaVWqebjpzhBRGHGzXNgcasilQ4LJAqsBIrfHGLEZ7RQ
3EXBp3Y9FPLQrdzY7tQo7xVim4L8Xzzeo8X8y2EYfInnoQeQ2M+EmFPHXWzHCv/Y
2Eisqu72wDXIIR7m+RHxWqu7w5pot7fR3juLjGgMYzEeuf1XJ4BH+3BdnhSjeskg
st5cMow9ObHL2Qv8CoMlqF51gjYR6WT/wurN4Oofr/gvTIpxWXQp2Lv0wXf1yDZz
uCUond5frs3P9nE08UOvu46yTadDd8l+6rDu95bERfhF5LtTLxjox9TiZDT//QRa
PxIk52G6HuShXSK3zM+aGO2wB3bNNqojwQjNMUP+f28AvRdDiCU1oLl/dFG92hmd
Ua2oK902Li2lia8Ftd5HaMG0IM0bm020nbA9AVQ4jZcmMnhQjD3mrnvRXCZp3EtD
In+Tohx/CkqaOUOS1MV5GYCwBFfWMkD4j+4/yXTY1fAraHwT0k+oANllYL3ak/kd
eL6ne39AffiSf5xmMwtd3rkpxYEK+G07apjqgj/DGVOBnuZYE5zN/vXuLgGkylS+
5Kdfh9SZKonuZWoLLYUnhxDBLYu4FUL88RVhDkGxVYCpXCmzH0L2XX8QjGcSs1MQ
riWFT8U14OjMBKLbujHG8CO/NZKvSqALHljN1wdmYiHuZTjRr/aSkIuQr8pSy3Fo
qNARSMbvBiV7nc7RGVaZWjsqEPG9IrpMX0leGbiqzcr8zorXKY7QAna78stL91Ki
3jUtT5HrAJ1iH8RgRN3wabYWiTdftI6r+taD6PPkQgTLRgxDxS/UccsFjR7B6dJ5
tN3oKkwjlUF1nPCgbh+ajD7oOjA+EfVompgunQXcZtNztTAxpwCJfbegiBNqoR66
a4w207uizaa3Xp9lLXKuVsoOf9SybR+YH8Gbn8EbvF/Lr0BLwP6TxHSn7QZTKvyu
Eo4eTipC0YDFLPyIEWNC154kL/smeZNqr9LY11Q4FY5NtDVktNeSLkmxRvz7Whz3
CggTlCW0KMvHtfrPZuoM67ONA+tUOFxMl2aNkLe67OdbMAM1AeIYlHMlGAONQvkW
yQiAwh5JyM5SrWHvU+E1gwU5VJCVFXTgiV5dWy+W+Lrv5U+wINBZRlFXq8Mg53A4
OLRPgkROz/J0DkdhhMVMgv+rBCHQVyLsTM7fCWQbcLb361GdYhD4lyQ/tFb9Lqh/
LlZR5PV3YLHrx9627sWcBnJpZ7Rcn+/hGpJEG6tvldeuJ9TXZhfcH6aR2S6KBt2f
gZLStOo9WCKOI9iDg4+kDF54tZPIPD0POLb5zxIc9VKUd295rkPHxdfMDsxFSjB7
tX1Je+MHRklO7SJFI+o8zxCV1TehCR0JnQn7pStpUzwhQ0A0Q94f6iY0rKIiUqBR
CtvmZdy2b1F3ZLHQUYxks06c3xym0N4jZD22otgFGQr/6xLvjBCxcNchqv8Iirfs
q4y26aDNBCsMRP0aCIQVx+vsg1+NxkP0E0W7/6WDTJLVFjIw74vFbD9X5W9S1luu
XxMuzyNzUl8Vw9Qcg2pESrkuVgV1ppbmWD2h7WQTGcjLHevGWoGRBLkCIrqUz++f
6/XZiCyANzXFjlso/60auByPX0OoTlkgJ8gsVeCIFGfcn757QH5cNHOTSe0ydyiA
SoST3J8jNBOxK+gvN+QSMI4CwmHpygk0sZfN4zIc435oDW0QoEVNQvkkhMgP2u1j
AZgbRFubX/EO4SqSc4i6TMqTiL2pjRL3Sp4D0VdLHyxDshfBl8DM9ocm6vXXtTMo
wlvSp/KDjlchA477JqqFoAOam+RT3yolo8F0rS90ac3FZVqNU/AgeMgNuUUPXCYh
CeIm2S3lH9pbntxx7TRxEFzxM7EZ+XdCaqKr7urD66ds/QNXFcOgj4Hhh5ssU1nt
74gjQOSfE6TIuyFfIkdSaLKlYKuZvjfrf1gXboNTVTiPM5O1HXnG/OHUBiFvx3dS
+274xndWkG7pcsZg+w6KX0pphfFw8GUvqZpN5npcVxyiDt0lM/4EYo00Bf46frW4
MDDuqc0ik+NLaVmzZ8WlmzEaudSiRx/jSq4RxyewXTgjBtrfWvyD+wnra026CpDJ
RB6VBLywAFRHhtw66tzoi1PufeqzYJCirj83cS6Z9sDjhb2CqAjL1z7yF9ltZIvz
9D9/gOpA67eJjvDS9C4Vlab3HGLsG4a+co+NKvTFoacKeFYVTrlhBna4J5tsS56A
ERfvL0X1jN5ZqLwPtPdEdaHnx5kfUM9X/y5AtTjMtCBTG4Y1iaAEljQJUazp33fu
Uxrp7D4E2m32TEL+cItXcPb+k9anJaTGrq8lmXC9bVIsH03OLy5sLZziYh8QZCA8
PXDX8ZiSEigEbCdFLc7/YDdaHySFCgN6B3tGVoC0O9tL6NZcoEFwDo83Ew4yb6jr
VShexpt6NIK1q47ZS9OSjVN331inQtTAJRSXFBiM7gM7diE485i8QqUDEN5Ivdp/
XShZFqFaeUAq7rvhgS04Zm2v8CcxknMnmzaFDQBBlszKd33s7kOEf1skoNQeqevc
GRsBN6WGsbnbqOsmV4CkmzTGe9hWCSkOmLHu5ARcOBD7X5ACUbGcQ3qf+OZ2ScZX
v7kgKE/ZHFzswTTy97ufQvihTfa5GbLiqyLGwJHH4kosagHh26Fiw+8CLAN6uG4j
likiyZb/AQwPr9d4oRLPQpl1Nb9RJFESg7mg+Iq2Ob7tE45Hotr+wUKt0LKK3YUt
v13Hp9xC8Fpymzeiqvs2i50Kt0e99GYEYZJ6Bs8ELIbnprBY2bbMhVHpx9yY11DI
nQqdwnXCWvcm35cWHdKb1NXdo2734ME3BryZi6jSyNdkpNpTSt97x3cE8lB7Ks4a
iVNzbbuvo4ZBoX5lQqiM7G4MjRlAG1ugWosz96/cTFRNlg308gFTgdAQhN5/DJUc
0oIV2hwUCsnOC9ezdA5J45pFgNKMYpQGDkNP6tMRuX7VoZVC6D7LH7yEj6ozKl/M
c0Sn76bYx+5Hh7AbGXCr9ECXxGT6V2jAJztHhaT1vaUdm6DDIk9XqtDBkb6e4pKK
UaL8Lu+l3wqqpqU0eapGQtKpA3BVIVUBIwlWPj/Bl9iOlJlztQyGP/QtDAJJc3Wh
cRtPd7ti9cvH7dYVDdRq/GjpF01CqUo5SyshsvOut0kIPrn2OB0xHTiQ1GIoz9ej
v4bOI/lLYWasfOoxxC+QrSmea2YsCUB74iluMhWdOofQIfU0tG/BrfUrdMjZP0lj
9gINZ7eiOOpmI/821TPOkx9t+KZybpf+C0j2qMXUl7IKQagp+iFY3aYQTHLr6QnI
rzJQIsq7vGwSsKa39U0EgtMmrqiQeg5Yh7VYXVW29hO7SpWrCxFCrW9OdtGwaXWb
BXSY0qM2neNhpxU9GORbtVQXj3aBGmS/YCOqlimT1d4CKVDbfKbWKj3LTl0RYwBb
+FGPIiWJuPcSulWXOeh7E4/OE5APkK/6PzTM18XwVY9Ov1SlqktR1t4dMH7CZzGQ
5X7bN6L3+4cYIeJjQ1T+WteuUDETJJJmtcbVOD0G6BySOxTucrEEgrlPgTqWYC25
VaY1/b9DeHUYHOG639HtGdD3+L4ORPIiwpxn/QGzBGJxyrPB85hxMiS0uuzKHOMM
4Vb8CUga5RofUOiWfb8kkBwsXoG6F1latRAxTxubEcHg5ZR/CECT0WDEYndrcsqt
ktbfLOlAZ9T7/GF8CH16rrzE0s1l0iu/n7j0Ag+dbb5R2xYqBMHDnq2GP6zIgzyC
e817Ljv00fqFBkN1LW8f93ewcc/s4faIS0+TWqBE+URHeajDLqxI0xaAjnMiWPzz
DP4DamFFyzA1qrYainjlTXlTq0JIYQrcm4awMq3FgEoKG3OeWF1CpgvD/YsijL2p
1ZTKnk8AKsvWzAixjd4zqln5RH7biHduTIVdiv6BmAx6IXQTT54gECSGyBiezLyt
NeKEBHTljD8pKI1o3oHGiqmhSbQXoQjL/7hzHrrjQGwaovQ3aa3KTbexIFcbhTod
Pb2Be0VS1k8c2K7Sg8XgBz1xG/MuLRTllt618dor1k6WD29yxIZMpRtGLNlVT+Yd
rUB4wN2vcLeKDH+UZhDZpjkLHby1PbmeF2T+sdTZ+JXyOOIW+HKu0jgugMML5cj1
X/6QS/rN2Y3PYqid/kukyzeX1xm2C5ZZdErArhYuI8/s5DU3PaoSu6SKTHbKjwRA
dFQ8yt4D8bCfdoj9V0PPTm7xJNhZxA3IU2QhyoehjPhtimZvUs+SpqHZ/Oq5yhC2
HzCyMHJcxHfjii4m41/yQ93nuc5BH6CEUUM6wVpl8r4HhXZyvKhjR+dZUpX7CIQ8
gdp/CZ6QDRMxoruJcI1JjQnTMFv6l8DS0M7AJpNTwNVklcsX5AOtJkxoxdh2rqp2
a2qvF4jmyUBSMaehqpBYE4YA+i/CI7U0U0tHeyv6G+nSvq/5XaicEnA7rQYiS0A8
2trbcCme75prYxRr6Qvdx3+flAzKLS0vhqmIarv7YeMXYkOQYWKxBbGaU5crHScu
N8TNxr+1uXDYeI+3nqk1RADIiO04mBcSt0kUQjhGT6i/y7PVB2t4uyA+8B/xUNu8
D+e9WnVSkijlSATgq0nmMd6rGP8MESKiV4oJV8b44PSWbE6FUanUYwBFyomdhxKD
G+QeCfO+d0WzbDO1yCAgVdE4bqGtHmQFrs170fP0x1XCdqT4BcqBh2jv5wEkFE6r
gGTfImcmu4MjCeGWAJOgoqUEnm7rmfccoFurK5GZIFzMR10ZI9jocIzT9UoH3pSZ
hdJiJu6kP4uq9f8D2kzLYk1xElOhYaLdpy0zAbZnkWUqNgnp6HsQkfWXPe68ptbC
2OEjXysdhFWd6v/+87RlU/Fuub5Ri07Lg9bZPHb9oo/PRRu9US1uiY1MWg/LueRF
TYLNnnPVLZvxUIMv4OUUsDiwf/DPKrlasArcYk7Z91iQEPgUxPIo0Sl/J4S32UWk
R6AJ3b5sPDb/Vzzg76iZWG1SnHynwbnF8WceVDZVq0hUzK+KQ+A6onOrJGEBQtR3
3qgV2b83N5/5EAFGcOWP2SthjoPIgq19do43KMKInXblw6JuExBd7KkOihB75UwW
RIeOXZGzvjafg1VTTPeUyN7w0FrWqB+02vc3DrfmwI8TokRPGQmEPwEU4Hr3deRC
jhBPyuDYHk7Kw5xJycZnXpiQjOpPbl0w0wrqqEpkJOCK26m+diyBq068H+TX0ZA+
/FwAi5j60Sz95g8BmvK2+pgS3L9VmGOAbGNgIZScyHP3n7AKIqvp0axcSVscg6ny
wOeoJa1LRY3sWDzkk+QKhMVhFiZoJbIl+GiOLQrMf+3zzEOGxlwTOXn4GviWSSvY
nscuQLBHAV75TAPcpLe64mM6Xj3gKeKiNK58IvqhsaX7G7WvT5hxypnKlcGn06V1
zmXbtQjFog04cJrF2HodQHicvvUYpgCKZ/x5t0iNq9wlfT4rT2C+L5bwZcjbwSK1
as+Is14qWLaIJ/XBKy+JiwU6gcUJPS3oHFeW58ndg3QRSGh0cwnJz9gCcv4e1tIT
rX2+3hVqzIA8TU5N1Ez783xWyvtCx6O5qZWpxmijC6o6R1oRcUn1Np5Uq7uDHdUO
JcfZgD83feZqFqhWZ4luzlHXlSs8KF8wjrnfAQn/NKBU4jKUqdxHmpxPiiHoXXtd
s9LgHxierC/3UmHC2pJRzbITGVEUgLCC+VdOw9GXT6bmZtBYXlL9wnwTXl8fXRIY
Zwe8fxlu4ExaiMPd6Z93WKaHCGXLQDul2m46ztfInMo9ZO4tMQgRChf2bKUapdwB
Kve8Kv+Ix2VxAZv5jAJwJmwLWSpe1tU3RBtgaHhpWiNf1oWooA22q2Bu6DbFevDQ
OSo7UBqQbsDuKGPQyXXWIfM60TT3ggRYFE9tvDX/QWboyRQ9BrV93gAQboJwipkn
R69rdLxcfpYASi+bdrNm7byvivsIizRl72dHL8e0cFFfu/ZCQy4Zid7+GeTUyvae
ndv323S7C+37+PzENPxtiFcAcOQdr3nuQwpFLznYaqSVQYn+nE8u/wFV2exJaQSd
cblUd0rdspbdsOVbgCkBMiFwrKp7Xrhc9mjAwLTkq+gRIpLbtGe0tUHw8JWehunr
5l1AseCnQtsjT3CaE2YTjaARUqvnKzg18E2esfUCeUGVx03Oilqx/mKr8KZPtRJL
OhkCNiIa9OsMOFLa059pPNJaV8HPBj2PfTmSMWthH3qcL9hPnIklFU1rg7IxxonJ
DfL7xDgVNty1tcDbs2x3BxWRLFriW5XNa5iUNMYHpndtsxViQWLY/bTGxp6blpQy
HlNrU0v+we66ToRsNDLAOcdqE3E7vn9gpJxjBlkck+lzz6piTlPg6o0wCJbE/hSq
Cc6Snlu3Arb+10/MzTBuYtxccpbRI9z/C33zxbN3H8IbT1XOLTfDmBgMfEKm17zg
SWavLlPB3IbtMFDi8HXpN0q3RacrJkqJxfGXKm9KSUyqGgVgIA2MYi5tqU4X4fBX
bcWAINHeYazhcySZqXk1kiiBL4wvG5vgGyW9BY+Yj2v9R1AR2PJk7v+/JhzK2eEF
DyyDeFuMGYq1MGYKqCdmOCRD2IQ2EwKkU5fSJqWcL+73Gzj0IECoDATHOPz/m9ia
2EuV+/KhGGyAFXnzw3lXU+6K7HGsT36mqTlMgtuyS6PsNoaG6O37r2Udkcph6P70
EB5La2wlMifApJVejSw9WyLW8IgG2ISCJQMziI0m3qxTPH2vzzssU/Xo3OwkK7rf
1X6gFnlMeNj42aoILYldDxoRs1sdjKN5exL89cmrYrvLsCTkgC5dX46Vo9LVuDOV
JpCYJNmrWz4gWN1sks52BRAVA1OgZRfCE28JzvBzNtPMdZfjf9itC+IrvBWE54YX
/P9TTZpBnYEZjU5Wi4j5LlQDpHY8yMh2ldqAkEsTxlkI5Zw1mi3/eX753lpLrEf6
LiHfVJd5JOt6a6HxcFzE9/sIezQL72XTXgJZJ7N/zh/Kidix0oyUXHcqnM1Z4odV
Rbl5/ABxHHnUDIupYFpAFeWBsr6rooL3I244ZvQaR0n2ljR1TU8Y96q9zn13n+hS
1G+E/n0Ik89O2mNIBv6/VB1Q2VxvlxapGBjeVjsCfrAcalcnk58Cs7WVKkm3NYSb
iALu99lUCauu2woBH9eOGYPINRzM83BgDdPTi6//DfpfwolwEct+uEMfNcnTsLl5
NRV1RKOrEHyFqU0PcA+zu+IrkKVg+W8McCJGPjDSVZsE46w6VLp0keori8xq0kHm
j2DQ+F1HYVbT7T6RQAkPCN5NYuPNShiqMOANaMv9zDIlTMMxHusfRJCskpB1wGyj
gz96b5eFyoZ/xY7zt84cQWZqksARFgZp8RgYvZMlQjnKXs7Pdff4+JW9tQtiC327
ifin/wKGoy+D8VHpLBXCkqNf/FqPSO1zzloq7Mse7Z1ybfRIhhleb1unjj1PIhfN
wYNekMWF3soQe/DoV7JqOQmq01riGjNJNLNWK1jFd82g4s5lvWeBwNn7Mn3AR4Dj
GwXjnvBrpyR5f1IybMkHBz+/VXPktRmKtP38BsXnlRTL+eQhDtzrUuXPnRthylwb
RM2xCyN7VjdNJZasMT6zlrzuLAw0TIoS0C9DIqxuEMHW5jZc7Qac0YnfiPxRdgLg
p26Bkw++L05IS5aVTVq1a++4AbqVLxuQN2XT3577m+Q5+kJc0bBaTiaZ1bmzZGcp
vT6/azy+9BKA4b5mkti5EJpjbnNIOsbX7f5wTvX2MO+Jc0qxCytGAB0boGQh5JgU
YJXw4xBgm/ViRWLH7Dh11MAiZBoxZTMNBZcEdYc6BkfE5XXyG7NpxF0dXSDKemoB
UIEgvPx2e2zpVCyq9R8YbC+RNZtPlu1ADjBaFi28IfTnE9TXwP6cHpXnw/NC+1Wt
uO222o1wZ6l1otrRb45OV8CeBrWwqqGVHJCkY6aTZ4IX61/H9uYuPt07NV9N8ZXG
8qVrCkGbkLSMkP+23ksDZACDPgP54Wf7k98OtjRUAuDSc1J7GLJQsjw7GIklHUBW
2RXboHxdu4UI85SjUBDzBI+48n4RBy5mQoO9+90WZFEcmXGc1gReOv/3R0iK/oiG
qQ8sX5rCzGV94OxDddtZSMjkgvtJRkL36a3879J7FgK5ro7p0Jlzyjm2Z6wlkv+N
nLmog8aU3W9GSDQi5qG2ZaWNW00nqS6C6DIQIoKfUU5stSzqxrirpPs+mbryZhkf
FLktSvm00IVrMANynL9W7y2HpgCyHW+XsEIj1QCEIRSN59i7jByQLpgnwhgWhqdw
yDrX/KmkmJ7qg26lk4COtegZSw4tk3z/qTpvRr2RaTfKqc6th/ef5Xfa7rQUk6i5
Uii9Pr1D6GaOQk9V2eFQtloQx5/gFtrcqtEzmztor6xCg6ol0XPZYh+XooQAoO4h
rGz99iNjFHWvp09hgeleusDiz8kk02Eq76Q5pNKvOnckAkvBufafFWLAIT/GN6Dl
Y1BUO2PzVaiTQXY/Til1OJacM9dSVAGN0WUgVtsLD9DYJr99FTcReOxdzzEWupOe
uy8BdmXeTH83eaiwSKsGdAe2/LosQEPGGzuOimcyRa1E3kwj6aKwz+vEWg3uSLqB
XqgV/MPo3JFNIePXP7RaEecYSoXlKEevkooC5NJIbwIf+zSWc2blMKZMx7NiSKiJ
iKv2YJWZ2ztC9YHYBgLSk3bG3odlypVF7PfTZsm2AWzmHohBy2qTTzNws8SFb0DJ
BDHJTUQaZdWvNBF2FEWf9rOC9MMEvUwY0swiVlYy0wqfbRbHzJXIO32+Xw24uo4/
qC8AgOrxEL5iU/bPi1iqBrn5Cjm034S/0s0ky7FSJeQ6uWoyOjAVk0XkOMipwVq7
v/E7J5uaA9CO0zr2VOI9Rr1bMwSNRwx+MfPiaXmwof27dO7y2bSmFLX0zXkuZR6z
+h9H6OPNtAM+XTTs6vWbTtT6BnnXBLXLSk1k5lBIVz58slQrVSQP7vWpP49OoURu
w5dywkqdfCuZmXT+cs7RPpMn/nw4T2viyulpS3kumMQkDPtuLL0UJIvG8lEg+bhe
45SK73pcqakvwLJnVOVC8upne4Vi23CSrxIhheWulITWldACEn+GMNzz50yXzoOD
wQLaFMKeLYjQIJNZLoN/INKJa27WeMfQijB+A4aG4cpKmtpAUHDM9/2XhrcMdn4W
VXMwvd3OkGscKnPz5d7AlwlJ0Z5OeU6nRR8bC/4VvyLdidwRMWbNhB+bO2KCCoA+
ad/OOTt6dstqUINpfnOQzjgczIak28HDTQv+EZOebxAT4QoE3d/ojbpPIwtstbxI
LpA/V1Zcb12JqpPWZygXBYbW43QqS1lFSSvkHuwwxTNUgvOgY9Eun/Uvack1+poQ
09czv1NVRxkjM6mx12BVo/2dehH7gfv1kfVOZaeQsM396B5407prBa1Ve9i8nQa0
X65auSM8uQZ/SBJ04zjSsIveiP396ndbHPnV8vXupLBLJTbCnJQVugzolpJy7/jH
Z23uZwnpcLk8ewh8g0YuD5yqhOSMM3TaO58czAO4/k6zoeTduEEGOmahHUG/Fbom
pNM3gdyFfbNKOIzXQ1sU2f7UHRoqq2e1BrFm9EDPjfmZXtOXysarzSY/d9a5MURG
e2GNvBtOA1cff4+JtsfBTgAwDGEXhIaGHQIF4Dri7iiEa+Mem2814dLLDUdrPu2n
fcZemO1IBITcVP05LhC9sdurhfhkpkQu6fzuMgIe+7TDAbho7s0UABXyarX58dNz
iPzr7jle9qufrtDrdUs/TDKEkihHprMp+19SPz+HMZOrwHbZQTB35KsUww0MoNiS
y20eGjWTA/Bn8Z7+VzVS1X8FwPuDIYptLn4s7fELUiZNOctONiJ2cd+YmNmRjSTh
JlKbMUxwj1TiUhcaVt0AJsBH38vbc1T97IXBUbgnMyHXfv8GxDKgRjCohV07NCUy
3Sj5lVkwiyFvQ9T5/kiQlY5R6lUDElv6YVMntupHcwkRGEsceqoudNX+QrBlOQcJ
MYqDoQR9ROgg2I8AMEHF49jbZmSL85RXyvl+HDhcq13kRJY3t+U6Lo7GbARfabzz
BkNvEOa01iaaBHANltQrcWEposZFY8SW2jwxQNopCdozIQHdIyZehtNqCd9qJo9R
VTQXeJTsa7jGPRehowwYxXyrNyOIiRO1b2KOCC3KFxoYITNkRC5GCKyykh3pyheO
Vsr+Av+0k8iO0wLkwPD4ApOvMXQVlnPMRVSk4m16r9OWZ17FaVTQlecMhiOpvqo+
E4XqwAA49Qhur2CdKzrVYTIraT4fHgbpHYIfY0cQ/VzzQ7aq8ztdLixMzvufozIC
Frdoi60XFk1twI6HW+4tztBv0FY+CFfdRoh3b+edl1YCwvG7P3eOz7tExOcEehbc
UR1KWHmzhFxOKPB097/HgHm1+bHRnscikH9vKkF2JC9pWijHCHTAwtC7XSvzAiAa
Tae0D7wxDqq3B5xFbnMxymMtFRE1kYM8gDA3rCYj957SjsmUK9ZdG8yT0pkE5qgD
BnLWfdzK5BP115hX+UD5lsMi+ZLrNATkZHx7M36Xng3VMUM47UpoAzqFh40h72xe
OipNHr6XPb7RxlZafKsXdgqtYVmUff5yv8xlnWapLlOGM6jSbCP1OFXk3+SCF7SL
ty08JvDN46sJYOwIu6bktS4LIf93/kojAFR9l0EOFs7nWFci3cPqNK5Zuy2rX0kX
v3SaVF1a3jgbCgYlyb5QpF3d9tt4BtIMn49n8goA2opcB0cNihs4kdukDI5ewrST
BAFSFw9tEvkpWa6z0K7Wosxk5F4hcXoy7mlm8/uz56/xPJ9262pW728NkVy0XhBY
lfrXJAHmpEdCwzUXn7zy0lkkFf9JUHBndP497aaPu6lF6xRSD4sH1mz9TBKpaDpX
A0J4A++b4M9TIMNXzLXHCBbd2ypSGc405AD1GEZPTo+XnzF3EhhD8y8BT53yB1jR
/V9VRNedsrI6kyCJTtRrK0Z+LoxyrT/DuSRYXKa7N60e7G2sTriwMoHfFHYeyYNT
cRTaazpm49aN4GM7Va67ScV/Vh3J3h4Dg5K+kIypRD4er21eQDfeqWC/gevW3goS
RD4b2nsBYQ8m+efFT9k5Uv5EGBiQ283b2GCfzM84E7U1cuCfFI3Atdlz4jWyLT5L
C5NZVPXHQ+hV83wEaBGzR+mk0mJAbpAXkmx6ZYqwd2MmRkLVCfZVZFjDlPAvL9o5
Qvc4x72v8xNv5cQMjTf4GPtwDvYq7HmIM1GTp9YfMqzYyefsW8gh0Mo46ngGbAD1
8ZtyMi2UFoYgDkIzyj1sHKHyCJOI3IE9Cu5I6y1m2pLtqSTYv3hlnJZlebFTxt6t
1FwLA7FxKLolwMLIPUeswPely2+oCuJoR0KkU4ZI/kQpChHrNICdl7uWOZDYTUsV
s9Io+zbOXnLRtJ7QQvcRSTDb9L0ZFUB3+WsxIzQQ8nqVgt3FFQR1pc+MA/WHJAKl
Q8UGMggJm30ixspKfWTIGOlyti7WgU7HQXIpxvlus65kgrbYl/jxGxr3vQJk10Wi
pX0Y4HIYK3LHUCWQqPDC+8Q3HrXxzfOv/caOlByF5Xx2XGxusnXEGbaOf1GaXwoA
ZQ5NXp01Uy1cGJXT4gEH8X0jvCA+F2txIhehB//X2CR0LYnwLU12B5UdERT7tnUb
zESEgD9RyW1L3XB2epcInc4gyXDia2MDQKHLDjMxGWRkHLof/rM9UwLlihCKsCql
V7A/Kp3pJBLpKiXiyTsoc1ItJMz7HlXQ2NFTfQyZWfvfCcLtEJgmLsxaDa0/e0TU
0MxOZm1yvz+RaQe9DAq+8JlHL6ttKJl7/KdNr+a3Xfi5s6kfSU3GiSd/ZSDaedg6
ZW0C7Q666vYnjBEkMzehXMFuOQsiUpJcfA+wVzru/wKOHNnsHqwFiLCzksnovseU
9qzI6XwkzJ9jsUbLpJrtziuXauSNNHSBO7CXDmARmEg6bK5u6DWlCPaxNx8a0YOm
c0e2n+KjU4NucfoeTkrZXye1S5oB9WGdVwrSm2iKD34s+lSCv0HBC/byt24YZr6x
uV7VIM79omaAz59EuwNdA+URz3aLU+SfI0Ws++LG5rkqN9sWOcW/Br7QT3KB8va+
WIQdS5UGMLcPzrSTB+d/UTavCKALEY/DxMWN2YTjdH+iROP554Ony/Zo/ike5aPX
tnXoSL7ReeT3xy8RoP8oZi/XGwhDNnwNxO0iavk3cLQb7VMTIJ0vIRxlCrSWA2Z+
8Y+9kbXlGqfLW4WxHE9Ui0G6YumEF8VvNBlO0JBVgMnPf90tWLZQYIa7Da3poZtO
xmo76hX+3DjRSkpw/zR1HTk96Z6/Z50qfLvHKqTxhtGRDv6EdIO7dQMaqb72TJ0J
6MpGVPt2jbm4s7wIzDsBmFWJDlsCTSHv/AeNy2vgm9Nz/5Ndgh5oLgXBqMo05GM1
5+EnFFRPJbAc7c6RKRjh68qKcokRBWeF+bikuJI+N8FC4r+fQpCqHCdxIpZ7KrVE
J1xnPNpVYou5TeJTKCPXLLKGgVQnorhO/EY7spjpLQJZDidMdn96fa2eR5LjipoL
cfapZRddv+S72UXu5eohqeQqdpd9MswMZL/AjaCr+Y13/esSECAlhHnmf7SFKtas
rSBuahWOH5XZSu7z8cNMrbXgBIrfhQIDTeV4tVaA1DhkCvQLfApk2Gp+9u06seEN
Q5oiFY7NRmvWpzVA4nDK4R2MVA8iZVlVClWErm2ugY/e1Iccs9gH9gGdyXstxnZr
VwoO6BlWdUb7OMD9OcVU9zsuWZyqL2P5oEy1PQM+9bq4qqOWXF+bg+XacS8vrPox
9UDPpZmpKKjQLmf/QT4qAJLZvGz3qEu3UZSfCzlOPUVJNUD5jOks/VLlMj8G0LkE
3Img3pYPbnq83MzrS3JCYJQNzKfPXD8fz4FdWRXuvTSF1EziWrCYNOkVCyCY+5MD
zJeuoLq/DzeehXipr7KsxJj7HzgdufgQ5HAhp3X+RnnREeWTAqGpmi8tpowPJzu1
s7cI8t+lTlkWE5PgL7lpy3odT31pjkuX/DPBKkLJby9ieYcfTdrsPshwqaORwTSG
QDI+/nT1NV53luzpLiF+m8awPPvSJCUb05YmRZ4iSOmS10yAcf4nn5b3myzcVaEH
26yliia3nmZb5ZztsV1DAHyaMnC9dbfQ5RisqO/MXR0R8mfJXN2FBdpPaTgLI7mQ
kRvMfRtavFFYPYWmqRpHjLxuWT2ybgJHqK8B5FeSJ2nCeUliFf3rD5fU6J+ewNfG
EBIG2NYDtEwgbNZlH6MgqLCBjY2oNkdyOIQ3UYe4VWoDanGvxLOisKhVKjip4kIQ
bGlbhvMIFv6CktIVbP2UwN/UbqeTe/NkhZ1nd6SMXIKfSWHbNQLcJCQqBik6gxC8
ZyXGjByDJnV0euTJp6WxliBfovAvDvsbnCZeGyl/vpaXTWFE3vFpRhL4mpcgt9f7
HZ8Jko/6JRtShgLsr6Zxykw/NBIXyD/pyFPNL17lroNzVxHpHys09Nl7U/3kdyss
WI7UBqArGxyUH6P+gDLkzu8jTB5YTO7PiqCkFNC9b+fTN5vuW2nRjtMAw+FaWfrf
O1DwXrtGaQQwOpRBWtHz8/AddbTiniv7DRMpRfip4INYF1VOTVhzBSI8m2cDvqpF
2APAJGPJaadKM2avuOiEsu6H/Zjf6IMrqWHT0z0N1al0v76zA6leSRMa3/Dx63xZ
21gBm8KNXZc5C/2zBBsSX8VjgytsBxdE1x164pmItGR23w3G9TSN8OU2xfKSQGF6
agrnH4paIK8+7t1fA3lhAgVHCGYu8CRX6gqCJlNPJEHFnxXjJ+597LbgW7wcFEeQ
jr9UPGb7J3Q74KUbCflpgfWRSWnjxsYkPM04HsEal9unH8ZllFsh6OeebvtOG6ut
8rkA9Siy96Zh9BY3pr7nTejBAA3klZ/mx8fSo1gt+ym/LIWFbYtvdSVbHgJSwh4y
aTmnfL4//XoB0sQCnjjjhS6DCVgZQkryhbYCdoT7zF82eQgtQ6LW/Dxhl/cVslT5
Mn1W2GfrpWWtSKoxJyFTz+pL8NW47XUl67GGO45fr6DYOEcsHzphlUu5yyoNfJxp
29XRFr0KDSMS4CwqYjJM7oEZuMdqmfVyDu59hP7M2vSFgYf7gtprhEONWI/1prVo
MLE3lN8ykOhNlt7b0cQ1y0+KXaLvuD+5c6hGU8G7k4Z32oBQ9ZJxn18yCj6AE9CD
alFTC9hVC5fS2vMDb1X5R4LcVfG/zjVW3jI/u7X3cuFAIooGIXM5/iirYUMD9qiv
VoedCFTm+9wFUhPNCwJX+qzuoCmHsjTEvCf6YGrWbAMZHvdpTwjHZcDTkhx2wtVM
fOUIg1xIt+KQzJRvsqss89oJEJiN7uxp4bK5iPdovwU+s0/TRgJyCsr9Wy4bPUIz
PMPr5HNagoBQZB0+P2J2lr788P9amrjvQph+V0R04+PpKHrq/IJY0prhB/GbzHIq
P9Cjy03XO1lqqwjsJH/DK1rJzH0rzOSucx/cAX/A+w5QK1jmcflfmrVGhDJQFuDH
6JYINVyAmjJdo6HKj96QUXNP8LMbAIfroOLdg8NzILEonwCJYLc+iHMTKdK0BJH6
CrR/Dd0I4fbWMannaqf/smMDre6SYJjIsOyOMMScCyFGjXHH7Ftb1yHRvQ5e7+Qx
a0FGl6n7kwlBaDTZpecybM3xblefl4+5uhDgqg1zUnK3sca/lLYk/vDnWPEWCyHL
uHEfFIO3UPMjzdd28Mn1x9qgb3Y1nVDjmemXYtPaBJJFiOir6/l6zl5dJPx6mp5K
ozcJIlKvKODlaDsaBD5gyiOlnWn7ktNScIUWgIP5ASAzfYYZZUY+svdiQz2nXkwD
M0b7KFRzv7PV8FobjI6VBiup0Ac21rQ87dvKw+Agt11i3JjL13Ha7JtOS7P48XT/
mjs50iIVgkAKERs8Qyv2SczWcws9Vy7i3KSWW1cn4+JZvr43cNSNwpk/oVaRKLxs
op+GP76f4Em0whGvpVLksVLZlhGOPSlKt+eIiI82EeIwcuNP/ugLTc0Tu/1b1OjH
r72kC6XE3p4T/rnitFBnKR1znjQoT0be8GIsvy+9WmlrreMRNuohgDDVjXIrarOn
wmuH6v7+2iOsH52CH6P9eDJHlqQ5nVnICD3SRnfWawKFKDCHCIqwkEFfTBm+HSuT
9vM62tRpa2aXzsLzexUa2QEnJbvfOW0IbDIHfP22zpC4xR6BarhvwKVuiQTTQWJF
kJ4dAKGGuMKtuFeiEopcaFC0GVaJ0BaemOW4npEZ6wWb5iZHO4xVFi9R2MnUoU98
b8JrYUDJMU99H3z2g6L1LU+OfLr63GeVELiBtNYO2J6JGnVVC9Flt/APDy9WlIap
ep1levFA1pCpSlgc6NbmdFXXJuXpvoIlwJBo1SphXGGzU/t1+uDS/Az2t+yW8hTR
2TSjWhs85Ugef0Usd1L6++LtgkfMGLspZO2nQqD3T7DRVwCV/WfOZToSbdAb8t/U
1TKLbgZTXK6bRsnvuda8Dn+wvUJlQLHQTqhnq16Igbqve/ky1jw7svUJ7vZqbeZV
3jzv375XAQ+sNlLIA0tW/MCnBk0xrzFCAcIvqRssGxEqsJ5QwhZrWvMAG7SZI6YT
WPBfqTdHm7OLC7rzmVtXFzYGvHsMU3vmOLAlfQB1j0mboBtuUU8Sa2pRIjxdoWQw
7lTEE6a4Rta4WK+y55+wa7ThcHswF9BNq0zd4Foj+FHMA6ANmdhG1dOTzCtG3Vko
UgyMZvJ8FaBpD6pcj4rvoJAeZOj9LnUC6nocUhynku3vJiPDDjVyvCsE2jYCohjf
6oUGb4tiIE1OzShh+Te+ZJNPgxoVSF/dcop/10V5WwJMTNdcvyl57XLv/ysCemBI
e+dd3dx0BNzCanpUm4xwgYYi27w+0gLKo3mlIa8WZyxn8P6PvOaOTNQXb6mRhe7j
XZPu0xvsIrAA3K6WfhMLG71wh9dgkV7hW25H6g+/pYuHEquWH6ZS4p3+h9aCBTf9
+ow5sGA4t5/Pdqb/xYp8NDfvJJgu6iHtMfyJ+Cc7joAMAEgsGT7hDGzQnAGJiHGK
7J8KGa7EkrDzVuHJd2K3l4GQurh/YS2xCt6z/B4fnI0qEW/p82Ium3XYavPCCulU
2V/zhjCj0150AsYV2lFppdf0leZ+e+dYM2btDpZrqFkNYabeu2BQRh0YVSzzAPR2
ok96Rx+L34UEj9xlVkadbZVAS8mf271t75zkFlHaFjxDably2kDPB7fdzs+Zwi6C
8OlQ2bR7OEhLZGH7ci97Fxr7nOhJwEZd6EP7lvZ7o4dF7mpEsXg+qadEV1dUOD3i
b/70zQ+WSiMaDbBYhi6K6omMZ4Ojkn2dQWNQjNIIWnl0Vxjv5GfUrlBS2PxSmtt4
Zr15bMHvP0Fy5eGrvXiNv0AeA4uLZdeuLLUl2oeJaOw7AQ7WF91Ld08tiFZMC5PI
EmiPu5C2H8zeOi3sAtRArOefC1PLizaHxa0kyJ1cXx0jw1TSFaZ8IX4yXlC88cvK
o77FYpYI55ht2jkO2BRCSAFcAtgWXM6WLDNb6h+Zk6wx8gctH907Da5eV1/74yyD
sxoAFk0YxE1zpG8vOJm8tNEOoS82mNPsgSsCWUVe4U1vmpcUrBJH8sDNo3aSmxyN
Aw8VqOq/hSvoCDPMb0sqT7Ae0YKth0f7of9DGnDkjY3y8HUC7sjsK5yZhSPrpUIL
+b1Rtlx2amL5UfMulFZXZG92nghtdtYGzOcL0WoQDPxHA7WA7tTq5HuPP3GsbeAE
l7GmDNUq9oUSD4Xbg+PwyHKK+IaX1eiL4ZP55w2tBG6dVlQM75i13/0q6HrxTFYi
NYR+ANWnT/DZiFE5TmxyCqxb9cChoCZ1/FaWxDc//V5ZIkLLEu+FJHq9xKbOjuDP
Z+5C6xqCKgfcyere9JiPOl+QYLaGjmbAVY8hLRLEvz9eQZ0zMSAUn7N++icjb4Px
C2OeyaM1uSW+t5E9tbWEMRQYeslYaUxIFLcCVvswTwA8bLx5QzWR3RR0LpOKGhJN
YWgwAV15pcWFxzphifvgyoxH27ho+dIVxV+hnlH0zHF6x6zWBMQaMjsKHEt+TPB9
3MXHz9BMpm2lWjqJdire49zL8PU+5kfVnFiUdOgkoivGAwoDnS16ZRxsjGybxK0R
C4arErc34v5DbmVzxtNi8e3ZdDhpk18lJZkdInkzqb+2sMPh569q8/uoB8Wpnmdo
xS5ZwogEqqvmanD611jrG6gZtjDVB2ju/KRgWyQQBnRHHtoOs99zbrM4ZxN+j3Vx
DaEHlhi1HebKUTky+YO20JuP8Z34B1I8/c9nzVeeMQw8TwyXUwFLiTg5pPyHzXWQ
HxXiNJ6RME2eOT0LSUsmxr4VPdpBRdHqV5oJvLVOlktxCPeMDj98wp731Jbs5R99
n1cn2Jby8E9mWXFrllsMUvwIzy4L8Ur4mI45JAiNExH8La8pMW01QMb8k+F1j7Db
O8XOPfG2hMsaVaOg5rDHgMGN2LoaS3pIXgghs2C+Mnxf+45Cnm3Iox4Djx2VQ7Hf
5LwF26GKkIjc4lAMUI3lZM9TLt6DA0eIwHCu2nUpBD6zKRRbCsjdhmjnjN18DCQl
QCzDTpQCJtz0GDOrMts3ucJnc3yZI0TZujKM16ft9z4LwWcCOsAeOcrnjRteo4ud
Ii23wkJboQGbfxFNf2lRuTMRY00WoBgfF5EjPKAMvVnfGx6K/e+eVPzduot2t0NR
2Gsy/IY87s0I/AdODZu8pW7UjmHAH+kxgdysp0Fm3bEigNQlJm5P8/DU2NPg1dq/
3DOz5Q8bli2R7irKF7TtfJgUzvtwLA+TqAknoXnnUQHv5iRDeWmoNIJgHznDY/oj
PhRNjDCG/vFMULorx2tvZFU5ppyWC8zoERcWDUHNTWvBVOydBYokYoEJ2TALhfl1
dkPCOP+xLLlGYjEicH6R54bpyHjsv3flAhBmWlkM3y5sekhN4pTEUWlDsfEMzm0+
b/jca8F9k8FEpoXjmZEG2bgO4dtW2OTvlfrFZod4UoHEwxuqV/uR1AdFlXMI8+1E
GlTmSnoVwBEES0FJBjR1IDqUd4Fty5PyvZezBAm8t4MwHfMpjmkguzBXBA/UhHa7
f9yJyTY85q64CGspAWFBJ4lZTjUE7aTrwh8tLBYgUCYoI5MawHguMuJVFDYxguTi
YLZvDG2LCTsyHkGBSnYTDMewn/sykCPd0af/NiGUoFSWnA9eSir8Vk+sr6O6jxbi
m0tgtT82/JLC3CT//tjP153JSV0bq4wk/0SWraSK3JriBYPMnLE1LoAccgf1rpkR
ugqzwGxbaS7ZgnHGpeger1kzfgysDeSTwme2dX0TY0r4nxERi86DCavUGOZ5Ecr5
Nqz609TzCyV3oUzsJt3Vi5q9mvjRdO/7pfAyD46Le8IjEgErbLXCCMJM4y0wvBGt
4mo9WBV66S7KXQW+o+TqKeQUoNmUrkKRLW4qCvEsGPwWhWU48P5Sc0YJeaqyuTlK
wbIeI7wQwvmU3AU0kjiCHFUJPpOJkxzVAoZs9eofd3idyHtoRdsB+Rfs6FxUU8V+
9wHZ2heHHqxGY0tvAbDbYD5UH/MffO5fWowz04Nx2kf4b60EINmuavspYN/TaW/U
bxCjJt/bUe9FiAVlC4op/P0/BkGpc6SOOc/rpuk/xrKrqBEDTE/MppcQNorSwQ0H
AFdmtjx1M4rbZIifMgiAls3SgKEzw+Xhd2Pimk7YpC/+u3tTbcdlTsTJ5jZPqo2G
dU8rdV/xR+HROAB/XkLsW2sImTEmYbFagfnmKqfUbRts552WHt/sjMqhoQUOBUpk
Pq/PhXZJCRyzrDHlHCUHjJTZloeePRRZzJSrwoVqDR8A1di9pxlPxf0NfBm2/Vzw
tGvgewQLCVpDMRZQCwnLna70CFG8PxnZAooMLtG0rtDEFoMaONliGehxh0qcbhLz
7RbqMd5VmzM7Soog6C5Rw2iiwJwW0OWJcKjIvpUfbRZib5n9ibymlHGbwb4QwPFK
yTvzMQeqFgVgA4QT11Cxv7DnsQ/Uh/duI0ixrOwnMZlMeCgWFDSuHFn9EGoxmKD6
BitNTPL4jXymUprwSXh78VMXHKhNPi1JV33G4VQfyuC4/JMJrRUGzX1rnIyQA49Q
hjl2n62TjOICywMaJw/4wXDcUp+MdIV6WFCw2yqZ5ER8CxbMdhQKAU1Wi2JTUFCi
ij9DRdTjrdx+YiJL9HOx7ZKniiJh1fqRXeYi4KQ2P+U8j8OILWwdtVyFsNAdyJbp
LJqgXfZ3GnbEQmgIL4pw+4ee/c06Q+9aHAmck5/x0OglSBMttLBM+zH4ZlfwZq5P
HzK715PERbwJajLpGH861+3R/h3rn//NP5DpXmFm5TP0Cc24ROM6j20A1Ff8W4Ob
mE/Z5vZC80DbYRj13UL5S86PtZYDhSQ6n5TWLOFYQaDfRwAVRDfkKT+qH7KOmf5I
UJ+7nRnj+kavGj9rl4tV4w0RAFBKF7HVCBalveSRQMElKad3Fgk0Zjc/0a7aMJiD
0LHtOUqQ4Inm3+9CuALd1nhaV09ReUA7uz//u25df89ZSBaQW7r6zuVlMp//YBCJ
mcM9mn+nbtofpJPPQlPaFLQEo4Bhqi+v9/7TvCV/hxmwNXJ0PvsUcjQFVhfpvcAh
X/RFCVvlG6tQku75rJhS3oJiBveD8EyeqiloK32mhqGUs46ne66yOOcQQaZGCKnw
Y3ziwzQTuofOxdOBt4p1SxEeHWxANAdfr1NE6eJW3VLBSJq6wJZijTZ4K3BuM9gD
vpixz57pd4KJWBcDZp/Sx0xYErx6q6GLv5d9lm7khpR4xgRMuBe0yir20KyRQt92
HDl1q9hEorCnwq+HDeUzXuUVyhsuEthr/cirzk4PJVpdMInvBPRWXTONcwPDphgb
Nf8ShlxTVN6RpX8qHDwxJXzGstfDsnocYv28xmedCLko+59ql9tbsVOr9TevSoBb
DnORWTIvRE7NSTPUaRlwf5ljeJexraw4Xs8n9aLU2DpxTxfS1Z6T85hvagwL1fwv
h/hHtFKtXlMwgnM7tiWnABzI7xTaOTCmDGa1VVF5R8IcnwuBYAADvgUXpmIcr0at
5cJVpHx7xFxSVGoJ+goiQ39yeztgqWkrLRStCM/2z8jJqarW11dyiZwMCHBKyw8n
XY/yIRIH2mOWvHE4J8uhy4MQfvDtZIZH/AzNrw2eYuKg9au8/oZpAzn82agtqmiL
FuLP3x3blixihBaVoitJ1teX7pNwCKnJRhJseKMGrgr1Ro2YN50Aj/cgYEWyxzK5
oWoGS1SpLycIQv7HIaVk4rJkX71CeH35zr3ESAlZut9KdI/jEIjS+7gCZbL2NNa9
BTuAlqcKKp/XCGbcp3GQx1/F3okAikZe5+YcguybhOJgWBzhGkSfEz/Hi/Qr/wxX
e6o+p+QtYw8I8feR8xJoFeMwSA+1EU4ZUcrgP+y+PUM7ZTiJVtIVtWI2afpmZWHh
tKVHPmZOMaglEkLAyHOl+j98jt02c3yFGiuKnIZIiVCRlhoS8gmoueGNVo0AJyLV
Ocpo0IMFNMYLz+psTjSK/co6oh/fgLLBAZBLF0Pb8h0qEsBowvkJkIXynLZvYLdi
iXy0EKPdjq+O3o3KxJ2h2leEk2O5JSUfuYzsdRyUrZe1fm9nnfW4tnSGsuMKZcxg
P3hGUGy2wJPaXws6WewzLTPY36H7Sk5qoV7wTWz+Up0LqO0nO4+DHPa4Jc+g70KG
eGZKppJpONqW1yWqDAUOF5W1vDJ1sMVz+F0B41Pp3V+BYBwFeU/7OSQv9tS+tAc8
wse8swJGrwCPZxnYHdLlRtVoMnnuZREmFyKR5Ko+nYtER6Of/X0QssESmutG02om
Dkx2ZYCOf0N2Y0/9H5a9fK6WMTNTYIdzxsu0BTltDVauAO218o8j3aHbyFkD/Kr5
ux4rn0Ug88oZEYxk2BXEC4921lgW8+FI92VDfLxwQ/pzpAMM9XG4mwa3VP9wN26V
vQfsSobg/KmjryLKVJ6db/APVilQug4/6i9hS2NK79Hom3QUtfMQAAmMuL5+Uuu6
9KZGRNgqUnBRn2jom3TdoJ8RTI/LpzYwXFoYFfYkSNovTx9hP6Td1AtglDSJnGCl
AfTIsIaxyAJcD7ds0OfM6CO9G12MN3o0mnD975ygJDmEpmEZ6frBYFoF9tr3O3iO
9QiUDnSefGxrsUHH7/hL6Xt+FlOJnkXZqzW7rjiazmKGZ/Bigk82QvXfgrIm9cDC
NX2sV2QY5lVVBRmdUneDnMfFw4QCGHCFiP5yCBvGKTbHcOotU1tnCiawSWP9GrqB
3qIbUHYTpD+rohCOGgjOTGdN5n96/GQ7OsRYGpfgMw3CFcafQAJJIj50EgkY0ZT/
+6XwwFTbU5mMTY9BxSDE39NfmBklYFkGs+cm/+ZBtBDdBzuEQfVvGzA7RDK40vCj
fTd1I2OoTeO0SNj+L95y8iY/HrvvfzQTvz53c56MUi/B6TW3ZLJTZZA2I/ScTn+m
noHYGwHKQwvq3QH5iqkaSNMUvjh7k1hf987vRwe/lzMfc6kT05/8XTFICTvC9wT/
1SDnvT1Ujf10l8I85Lulwmev7HteQMOGwnkO97s5UZt8yMk9KkdS6Y4UOhUE4IQ6
putRBrfK0xZ2PBSZ6KaF1KjS2hx2C7gFsA4cuZgXhW/rMPbWnY4/VAqZKd6bujYK
x6ELSnbpV9wQGRYie6cD61aihbsHzhMqgt/bWp7uZTwVvGccCN4A2BIx7EXaVXE7
siOMwL/nLrVBZ+i39Fpz7HHe7U/cWQE7eTRd4uDfxTyaR4fcDR1LAAmaRsqRu331
h8xnPz3pUcQ/IYpqGzuvENBZFmrBhRA8r3tQB27SDBtj2sZaip99HlxaOT5q6te5
e+vULaNeJwosblRW/R6OaN4bICw5vbCOV90pNHVhvEuJR8W9BQqS+d6URO9D1ZuS
coQvGt0KUx5umiGqFAStsA7Fi4tN9z/0dm4oPJ4thxE9QFe/N00q8PBZ6RPGH8ZB
qVSzPSG0bT7Shj501fbKKGxKh3JiiVb4wBIqEY/je+d42Si4aV/ROxZvoZMIc8lr
qL2eghnV6ED5Nxur089obDULl0J80NDbIBeYgPJf5FM6GI2YY2b7xQV/czDQCbuU
u+B7UBvDgPCqw/yV84EmB4L7BOS5zIxyaBRvriQSE4Rp7EFaY7/kUMQowCjL7a8x
ZMw0hGXc4fw0fn0E+ONTbkGzc4gQBCmBSoHOKJGxsQZL+U9+Dl0wY3C0hhsXSEnq
/sn55mwfmHHMmo9wseI5XBW6QBi3w5pTJ7vebKYofL9AnTpNETmYaPXGcYTi4TvO
WVlqb72pdrjyYlOqhNEdTXQz+3IMsOVehZccOel1VRpbCr40f4vvspVRkmjEDaFv
p6DXW92Cy2HI8Mn81U/L+jv+snRIcTC0OmMpfIqUMDcbwRDi0S98Oi/COe+3gYQw
ZPzqWuUTLtaCCrzF6/WxfvtW7lKdWu72aq/4FTsiM/RySxnmdpP+qEVishBUwOaL
o9JQ1KX5fFrfjwCWYBjRThH3Qg9pHe+g/RuGUFjD9xYqmqIa/jKebSGVxEUy6iVQ
xy8NUhtl/fGER82iC8EUHe1dFS0m5bE0XMzSTEQlDjAjBagBHrOq2xQy3UhK0KEI
0uf7klI3wsa4sdmtpM6rLOCmRww+uEBQZgu+qJdSxXLSTTZPk4GNu18mnuJ5vyZj
WZ1GL8XT08YpYvlqJ5fGs1sbrVlcN0QUWiks6mUPIACmtCeInxLKRzGwlp9WYdc6
WB7137KY0yEDwyWd8arLLvXQetsK8rbo/QXbB8T3g9Z1I5RSYeL8GRsERYDn+tkp
nogVAW7smvXUaFHD5CoDk8wXDdLAjdFwXNLz2pRnCvnC1JfyURUK7KphRFxAA5p8
selbTiNCRr0+brRm7Mz22m7F4E4EJvyAE6V062xbaa6iEa3jABwbMZK+FE4wVBIY
XAw8vDkLno6Qoe9g3JhHQhn+HuK3qT9ZnvVSFBqZGjUtd2DA/rVr59CZULaINNro
TyHwWN9s+7j0BTe7xCg6gmS9rA2Izpq8gO7lQ01USHvdduQtNEf2i2XC8b1lErVF
NhnRWeXfepTA7w8iChH1+wyiy/19uPthwKA9Qf/d+lRazpQeyawqkA5LLfcg/Oia
dx44B1iop4E/YwSm97yeG/k45vI8+CMnCwLyfV07OL04qUnAnKC4468ppKgbMias
fVH4Hh682O52oUzrDkrHcq4Yx2eIPN3NX6CMIrRrrhRFO2N/y8q4xS2wIJhvi8X/
sN/+bVdBDaNIjS2vJcDAhs+m96cLl2xjjszT4gQrPXWUovuAFSYe1DJjHxqcqwUK
nN7MdTlo6dDG9dPXZzqYAuphDVKhLM0YipIb72oDs4Bh5tHkrCemyu1YL6Em1WXB
wTKB2883ziDoVd9X9f+KO5GN9WVoqdyy3KpWlAHR1KmDDyBuzkyrilD7v7cHGFpW
Awi13HIhRyeHaeJt+iThxIdDDhH+MCz/BsZ5R4mu5gejJ4ZiRIhazJbQdM9oAGKe
wYBx3pnxPeGHJ/MrXrZbPjMFif9Y1PbpypngOpsvwemoU923Wo8239EgGd79ki65
oacTiWP0yXpLjs/zThH+e9YXsvTVyM4tOeQOEpbs8DeLXOH+bKHYTz0PTgZZfEFV
xNVUSQ+u/1hF9+Cg68IkroMLdvNaFiXvf8p1BqrvxdMz5mVzN6f8+6SGp5kdTykc
ANKPNKufI2uNxjGpG+QnmcjXcWc6F23hWKd4AU1fiUMjjWNsczA+bZqHz2rUAxXc
Tfi3DpkBpA/qhCfElezDhcC5hmyF2iJ8SX+rS36mclNa6HeUI60b94o2PzMRrlGH
kZn+KLvsf7/zDPseEkir0lZFnzhWRf7BSldPVv+p5iRV2ZwBt9O2WtqHp0+WF3Ff
19HwwHoQ/c7i8I7WKaGLz6NCsJ9yOln1TMP6tE0aVhdEvbFJtc8xKBHSiDeyJPR7
CFp1lyC22RiWME1uPqivvYTBb4+06Y5Kh4a8Tou6NTL1lfaAEikiviIpFA7mvgpA
duBsDd9mgcezzyJetmV8tDI+By+ZeFEWgd+GEaz/WspjilbLyExA9OgTMCoiVAAx
xc5uuOoSor+pyg8gT/mtd/uHHO366KvwKfQfqev7MaRboax+1rTCkGJ1vgKpyWxg
lx8LHJT+sBCxkzQhO1MdFJtCLUyK3qaLIaEEhznKx/SPzrthYxJgSJhl2fSe7mRS
KKOBAO4t2etb+4K2sW9f3/0cRUmshwUg4eaHEIVumDR32WP7LT9hrGpCAT2pib1U
nnjdobVB/UTzg4MklM9ZWZddavErUk0yvmTVD94xugl32IPkYspfDYZRydbd8qt8
7ZV9v6i4ldp6/0h2q7G05K0PRKp70wkRkeEerQp6qV5qcfk0RHnri8DJ9dY8moNI
QMrpER4B3m5fVmHi5Z+KId5kigi6sUQMWwTouayyOdv9GaFyr8N7eNAqZ+bcoxGu
5ulxJjm3nhSof3blMawHxC3sCq//DzzK+3M+04gqKjuh2vv2O2q82RDOMtpNyRxh
+wGSWOE5Yj0oerc9PAbJ4yGFjQIPl1EQ8Ry8K0G1ZNtE0BtJkwicTSi0GQC7SCTQ
xwnjSvchydnmGbzRRcf1nYwaljG/3AOqNXMoHOD4/8s29/YuCIoCPTc9mmm13E9C
OR20uxFs8ug4aauX7+/sXQU9RrFH6y0bhkVFdvfoWDoOSAGDQMXxOie7uyr8uydN
RwCTOonlsIp4a7nkgM5S2lO43nVVLqi7Vy2Ccl3ncXGNKzNAAJXD5mYGHiPNWo0A
m/OywjnYxpJGnShgabYPm35Mxs4VxUZLIpFDB4GZleVMqfpwOmvDMzqWHfEHQ4ui
QbNHyqTp+PoI2gLzUWApgCVkJS+YGajIdQBwviuqtjMbLhl3nwHJAW3IgxWBrM9/
USJ8jTn2lfrat//slrGFN+SkCpjiXjmmfh861wjmC4ut7irRnYEdYlIuwCUlGqGX
taLRrls0WEH9jmEbwtz3daQA5UbmHlxavkvoMhFfArw4N6Bt0vjtLlyW9KM4c9I1
MK4hUnawOAGFmje3ngPwHOjnNxl4694zIbAaOCIIwi35d+vNU/qtgnmnzC/L+b6d
Qw+f2a5nwQJjJjH09SU6pa5VzfHL6ViZ0F/zXdu9nGTGwEHV0SY2XCJ+49aYKy14
oojtppSBY/F/gkZkL2lj7ZbNVDaq4RQiC9dcX6A8S5E4DS3WZ8ukkKXIV0GXrbOB
THzd3tGEey+jWxcrCvjaUf+15kTzG9sW3lb2utZVwA4WU57eKtJEw6+6sEbjVlzx
C3El4694ipHkhVHpkjsR/JLm8vL1ijamyqyKXcNwc/zoi0eBXyUkXsbWyQu7ghjN
KLyixV3sz1I3xFnl3NidmiOAlzOUCWIJ6aUDEKrEJrocbIWFcw+mR3HmOvPObxWQ
ldO2t8GSmDJwE7BxlYiL0tnaBX2IifS6aiK+PZ8/cvvuGCKxb3eV6g4jiGEQ6drq
KPeKklHEtiwBTmMrytqEx+htgGAbyl50YvefLUCzeY35UhKdQjY84UibTPwbPFtV
RExuAt0HdkMQpo9R+hMKep1LhC6+WpLRYXMpYUNfh9l3p+bi2bUmUIcurkhqnWFc
Y2z2/ApGCQXbPEfjjF11RRPVcMmbKWVJEk/UeYE08D+zxyfJ3fkzlXeymYUUyLSW
mOkx5WpicFcrYAYWCDOslR5UOpKhzpqjeL9t6wK5SkjCZaOwHm18XEgZETPbyaVy
DQl6pHERN3QJSPphcDLA5+THQWhMNHBhtJYO5YpG/WD7YKXNG7h7KkuqiklMQUYn
r5S/IFCbDgtk8wJODzgLbdq5odmobxyllZIxX38bklGRVTPsLSaAicm/kZYSrdtY
dF1b6cezL19C1ClJxjG7NXxf2ZzA9MkGcvDEd9GcUx36KTRVlY1hCAy+j9wnSzef
3oG/j26UyAuIZLP2YEnM8phI3N90nENIwOEQl77yH4PzzTcQpxmUrCPo0sUZX2h7
9lTOJxaM62c7mkw2sii2JpUqY3UjHMcvRy2uQjRSDKxcYNDwFG8H+RZrnmYXskZB
3xPeQECGFH0mOeVZIEJ2mkaq68zccdrYe+JS2Hrmma4r69S/Xa89biopcTmCbEVu
uPMdkQaIas/XH8FLVikiOSggbbH+Kbp67NbnzUmdKmag4yHA079Yb1WB2TKOTfNr
TuNDujmFeweX5Tht8pKS8E7kyjZ5YHYD6g+GINLAhOTlazp/0EZI+3C7Dbi4n6gA
PTZzTtG+8aQ/UhFYjU7UbHV3l9YIq+R8JFu0h0gKHZCThTdPeipNZ2AVCtH/AGfH
24Ti+0AVKZzkenofkPyjDH8HRZEIArp05XsX3+vxsL5CEjQ9lX66zA4mg59GNWC6
8yDW95fwaeD6gux8ZnW0pDHDMf1o2g9+RY76eTVplw3sTx8lty8G6Iyti1cFsBU2
LdP7qEcuX86xrUaQQ0cRAT0Hsskp2axd6cymzpZtqniA55TCBpWOj2ZlvTwPWSHC
aSqXzMi5t1CuYeBbPTTt52gHVO/O7N4jDG7YZe97yUC+PNCvFmj4mhOLWt5/4ScQ
bUEA1prYLw1eubK/9uygO5gAZwUqn/RxIudkYZ6fBgjVlOcnl7y13jEXnL3H9sha
RIYi5UB0k1zRuJSDDAbZvSArb7aPqr0T74Qgiuch5PJNT6v2IPLyouCjCfWn4uT9
k5rOLJrFWJj6zC6s2fHSrvp/DjzkRYvZYZavOYMbjK9D2Bj1pBwkfW7DuoDOq0za
Xj8C9JdA0vD2WA5i5QX2K89+LhA3NtYfm6uYry/KFddta737b26ORY7DLQSz3rQO
Wr3qJLrXu12glKjC+xcbZixj8VaNrM8Z2qdPY832bc923I9pKEiKcBEs88bl2Vkp
86iFEDYGBwq7EhbAyb4oNR4Q2ncvo58wi6sUiAyFy6odLGDnXQ35sMdD8FwrksS5
kVcKK+EebPsV8ov8BmOuvxdJ8BkL7C+z2lCXRmu0oPnEDXw+/KnB2wMYNR+Q8sEC
4gr3i+PStBLvNZyAAASxtvbh+I5GMAv+x+zkvPHXxSYXQNDJxM5cDkLd+njN320z
BK1PJ6DAyFGGwJAxx+l8E66Aw5KTLklp/EcW6+2OBXEa1UdX3yxidSQjlSNREDRf
lsG70eeQ51YI0aaQ6BYglbscy2U19O6tZPI8SXd/4OKO2AOh2urBujkrGfwvIRmT
kQzz2LH74P2mpfWMtMHJ32Irg4s+HNxOHTRxYjYOwbKglxLqs1vWMiLvUywTHJCN
POjYbjV4oEX9wjvigr/96f4Bz0hiWBW23CWW1bABym3L7aKiY58JzgjjJohgxVVC
hJenJ+TnEhmwreHdNRActtEWkj0zjRPM7GNIJqHHd5C4vHhjktjW2sfCzOmsKIm/
Vyw9VLP6uHyPg7UFlDBsmLSDT3w2YY8E3bS/LAb0gAMO32EGt6AxO6M5GlUmCekm
xAzfG0qaWapzdSbivyD/4v8OKkQXS3CGy/5TATn3EHErpx0DGM9hAcVejKsqFrsX
XEGJb823Eq0rSx7JC3L5SZQV3NEDrFoGH6GiZoaULg6mxasfju2u9Za8IOnHADYB
J0wsSF5qca8/P7wY5LUKf8fHzG0yyKqtq9dzDECPOZd9NFWvEkrKxLEM+fjZwPXh
Ew8YdQJ8ir9GEQUuDl4aBsxfcefhNxS6ddxohP6/EwFKrEr5reGzK2J/Rp39AfcS
bAwuELp2+Yp3kMn1yFYKQi5SmVGxOYIEUmJEvuWjZVcCB2yUG+UW+gLauO261yNl
chVxfJfIJKGweVwLTYtKJ2aRZc/W3BwGVt5UUsT75aGCZHRQ+I89905s4BdYhGcK
KzZ+vSXKKogz3+iUk+7sem/6vAYyC6OV2kzu9quW1KRm17eZP5ETJKRDr10uyorY
1wrJHsoRD25tmSApkee0sf7KopmWkSmKeau9A3evwsY4pBaBGNmPou7qldszIF9F
gufy0WqF50DfBN/5T3C1pV9HTeUdthZtLB+7ReMypAqAbuVqJMm/1OIyz0Lzyrcd
6yWfgHCjewjmcBpiJ9idDcAfzH8E/CGBynRSwXW6JYJFkvVDq/N2a0Aq5HH+ohq3
XuP+6xikw2hvD9NR5PXjJq/z4EA8yz05f/U1+PN/4Ob8Q57L6PdOkvIBNZhGFd9v
DNnLcl8+MLY1EXy12RsTyTF2dBU/tceIGU0P9hNFKxdjHWY0e5yOtNZYWrBQAVn2
xrWLaOV/QDPVEoWTfNCmUE/tG81h9EXacsdsYeXgKa0NiZLT5tCXlznECctBX65R
yWpDnkrqViVnD1Msq5H/A3oeacM76wxgNoKC7MqI8DUpNXA5z+a/i6Xzj/nH3cMQ
9cM/1qSy1/eUJi/Hn5r60S48UXXV9YHkQFoQoDjjEpYke6CpGKRO3BOOIJ8e+gIZ
reAlxpUHJXxbT0Otkbr/BaPqq8zSITbhMNa363xR9A7y4O+NlMkTB4GEsauwe9+Q
qFKfkJP3hy1CMtskKOD0TgUjyF2yhzm/IaLRpn1/wl+9DBhElK0etXJXhkytGgSC
vrX3XNyVVnwfwXUiibsGoezmhI0Ll6Ckaq52KyqWb/Dce0JH5FRto3di+ztPsXtE
QiGNVGhfryDnAu2d1LzSxKyiqvNOqoJWFqxMEHiWGlI3o8ZoHM/CK4Wz2xeTNUmv
xuzj8jzGF84T1Lpl+L+NquBrmkMcijRXnae6/DcsDNlxtQDTRUaV2nYg9gRBP3dX
xWdB50RgRg2oFhueNJjylWx6KmF0kb9b8tTTuES9I4YJmjZ74rQJne6WRKnW6MXr
q0/WpXgzqwfWwM1w2qdo3cY7m/dYe7hAsORLsVux6IB9086SxKERu7nVQEXQO6zQ
QTA92NcDAxPIz1/Iorl1UJvNom++VLBv8O9TKdXCZ7B7Q3fm+jYzOETMpgUojvkG
sy1VCUg/q0xP91NgAn0yNA3xZOavqWGkdaN1oLSsBWN3/BWJQ4x9he1oZxITblYe
MpaiV7TdelUoOqioYlOfaEVhE1/m884OakFOILpN1VyagU8ym+96sQcV68ld8KPx
nhMqL6/A/yCy+II9CFSG+2t696USBjdBkvLXoGd1y3v4ytAFmo0NwWSmZiLrzOhp
5QeZuP00N5gttSYpOx51tPCgCFC/6C6tu4KlqJgqpNKEFe2WfmWdQ8U++qcwd7tJ
P8bxWrgvie3OTqzhx5zQF/cF2Gel51Al3sxjvcQOwSciRuxFsCY5rYlKiuPcXpcM
msNeKkTmk3MceAx1OhiPWbZRy3xdo5JwV9pgaC279LS3ZWjYTtSwolmZOkPvhHE1
64ZlHV65S5o3Gle7a3TVyjYw16MZrU5Gk7GZsmSfEIF16zvZerLbNnPP93Ycc1M+
0SVOMsvtzfxHfzifN+SGy137lf+oH9G3t3trr3trLGtAe3RTenIZmmVRobxRdJCz
x2IynSgtZkeUaesF3H8q2WJcPEVlErNdkz5XV0hI4zFtHXjY1BDwgEb+BznpnSUW
413rCDSZpiIk0M1guINr/EHfpIao7lMYmcl2zvt+WSMygG8Pxs/1DeaC8m4T/zzp
8cMIv2USjO6P+YVOcjwHF2PLphOyvGL53hhkpFc8IYAZBzEguYOazUYpuuBPi/h9
OxgUjHc4goRUTRZMiPTVD+qAJjoSf8YbYwoFKgXY3pE0G1cGXAkrN4OfYdXYfnGb
cDBo8JtIa2bPsmVhKlEpRw7JUPZiGT5Mv/AMHr+CrJgIbKZOqkD0QEgK17uqXCBr
PSOMPOghO2ELA8iZxpo5eeDQrq6E3YFNir/2FMsD60vKIGWMSttfj+o7WnSvF56v
MhGuclQ6XP7HUS5I0LcpNnq+HMQaqBn7e4TYyopQKCiUuCOIiE99mYoH1UsMO4Wx
fmp11qm+kcTv+sCwkUM4IrsPI7pZp6LxiV3meJslzU/UqGWFFRLDGa0vGDW75q+1
k95wTKL3aguwaPGfPgikc/XOSYd+5X6Htf+DxYpk7B/JUo10ndtQFZN9M/1rJB1I
ICAzb3s01pP9uWHeknlsgZAYKjUX37HqsFY/ikSq4JWDEWXjljrBAAc/exHZ6URV
RxfEoXWYrvR1nku88eZv0Lf515HsU+bkfH03Necyj0qr0VpKhLeklqq2siJXDHUy
hql0kzI6g5751pal8LWlhBXFRUTbKOHu7ofTGeifEMYOBzGZT+ZEjv5PsbUxhsqB
1YBFo58wRGVqzRQNYq7AtXg/kHGazUobIKP4fhJWT1ZzwaMX6oo87j0tKLgZEnbR
zH/XkBmW33hUf6GtF4ErJiKKMRHyv3Y0uFrYxEPYooG1CRGEQHw+FUx0MxAwh7gK
ZRF8FeEEGK29buNbQjtEatQ+XUbmUyrCT94VUKyDm8M4kWwbc67Rb5almGAM5xUj
I/8V+NIgdhJbel5pOSC3H8vp+zJl3/wGBOUltkV0BbCSAuFVjWpRnfD3fjoSCVzQ
XkgKUHDonSu7xGC7rBS+IS9dhUMyNIgnCBsi3AtXLSJczfAbLSRhKlM3ZIEV2HvE
3kf2/uk6V9XV0/Qvz/og9SmSiNZdx0m0GodIvboDL5T+f6/pV63gXZ1YImAGfHrc
MytJHuIZX2XoIHIngQQVjk6LexepCf/atiwk87CYYaUANIfjmWVeKvrY0GsNzsKZ
PgvLuC79RNDWi4Jy7Vi6acgaBSwtGku+xME0mXbyUWBsMjFeewxxdTcJIOxToF7d
ijq0ons3cwK367Y+6NUQGieuSIi75Cw0N5w+d9LX1DUKvFD6OsUM6Y9PDgAPMSM+
Aaww6MNskfbK4wXm7R4R4oe4mOllO6JTlrj/tY3Xmf/HDd+vQUGH6LiaC3KwV+Zl
/0HgYu21BxmhELl+3Hj8akrtcxHkCQg+p+hySV6xx0zSqxuC/kSsAiiIbpyZ+FS7
ICEazCoNFNEyNu+A1J5dlstjg2g/KhQOHQYkM6CQM8n3teWU7MNQ4Cscudy8b1lr
kP5ndC3rF3We2u08ubqq1k5ODdHiE3fn/yTL8A5JD4fBg1cqQ/v1ujt/6NPYr9TP
7XLwC55U6LXnH6EEDMyjl1JQM3jU8pMFkFzsLKlVI1kZiVQX4xknUIosD5NHoL7N
cCwEcF1kbLsj58jxPahZTQlqMkE/Wn5d1PlziuTOl4x0SeZNpZf8fqS8918HI487
Vj1Qnc4VsMhVhlH4cJQrhu8IIhBHb2soStToyIxRTM1JhfEywiCPNMBozEwV2D96
zOnhmVS0Qf5P8RXoGqP3Tsa3/fqks2+p/P3tRWIyhZxW8OJblySHUaiCfV2DcGCP
hv5tQ3D1NegEyv6ZxzPtc3i2MLioOXLCgLUj1uz5RA5airRTp9AtHQUN7FZs7g3u
XnNZYg47fiGKP1O+wielQ0Q098ko7M/iEhVokb082SRMkO2AB3KHPigngC7UPGeI
IF6J4zao+pTAgWIbeIUv74T4BWguobwXOHMWBYS0/WfKhuWu/zZWZIShnNhwCVAO
mEbILs2ijYlX/pR/0NY0Vnho1Xhcdp0jCeO4/bswsQ1gx3THxHkybHnLa+w+ELYZ
jB2ZlYHIAirk4Tk/KvTYRXrxNN8x9mCSmisrvUBHQszpkV74J/14H+dT6K4lk4af
QMj660EFuGb3X0ekOBnS2pMBPCNaaPBF6twwAbSbJKwhRmpT4MmoFOSIuJxvaP6z
7EionVeHIyLnRxk2VfzsiBYDuKIRmDAD2VmjSvy4GSTtQS9i27PtA4EdNMfnjf7X
ONBtXXALXtyxVjwbbUS8r8Opnmg7ECcJXeEme7nw6LqBz6ety74QkjMo6v8zYota
SbemIBo0q7D7wvonvw5oi19K2g/nQVocI6ACeN5J9hLIE/rPiPhc+evLgvQEa1hn
gPpaFEsRp6f26In3DR5Ewon9n888RF54bZb/3jw8+NeR2xVVo78B1TDjiau2coZ1
k0eJPzjDtW8W++W+xj+yY/o3WrR2zSGqOR+hC3d7tjcs6wKpE8JeLwI0md6JhhDE
AbHLBsjhKls+pdF8dIJSvjTULreMXvFETSkwIfi2FTwfndpshBP+849D8IhWK7Le
h9WoDHLO71DYMr9tXhsqdNbdNaWbwxEUuicXpGHN/210mxiKgl6mZ/mJAsoVMZAb
pyqEC/BwjOWe4yYLbvLiyMAdnfepKpgLjqFOmh0HkoK7C9fYCgMMa5mtsje//OVu
XLHA9rN9+jJFbkWWFmCZTNQZguTK3s1F+8EeGUdZtkviW5GrtaZWNjJcSwispHLt
o+STJ2ZJyhedDEVvDEHOS3ho+GUElgP1uQ9KvACk/YSm51r2pazfPUyizvB0arnn
jeFXHqBrDsng3CBxxuKU5S4sDQ/tyodYfwxfadN4zLzmTujYl6dO3MYl8bXXN5j6
xtNcVjrTlopQBgQxN1kBNpRVqJaBs7PDMTGG3+bSf4DhnI93SkQb/xWbkPXxNlot
sEZ9XUT+qvuaUnNtNrIjJmXRH21Qq6WAZPFUo8LwYEplUG+ii53BGDV0KPK5ol/O
behxPIWnikgC4m6MpV/dbT6lpwIQbVGL/SXoGWR9SrGY5s+EWQcmT5Dz08CnuS1H
1tBHCglJ8SkszEyAy4KAgenv5kg/a39SZB/qe3eD7ogINZLmPSWTQE/+sdQwIaAO
ihWFpLYTzOfY3EIsjD8Ih9euixrXiF5TDfJ+XNaVIdE44UKlUTdQPAQeDiNTW4KF
6p8HbmyxIsg+ISqw/nxhygszI7EcRajZ6QXqTFkgod5/F+K5WjeYA3Uh5jOfJsAP
0/F+5/msu+lZFHowRhewgNUooodTTXEmA3Ao8i2w+eyMct7xFqAuiXC9SeJNrxj8
Z0MJ7tsYZvepHVEvreiZ+mKcXvMCBwAQ9OCbwsDIQ9DSLrUSEE0vhh6/pR7RKtk6
ez2avKmnBnlMOZwVMtlkfaEOXVbfVccbsirrprGOfO4EJf4Ouko0d2twe7tNc5UQ
VlWPm73r4UTLRX2nsrKxH7FIzzUpsTdYaKoTHVKc6n8wja9cTqr6XkcQ5Tt036ur
zHRKLh/2IqPoD7zaof//x4Ot99YWdAdOROWbpd0nB52lndEyBtgA280NQixo8/r9
aSkYRQzN5SAENnzZ0phNC7+Wf2ICYlPhBVGU6OI1KF26rhXKS7X5XDEcnByFnoKw
y0nuLDYNceJaceq8tVitIvTZsuZxUQnqkaTKuZ1ooAIEPvUWX2Ebpfc1xjONnNSU
RUu0bMEFY0rRCI5LkIjHhysx0X4wcYODvpw3lZimZYRwEdvqG8hkhVQb89o7IXOu
qxxNQ2m5q3IQwGPCMM3nXg1B3tRg1W7ClT44xyBXau05Iwt6wlSH/G9riLgOwy+j
9GHZX240OqxqkgxDUtTr62gfijkVdm/ap0TgouX3HKIjBGfhPNVwyPsak9nYsjXp
Dw6GhQLOu4rwd3+ty//IMe7AI4D0/y6FJX7H29fRAuOA/P2cGZnoJA80qtCz6R3k
/Ld3Hp2UIVfSLSn2vkPGyxDJV81hBCrz7XA6brtQ6O3xslJQr0xyusg+Y9U90EO0
B2iWVu2UX3kuYBiues0+MfLzfP9WSDDxL40t9s6G9bzt9S4iR4t1Qfqn113IAcha
uUNjjcW6L9wa02iEYYGw9OgiXhEVFsyaQFk/yjo1vO7w4QxLJy2EL46SdL4T0dF3
ixqFmaA6CWa9wbyTeZARCdIgT8I5TzwB7wLD78Cri1ccwWJhnVLfJdjLOwsm01PJ
971jD93XORcnhQhHBWcoyOS7XYfAxdIJ7x0RsIcPgJiJiixrkpglTa8MnFlDL5PB
UpRYi+93OYwnk6yEskf50RN1q3jQsVpC13Dfkm/k+3tWBVE/uCjcX4/u3BDOylJ2
O+CpWjtyWmH9XhSYlaoJKZp2ebYqe41SGPOKQM9mEzwseFZ/TxwI4hfQmSx1Wvgm
y0vnYDU24FCHmUuJ4plbzkph6opKgNdmHvb9Er+LxhN/V8ZmqVk5U1Iju2SmhUr3
3OkAo7BVhIMFaLq0GQGtEUfwcgQxv5ZIc7xZXgs/8lEP/oJ7McqX/NZYuxBSv65D
VmCN1pm5hRtvNHXULlFMJNOaH+FssGQhW69AjsiTcL8WCGJKTXgz3sous5M2hf9I
JbUAWuiVen7eMKDpzC4QTjnTgazbevXuaDmae4Ck8owH+r56KCPv/LlWJFEEiXf1
tRhnGTWcOwzbMdepACZ3FHtqaguorF9xMLPcA2LHWsZswhdnYlHURPcoSZbVfmp6
Jg3yzZdxLN4bT3wRa6RjTmBW7qQQcJf5GokypKEzIkRXIHcdgh0RDyRZy4mU9bxL
IpiR0VYiTKIHMIrX6i4QGs0yrdv1pIEyov9nbBzc4jU1k+bq24t8Cr55QRjmJpFT
fxZ7eFMx6QWSYZGmTbrWJAeyr3dzzlNPbMEmyQkEflN5jY668M4UFLp2VSHnl7Wl
hyIIT0Kv24aNZQmN8c4XBBzVIWqndRN+K7jy8MclY+/CzWqCmjqjxOhJd5CG0N11
kOvMJDy9Vg/F8H3WDhLsDHZK8Mzkj/b191qO1LHCnxNKgvpGfZnTVMgka/jeSBPJ
IhI6Cv7Kxpxmdr5I21oUiOhtwHC6+rp0Np9VIg/ugZY916IbLCqddaf5x8jfwJ53
lwcxkvTXr0L93Nty/S9FAXCy6n4h8N5hlp5mCPcczsebVObi2ri4/9O0TJDymhwT
eBv7TYbmDhrtJHycYK6rzBYoOquUEs3nSqrzc2hhyvQArxFV+G15cDNz6WXkqIhQ
0dHkryhAxRQUOS6J82DGRJ5XS02ZLPaosTQXjCejM55OPCSOEpHVdRBsA8tmDUUR
z07ikO7QlOzfEfXZzp2Hp0yLBcJN+LReXe4VRNCISylqJvn59vwy8odpVLxz6+cZ
LuVVBBvpMHBD3Lc23Izop3xPX2BhxyjjLQ+c07upTT7fqJ3PdiLyof5dFEUQMygh
dDsFiU3mk3yQhcHX3sJ0W+9DilyM63MHjlYHyQnSHZo167AtWKzcYWW1SkFM8Oas
lmzugF1We2GuUMefh7kCZTesLePJmuzMwwceqatoDS3xHPLx+H3BDwVNVq1rAzlQ
2wat8QtzG52r8kz9lTyXc0VOriMoWMdcojQKlUviRPM5pmlQlRM2ExpwBE/xQsUY
z7BGHcrgxp71lCDZ0XyuzRYytvkcuaMIU3Lf/wZ/T+Wfk5Ia57OL+yvPOi11grHD
/xRb//lShwVBnx1yfVwKSsEhi485c3VXxv20e5+qKeIG+lqbsGOwQUSvoLn2Tk9w
uM7+pQbR+Ot/3x1w11crZyGyxBrMfUjJsDi6l4uoIalTza22zP+k7UybnZlBNSo9
6rhjbj5j/1Pk70fAzJZzQ0o1bzrkRp4cbqCudKGCUZY/PLfNj231xpPQvYIi9KBU
+UZc55kjZ1LEgOmkiGeF0JwBxnylF8rHKy0VVOXPylwUuAP9TOxt/VSTtZpqsPNr
c0ijUrQOufXgMHKLn1luPBN1kZvFwZJS0/UdYH2aRJoS86szk52ZyDLQ2AA+oMKF
JP/M1dwUpdU1Z0wIR928hSSA1ObpLEw8aC2TPVVFi64NrYPFljg06NzhKqyRzHUs
YkIQ3ysFb/snGZRLKIktdOOaO46py08gkVLLhWZsDLIec0DywfEjf9dw4dVNDsMd
y3CpBvtNDG08gIWqfCSfuzvpsfBfgT7QdEcm/YBkcZwyf4wHs5on1KY42VXgukSW
h7qbrQEoh85CwI0jMJdbwN+6vGvcQv9TYGOR3TBhhRtWkyZjT+y2C+M/CHNY5QrJ
JjzoF5rBmzrTRdk2q91lpOSWx7QEq0lAULNmbH7Vc0cjBpVy+P22ejH+SSw+723v
K6CdruKMyR4c2GcKSjmkrAmokdIG2xXVYJ8WafrgG6NqR4wgqR07xTx8XqCD46mY
y60ie+hx2d2E8aR63ATxbt8zunxq7b7rk02Sz+weMA7tf2neQ/YG21LRBWeqaLLV
19n9vof7Wa5dyzQTSgO6dBx/FlQ7OCs3S+UKTNIDKTQr1tAuE3orKUNHQ4RuowQv
58d4mquO9bZkcuIREom2RCJvgOzEu2zFlMvIOTYIskv/CSJVehsQhoKO7giw5sDf
e6OF+dK2gLrFA/WSYvi5lXj/rrFLNLDQoWbxXxSWD36HXgtShdbiCqS9JGmOoIsQ
TApUhGhhivNn9hJ3jk7u1TUF8eXeEJgVbALFAS2aGK1jlelDvFkgxIuve1GRY8Bf
QIABSOqdxhI/jtbehXMuaFHDi+HNwTVcggGPsB9xRwncW+U+G/ZKEh2X2z1Lkjth
RVDP2E5kyRN0HYkRaKx0W2Lfz4jQC40UhUcNCLdN/aabXesLc/r99QRKyx8QAjaz
cpzB2WysK7NMGFNg1s+R4TwRhhv8xTPj9ZXQQeaXWqGFvR+ZK/VIB6Nb24Y0mGFM
3srkG+3N2tA8f5GlGPQN1TVa81hGFdvyK6AiYnRdk5xZcCW5edc/vQ59PmhrOz/W
aN8WonYhXRgUFCcTVUBXmGBR8ixFkH/CXlsC/0fW5IudIMFBS5mggDgRj1tu52u3
b0Rtm+Nxj0eIr2KXpjw4p14whc1CI04EVSeit/yzMbW/uJwH7EmxXg6DlHFLQBBM
Kz7YCP1tPDbkfAx0aa3fSW/rZVSUrFkYb4hCNjqkQwTvj9W4Rz8bniYvpOwoCNPX
Vl+Eko2eFGrN59/qyy8p6nsNlrJcu5mWpdbrwY5YKN9tCEwG+dxs4yND4+Eo6o2V
/wlEaIVtN1asF+mIr9V/1b4ZGDCJyxpFknoZEBgvUUW/ZPuMngOrSgc1JW/3yMLX
3bPtPjXB05yH0FFHGStGqlYXkpZB4BtIu48caJ/7T+wN8+yI8mw95GL3MG3EexDW
ug2bB5DZzSzk9EmiOZ6/9tr9Wl2ZJKDd3I3dbJjUxbC9dScBKWmDdR+EVVVINjOS
y2Gl78GGmadtGBpEcyyQq9X3rkNE2onQ+abghw3ZofyvCYLfCP7mR6+Jhsl0lH39
rIIrb3Osjgqf84Hw2V181vKbvhDGFeMK3GhaiYtD6HG0UJBHEvEIwNgtm+MmCyOL
twB8O4/0YRGLmP8Yke5FvTCReV/hySnV7UJKU+KqCFIcxbwS5jr/GlJ+llDsT4Nu
932SHy8jFp79iqgaLrGqECtEOLLnMjXFD/mvUmYRZ75ngQkYFUu0WfvAnayWIOoI
evQ6kAStho95SFV2ru1K6048qKE5kbBW3cdyIEFQJO1bTm/oWr5ouhMq9CdETr3y
fQ+X0Vs9CyBMA+tnTpj8Z6kiUbALFld+/ibLJZEyinFjryvYDprVeqZ4WLUn5GW6
IzkLewOBXpMyDD/U4bfJEgx7gegdGshpu0TZh+suepdMtEilFGODAMY+f7xZ5Wuo
wqhnUPw2stXg5XyyZr+WPAsnwSIXzI+iSOTznis+HBWl7lzsWrnVyPdNV6NvPIT9
NNqT2hzmSwgoaevd20ZfljqlRQ6FZ+cY91PQV9FkbZLeYlWlhtZyld+5yKnLdF8m
STfpTDGWiS3Te1Uvbnm8G5o+r3SwTdOeh3qMhiHx9rmach5//pGZvXF9dLYD4Mw6
SV1SvtYy6QyLhZbuN+cbgOu/bsODmLhhIIfk99JRfduOwu+Rj6vSJ61IyTmSkN60
q68dIM8AqElKxanLmZY/405PV2J5gDH3dcWtWgGbZ+MhE03tcyUOV1z7VHsbXG1W
trVpyNoP9epjbSK5K+HQrvcPVELWyMs6szXFp/b92n4eidv65nvcaMWIZ1Vro4fw
seH1gFsUBvSJ4Wlid+xhwCXBqJgW02nXodO3zW2dQUVsA3yo5bqhkGp1qaaSrvkI
QNObsZfXI1btL2Hpqkx61ItpkbbxKriNAnXLStJHM9/X/ktTNxH2aUPYpD5DjXKU
1lxvpAuLwp4YhuvO5DLPfFGSXQ8UGQbMfS5g2naycZ6iXRJYapLXC5T3xC5GRlDT
A+SZVydBQb8wl/CD64CypABdype24CHYUt7BGzzxylEIVczvCGwcamRWYzxtZzbi
zpTikwJCu73oXJ7uve6KwGAa+IaV0nsh0WzKOhuzd3RSwNeGoFB4i17Wtk/Z5n20
QgYEJ4FTYthva9zNQGtDzCiEILwEEQPWpgq2szp5f6Sn5iMX9UUSGs7/AqtOoA6m
NFyysCr7V5vRwBVrQdAqI9y4CGOT12MiZ2goknI1UD7AsXuIAtsJWT7HDcQIdjC2
VFxLHu5tP1Vuq/5Ef/74XWn2ZNsw13Vl6Sw2OvSp0++vHA56SiQ7WU+ppnpn2t9L
c03zehsTdZb+VFEvu7ilNRscU179Ak3GCxtgy9QzuMpdyWpoCsuNMuAOMhPCplcK
15GQSpOggzjXoql1GW1h5i+icp2ROc8SI7XP6xbECWJ01s3WyOeDX3+vf5VJTrFP
y/C8tf1CGJ/PTSorzDjdykgq5EDrIviNVqBy0JEGrGMzei5D7ubMBs0CMjv0asFS
qrVBIciSK+k61Rg6AzYt7Nmakyl4LSfW2VOHRvhe5AyCKO22bMyagy9IzmNYEl1P
CrHGQ/gmQRWfR6BBh2iMpnlw9VfNQWr34eftn8mGFF+QN0NDd761oI0Ywil4w7Ic
VgYizVTNMWY8ghwAnFoIX2fEZd3yNQghnXpnW6774xCaYCDrG+45oHGn+Lbsn7oD
6XAYLnksfRSiYjTy9Xt+iEX/j72lAx4NEoXvQ3eQv0c8AoVz+u1ZrLeZuPccuhD/
ONsA2nJGINUjYjQ8dHIBkwMSy399hDhBbB+Pr5h9lX+OoiZolpLssJX1o4a0RcQz
PjD8XNOIxlMDJ1KvHPCzyhvKhknE3TFrsGYIS9lz1gaWDOK3HVXt+ecr2Gn1aA8v
odnbToDQN/aXDXgopQD+oBkiol9TsVXO9DKLAfKl0uD9e6C8mivZFE7lyhwjbVqt
7/gQasQP1CZuS95Q+MawA1EQ7QlrG6zXTWxm3DQd6XSVtWd7lsOtsLadzai1OrTA
B1pK6NwhUsuuIhFZPZnlSgIrEQO3ewVJn+nS3l/aJrBnaZOJy3UVc6M+3ph6zcZG
sSuQXJCqeBWS8Drxvo1yVwVSZL8dSIp3I2bTVdRD7gvffYoIb8aAmCtP5B/PEqkF
mgl0TxobLluxo5kG89lO1kSS6P5lo3cy+AGX6hkCcCie5AtzTfpqVs4D7nLpsFvj
CXkqEGfXm5+D3VWcyxju504UW4ch+6Ko+dgux0KcVam08uKY8s4ENCbfl/hByQX/
8qyG3XaoDU/I7/eqGZGVc+RSHQH8UM7UWB4B45EQQg8kXhJSb4ViWNuJxiw2l2ud
/GbKQhrK0Y7a0+j1irqASCq9SimyudQVigBSWPUCti5c0pm1Bl6RRXCwiLpMpPY9
+SVR0Ea2qSx3syMhpdm1e/X1FqwFO9TqKLdoQWQKrtt2dze2chjdO8O0R9hVM3l0
fDz0C7qdoM2bRuXLgUn98Fr1Ivw/gqqZhbgZxx7q3p1UcLBJWERYD1sBoGIOiBho
C8M6yz40ix8n7yZ2AoGESUtHFJw0JmbT4Wwtd67BWUWQ2qnyh0hEL00gFsnQqEa2
gHmfJ3KIVGWgTYhcReEG8kFm5xNwMqGTLZDZDCENthCpRZ5TtSn8C4qHLPs4ll3n
mpXwb1tQ3T/8x1OWbb4aoRBBuuvamZNE7Y5rULX0tbxB5BP8BQ/ZZF5wUp54y+/d
O/m9JXT+OHomZTQqT7Rz6zDcaLxlNHsGSiIkA0J0mfAn3EJucgGvc2VNscKeDhNO
Qi+ocXStwNHI3sSRMUTzkplgkhUbSAc9hLcGwUnt5e7sqMtOqKIcxXICcNxEYNeV
+d0gF1ZXzbbfzdSbOyZoFRt4TQeB9ufhcft8Bxm0aKMgoM5jn5tvTXq6EHI5NGOe
jEc0Wu4gd/MAa4Ug58wgmLnaz0b6FX/3LjtH6RnGvPN8OJReC8tu7zNpuTd1O11T
brHuUgXX6uPZptgAi6+phVciCZBWPTE6x/tAq7fb4cpOv/dPuHQDTlFAGhhkQBxk
rjvL7H0u2fsfganiX9TWI9+vq0o32tJw8MPMk1ycgalxYm540AvYgW5Mv/kJJksp
eFmWmiS8I9WN+D275wKKpBmPjcqRhiAh9M0EegD7kIN8xHzJ0kTgDxGjXudi0x8Z
/9k+1jstRVOCriLFxR6rBf/x8+aifmnzP0bhXJHyQS46msdPWBPf2udvCUuh/tqz
lffM3k3Fe9XNj8l6Ncu/yNDuVEWFDNxcYgSE76hrOQf6TPw9SYu2dUHaplyLMKJE
z77CiFk48gLZbf+Qhxmjp4PprEapuwJLNPxoAx7o1ZXT8XbuTUbfv+UZv4aCpu+F
FVyfgEvTxl70iZ4fqLi6N5kMe0ovthBgeUGjj+oEmEKSjFY7b7/eH3Zu7JVJ5M6k
F5TUsSY5LFW2Mjbv+zg1CSnknAl1wz/CEBzIbLEW6L5cwZIX3D81qnkYQvuXGs6v
qqy2wVJpTGrdyrV6u4RSKrB1F0plQR5Z3OBhq54iC7wf/+jiBYHN15bx4nO89xsn
MAdH8uylDfkUyK9+n8Xxum8AtRUn6nexMh2xH786dbOirZLAFcR/f0/XR30ujrDZ
EzbCtkVLQ+1mTaWE7sSKVhxcrX697+VoSBTbq6q5JAIZkzyte4KTzG+xkoI2GL1z
KpCnmgiuPFhaFvcboipk1kspQYv+UIi2DL8fO5IMBG8nbUMu+1yqrIu6aITcV9Yc
pS1J8+i6oi5RvpGCUWtfdzqipguWnsWyvkEsnwSBZpGY7Wh3LjXYlbDJ7aX1wOu1
eXlllBiZqDKbbcZfmBa8hZdN2I/E+SWtN5xbpvBIdn3VIILjsm/mgGcNT2AAwQC4
2dtdznY/vWQ5G6DgLxfPzH3RVyeh/xejdE8n3xMMFMzrqYrftcUZVN8hIp6hcEND
AX1ccYpmZNOqYQADAIffDsbF4qnQGnuGPfG4p4FUnkz61KEBuBdvQuRKSy09rMBl
b9RzbYLMQ/vVYdtHqjVl76E4bFOcX665wY4UzLJzc1itBYBWu3r23UTFWa3Rvz+R
2CizuwyVLXOhBDsuU+bgPaoMfEnBjzp2qFXDQXw8tzAH1LN3xr90N8VYMNGk3yiq
pGDtf8se/x9RXQMTREQsoUR0bPRJsHHzLMfji7UTSf5Y1dIWkwI3E7mzi4M5h5QO
Etn0OKvD25cdjUeHoRKBKhLapkzdIEl7OrlIBuQnnIELBE8QgH+W69n75uzm8NAj
cX8Cs3pmTezVPvq9l0+NoXx4RRmCnjYj7RwYccCboAlvcCCkdizg/EWI4OuyJf4K
pwF6PWfIpCTqGuND2pKkifNu3KqS1IEJAQiT6hTxQCRtNiWVfzjw+XU2t9fPqVCV
Va/keYIXOCdvvl0CBMGzI5wk4NLOWi1tdznF7VMjqzuk6yAab68rqBpEY5NzOvsn
AazG82nb9oCXOFx7NemEJvpfwZDEUVG5OSdlhhRr+f+/c3it6dbpRfkPfz3JNUxP
uhrYHUWF0s1R6jgpeAYTG2l5iWKBgHOmzUZICpb+a4uRd7ZKpkh96JlWi1I6HwWb
0owJ8W1B7ylpbDafsDYylTpXf+U6Fnn17L6vL+8ox0Jhwg4pysdL7q0ObjrrRlm3
z+OYzXTPItAJHjJI8eJso93jw3cIYw0XH4AKUvSipFXwsk2gixxsgSb8cHEW7Ozk
s8QK2YEsrBpvXzrZp7/nbypzEQ6t1hj0Zb/WCBalwZrTE7/jb8k57Ppe8yJ5JDVQ
C2+w8NoyVz1gjLVoq40BQaD6lZXU9VRTWcITSL99D33thDVToPmUhwcXGyEI2LaX
3l0VWqMCjBI+5m2zAEShkfsB2LR/jfKKAfDJNTjHOvofgQS9tDZmo5qbjdWsbO7r
0mD7WV/HtHxRYfpH/U0AznqdrRdGqFiS++oiRGvha2P5GIK1SzxMhBzcJJs+b4Bs
Mc0yEB9cmFr1RHILNXSyI+4H6IpsDcHxzx2MvfZiNVr6ltuVK5rGD+nzRzw9h+3G
vFUrcgvOeKoCsM13Ldxhuq0gN9doRP7rRQ3kbea14aO0xcTfmocmGZoTz9Sf/VnF
HfpO+FNIauGPVDEoiFsNL8lKUPEPNp86ValuVnPMZdBNC+9eJESE1QXVsOrOA+Vt
bDOtJ/Fp4jDuL7o/dn5hDAfMfIkko4fpSlw5GL8/2F0S/EA15vYo0EZNHZp+xKBX
A1p2CBxY30zPMaM3u8Hc9pyMi2yx1gWcSyZ5t88t4UUzbkWPjKgFqq91v8ifsTHm
J4MlsP27cHQOpwVR230Lj3H+RTUAJfVMSJxd7c90wUNtvm91hymuhCw2kqnfulF3
U2hz1NWy0O4B5GL8teOnOhCzkg4rhdvGw2nRSasEr02Ssa0LdZ0Umj4iIkrnxVjG
yXC5DC/RusEdRvk8J1kpwUXoUjH0sq+Fq+fryNe4SRPErorKPgCjysmDIXKuGEvM
CDLdesWOxv4CQQtEM81v1VqV5oOJEs6PvnEi1duWq19eJng0TKb+GDcovo858IFG
N2Q5qNX1RDk15r4jlLA0/KmkhszS2tIHIE3/ris4olRvp8UPpMSuX7cCrdREeCn/
xw+UYbXMof3EIK5l9Vz9PpKzOKA6bObxeGpvAbVVuH/Of517dOnF8gezXJEDxUXm
WQy+YJra4W1HJ2EACnWiBcXfR8ZPrnyCvNFc2uskCh7Bm+tt2I0KatPUk+xajO4F
xyJfl56FsOuC9x845EbUSGR9kAmq1BRlgENtKecsutVNdf9jRAztttAEPlIW+mQj
gTr3uiyURfhlC/NRMc/6nxGqovsa4X/WbDjzqZ0BcYzvk+al3odkhq7pvbF+waAu
peViWwr7UG06MAfzwZ2Mb4+wmmzq0/PAi4YNGumY2nw5No9Wru412XyGCBrOHS+4
fxuDmpeLbBNru0lSMogqOf3Do1/ELcjfBB0/45ABFH/nmNSyI35PPkX7H09ukstK
FaNYO5U1783fnZRgLnXD1osRVzxxquIoQ4iufhNccQm4CcadNSYkvx/WOGs/bC+v
Exa+CWWi6vpaPR5u2HKCVO4f5EWozdkTH5jyvQPNroMBdIUUQI3B/QTYUmhuWAoz
hpF+XGxH/I0oJhWVGkSyoCC6bpgwGVnz1itCIDcYDDegRXVOu/tvObFy9bs3toKJ
nJcdFmREeKkm7HaEhcb1B72tht2lzWxVi79VJuiXNMp79wV7UkRCGpQJqbNfU7F5
vTsk951/dgwBsLc5SDpqGp52Ej8ZAofAE8SLpPRIYHxwlyVhmJtFpi8VDFBTgFDw
vla7rpxSdB/F4uyqky/PnA+az5Uy/uU52CdeBG55pht+uQH2D3SOLLf3csR4TMWJ
+vv3y1tTYFJeydzDfuGbo2iPTN2kJXEOeZ0ZLEmWu+bB0z/gCWWxnUvcSqdzmwJc
L+gaked+KkVaLr+04CpJw+nst0oX3d0xy+l76+535lqKeTQXscvRj/ZasSWdiP1C
Nq7oHQRxDI9PCn8LU2FB7/8BjYIK1Bk4U51BNW5BOQQmUfeFEB1uve9BgWN4sNrS
lCXyiN+H7l7mRE7eyDx84tsYJGKCh3fj1+U6ccAQPzbN8UPSpxhcbJEooHKGcxyi
K8OQVyCuyfuolsEg2naY/mMkJkMUKxcN/u2VanP0wTHI6Y3gvbTR39ibS23gyODR
ZROgBDAn8IrwVrOaOl8AY+kPkEVz3XIesXx0f/eQRZic1vcz+7qiofdTLoQsFyDe
7hLBeXvQp5g+8MiB91oqiZPmUgWy8Tbd1BSU1cN2yWegxqMqTe+k8ofdp+X9CM02
Bi/birmQVzMvLnrCPRLCTwnAUiP8XrDMviVUHacXTXlyhate9yJztH7XYhvqaM8a
oQ4fugFXupUCE9pxI21eRWMSSQMPaopGEgEHaI/dsHcn8BB1TUjF4af9bmSIu1Fz
4jCP3MHzTjlvbpZ3E7THHWVlproac54qCdR0MRdZDmIqA28OdyPztIurb5Tdz2cx
zhEpMFjY9uiVaPn7vZGCxnwaYu3FBwFTqlD2LfFYxlrPLFn9hXm04esbcA2qpXNe
9ddm3VS9sqc660dTgHKinjm4KvmIFJ84Ci2ksjpzg3HdTB3z5/v3A2CaZk8jpJf7
TEWT+b9Y+rxsB+Jr6j5vRCST4lZE1CQs2pThhJZNDrr56bhnlbPZdo5nClOamb1H
2mrUGKNZ0NGhB6sHqZEhPNHvkgS09gDTzdNDTpN+B+8LT/pE4rtgUxeiOowxMdop
3+nq7Brq7mEEzl70FjInNB2fjZ9zJBaD2tOd1/iAGVxPes45Nzm0yGRcJGl+03/5
qTgKSjJZfjlZw/ff01MNFU7Em2LFzgKoopqXOUZDXAXXzx9QPVC9GQcC3P/FlmtF
rJRvJcX2Cym6c0v2YhgDq9DvhzNDNmj3w+2permvbQyEaSsYehcXmYAqbPoQkGzl
gdNGKU9O3P3geTA+DTEGMS+VeAsyC9NHaD6O5P2SEemcGy/D2lo+OR8b4qDtZbhg
dlwTzJ7zMSJ5SxyIAA5BeIm7USBtiSICkURMRQJq4sDxkyukbE17nornDdbaj24V
QDw90w6uFMlt1bkyrw/MuDy3rwZMyOk7tzstklN76sqP860aOb/xBHkKC8qhj7e7
Pjv6KIB6VWDXe1S6dspNG5Pj3rfMLcz+kpNX2ijUpSAozCZ/bBZsR/Uaa5afRz8V
zcrvhruwmb62FmNYiYnipV99TG22oirOEPZ0aqtNc2CxI+v3ZUEpNM9DtNV/aU55
yni7k2u/P6injnpOPqtCMYmeo2cZrSPjrP08I29CqmE5a9YjrAGsabNJq8hk60At
SdH/tC9nG71/4Zh5VudqLDneanfeoVtVvaOeSmgfmvwZD4ZFdm9j9xUQrbWRmIr7
ouDorY6oFmHyF3aA+e9j4eH1VadgwZiIPCkm27p0PFjpCg+n2EcYlFQMKEIbs7OS
RMheEYS2m2007IExsXBNoIA9VDeVOnTamEGbnK9za6ZA3oZOck6WBBRRvp9mQaMP
s9tykgUYv3NOrw/KJ5wIz0KsH/cRnq7BQXuKNeediCDwiKJryq79w95Q/ZxO+dnn
11ILPAS/wfDK6aXLSKSAIVFl2K6vq+XS6he2EOU+oXyl5pmvZRhGUQUdmTpk2PF+
5mWKdzwvM/9MsZK6q7CNeEYw/IpUI6/9We9bLh46i5VzJFhc7O9lAsjQvgI9fNwB
XbCusp297v8Ujsk7GZqmDuegPaL3+U28i4x+OQkOrmDwvI0COn4tO09hfYDO4ezy
Yjt88PjEPrf6l1PkSQ7AoLlnBdapJS1GELx9aCzQEvTsY3KOXRqdWDo/351rwKDv
ZXsnsSeoO0/NPb8dOz/AcWYPsocmC8NalIzUSFFJDgTql+hoJtHC63G8O+Lp7ef/
QIziY9Q46jv8BRfnpIBDqmJc1sKe2lc4YbCe6b8wadyFI8BVSsUOIEajYApUTKop
Jz+90Lj7ZibVdhiaoBzxiSdGDs0ChU5ii6s0ai78yF5mrU2qp5K87wl6jG9Q3Mln
lA3WgLuYAYulTWOW6vihM8Fwy4K1mrHoCGyX/P4cskkT7k16J+q7hDMJnQV9KdMg
heZdaV46Gp9Pm5Wo7RecES9VfzLvFRk+4TC8OvrXKdmCK+4a3PjB2Swg56DwVrEz
Od9yd46MkQqRZG9racX4qCHzThP2ELa+uUk2dasFOkxHeS+q81cRDV2IWOVr8C9b
Oa5eNqbnp5yGdrNl05dcMeXotItSel5WsFhYEnIx1+gznZslaWiZlkmlnHkB8otk
J1SmJANLbrL5uycvwjtxT3udClyTZx9atGX9aJ0ELV5MK1cKh8FoWmZEHjCJYoC4
5UHOa68jNMz/LKEx69mX1pKl7yzagNsvCouUOsBta7d2EL8wxP+z2R0mNBw6DZ11
9rNAEYA/6Odbql086l2Aw1j5q3Q7VIWGzxBFUeHPR9VtdR2EKt7jjp0gGI/4Zn+6
QOPbUvrhzEW6Xd1u1bBGd7lYD1JttlBaTHgm2PdxZXAkJeFsv/nVlzR72QrpdiH/
H71vlc7J4uBGZJANfOanRJFnjLzTdR0Qu3KnS3wjVa+ciWAR5Ln4eCwySxUlbpZg
34FOUBddx4RwXlUfhBRvqzNzVwlpzoomcWPARGTbGi6REUwfcdFJZ5JVGHaupQ1I
dl4JNrLr0KW9NS8cv160t8+iuJgl4qEfjoQ9nH2USpZgCFwehsdmq4OW9qrJDYOx
czkZ9fWVoms2HhLFKR/msU/14V1s5b3WsP1hxLQSlocl9cMqsYhPRWoriYbVYSlc
KZXRqWtcDf35uHLbg1JGNfKy9xd84+u5ZitCS8xpZxOP93O0q6Q++T1li1F42s4k
DoDaNDIG/YHVUlkEkO85iIbomkQ7aTsRhBxOOvjvi080UUm0/Y69XdYvuVufkDaK
4TEjJfkVMIjJqNL2/PyM9oYsamkclCGKjllM7tNbu1y5xuBWDcIN6R8R9rKQLmU6
a9EGDmjUO6blxZqfrSu2LzMxLsREixRXbZpIEXPqI/Lssbq5u2r/zZXmkM/SP05t
HOpz8AqhxHijXIY7tND1tD/0AjYzRFuVfNXdYqbUMMSzOI9k18sTiti87+lc1q+r
QoI+FGnvYHwSqVcMSUl+oAxsNH6GCUWE/G1lNtoAQ5P8K99xAl+/hCtSZkyMQta4
GVjPshKzYlQ3UCPla4QTuGCuIfpzM1kqaVxMXC7LWhWAjeCYCwVYKrW9YYOnDIX5
U9SCtXLgkpdvRWcf6DHOZfeXUkEzdd59102eCDKK2c2Lm54Er8GnRv39HOgNiNbb
ZU0mBsR5Ql6NzXJgOKW4bq9yoTGV1bJ61TeTxPQAOiflNOO4SmzsfVWUQyha7FdR
VzNoKZGKt7le0v3JQut5pkT/zlMlZ7z55WJh8shkMS78Z8os4r0Mp7Drq/2cM7Zm
S0/wGjFTS1DI4CxjI2/apbxDqksxuVVfPqoOChoHMzfcVjIXvU2iDhR+LdWC+1ha
FiIqvIkJ3YSCmpZJLgBheDN9dXO1oN99gn0gJkU11Tmt6xtwhQ+bwjwKz/Cy9Pky
0PQHIFyBSjQmY8qGKgZsXQxGtyeJL+PlqBffVCKBsW60o+i6GYRusNsdhZk8GTs5
xWrcrkgMlmF9ZyW9Lao53zSXeAlS4CcWbyFdFgZySS1hq1JfukROdl0u8+TEjLcT
TW4l4x18irK9uIQMTZCNhZaSGPWsqiAIijZE+neVlEIkwVWDREagqCw7GH9MOPLx
wG9+I5ohGYL0IV+5ysrzfl93NNdFtjpC0Jk9QSpFiZoiSgkFdzXaYaCVUGR396Jg
JxbCrL5rF0XiI+5zZm/ZzfZMh3QVZLHMcjH+Jv7gSEylyg2p6TPYu3CrpgAu68q0
EBfcQiVmMsItw8pWEcFbk7o0zqUvkeJRZBu9AldZ/Wh0cvpaXNhfI2PCklFpBqQC
7l0qjVCXltDrm6fKBmW+s7IfYjqkGo27N42epHv8+dcq/0pSQNzhijkzCUnFMV48
OS0g+64OvgLHBicAsp06KIjitJHoetpxvRsm+x29JueGDeW8lr7UiD67ftknNyO/
WOYVuQ0TKcEvC7nmkFIeGBOlqbYGUqSzyxQHOxxzfM5fJM+Jlmrq6rUHuSm24bMM
Ybx5uW6EeyyIwAtJ8UhuuqhjjhfIq8ce8fSY404h82h4PU83Ovf/LX9ix4cGr7/N
1fD6RpXhK/ulKlYBDbo7wqJHnmdeG2T47Z6OZR74sKjcp/nzTGIzotmMX+NXpoBQ
RVCZcMhVH/HM+sTN09nWRqYVldq6JNKMTpcS3G+BjXpuKJnX+9VON4P0RGBVoFUu
1mGx8FA7ZIq/FFjwvBLJJD+ppTLiySNAK0jdv0JyeRSgTuI6vay2dkeJfZ64Sghw
N2sfU7AnY9Kn6upipWKmH1skoFJO6fUdKmAtdnbeZECvKz1CNz7OCltHln4sAtj7
seVsR1PpgLnB5i13UTD8K8Cj6f05ZCOMPMOSdL6eyKQCahvqi3poeo8G8NdQt6oX
+l5ct5eYrh5r4Bq2SpRfzcodaSuVr9QJuNgz4EOONDhLEe7bppAVjKoWI5oeBmoc
2FT9P/RGOaWFn0Qf9KzDQLaXKQeZsQxZM0MBT8tncOwTmEMVjhpcWub8YMdVVR34
x8OEj4syvcxnqQPs4HVYziHcNuVZb7Q26sj3Kp3J3o4tHJCnDMDm7+ua4PNzJlVQ
mAk8O+ij7MuOKpHPooVrlx05oAqAEvxU3zvnzvlZr6JMeoazrXDo5JJudKIJxFqA
6TeoPAQxL8Jr0lP91OoPj6q98hJe1DpbkbnQTnTAcCSYcgj7bW4NcDgTQ4pfXuIx
xp/lU9/YbAPKhhuw7itUf8xMA3NXASSzYruEknyx9fzXKyip7UxQS1IkLes2aEnj
qAbRl3FbchqQOck64KaN5zTaoxruo9iHvO5l3ecPonmh1nByk8ObDUw8ahn0mR9y
otI1JIEjAMc6XIMr0iREWYQ1NQ/4H4+xARjgjquw/resJPFTrb4dCPUp6sedm+VJ
R8MCXGSmGxhSKCWJyN7p/8LIsjAFLPs11XH07bjnIfkd3HNc45r3g80Qg7VCOOMB
5biZfgNbtSuMjYLZO5a6n9bkV+PHFusOnx7Azr+ga0Gu12O2DHUPGCdppicn4wpq
1wzHxJO1RQz35RX9RPjMkv+5cEQYav/vGpx/6RMP/DcguGHnfNlMeaMezttQg/iO
mMHJpi/mIvJiZ/ffN4s2R1uTD0HIdRoQ9r2B5Z5Caqxpz/+DgO7Fo+wsvvevQy6j
NQ9mtPaNnWqXxxliotb9cZw8LS6cqJQM5nZs2sDzFyAb8FTfwB4QWaIMutUZ/dnh
fs85tOSRxLTqZcHDg1HPsuJsQQdInFvUnaE2jBoAnR4IpnYlDywQcIKWtcmArjGc
PxC42o34IhvFL7otAcwkKpgu6ZW/d+yH1KylMgfUVS6FCtQNrp2/HagPjAvWXrjc
OXYpw46pHvFUTlU6iYzyA3sDGd8dC+Kq0FAEfvIXpmnV0nVM6qp2BN8F2mblQu3Y
6HUlQb11y7I+JxdeeywUHd10oGazM0B/ozOSQDEILjCaCHgeFlDgj/ZBVVF4PQb2
Pwu1xwzvDpkyz7vzz09Q58ufDxruU+3IyFDEbbYtEl7pxrL4YMIo+NAbMVhxbUmu
WS6n6v/dGC894cyMMabTT+vMxb3UGgPLRIgn4bLkae7xfykf/TdpMCgfS6NfXJdZ
URr+g4y11O/ir+WJNsOmzliZc1AqOdsZkq/4QS/tOnGDJYjLtO4NzjZJkAlNKIsu
EHTmK2m2LVUUNmoO+4RQT0NFEAKnLltoQQtp6uOkUcg2CXRAz5j0rTMzT5njFf/D
htXQKMx0WzwKgtZSL2iMkzJ2FseuBCBrFVFPl2OTlEFdoUaNh1c+cw+3AsO9dtwj
8LGzDeKGTxupE7mmeHc7Vq0bwB7GM5J7AKl2TrafZcLKwYtqmFKEECtjMozfe2EX
J/+rWojFdOtMWah3NAqJ2GATTCsGGqpyzKHa/On2AsCsfhM8IhEFQkaINMSciRdZ
oWXLOMq4q0jX7IsuedQYNUxqb4GxMT7UPcsPowsh7X6mTOUE3x7CMY/bp159CgRz
kGgIxvsheVRUjn2iCGk1Fp1jgGHhtUeydxNxGW7qzlpOxwX63V2q7nVXh4PKabYR
1pZEh9VOIZLi2BfMjbrWCmdY59ghWnqBQk4g92EF97zkiZXWw2lSodS+O0Bz284J
7PGA08hecKKsdkrLdJz9GYq9Y7RVFxEKfzhbDHOyO21HcnAD4dFpaXoDvFnWQ9mL
BzH1fFP03l8gby7iq8AczMF83T25Bt0G6tW2eT1bNUgjH+DdOxlz2byVwMTQfPyo
q/7o8hhiTu1MUdgVMa22V5LF9+GPA0ddYONp/R5jmNc+4eWAiFdBYTQNx3erQshN
f4Zt32pLq59z/wa0GSjFtYoLl1Ap79RLOP1HD2FM1cj4R6u3786LWeu4PjxY8cvr
13AstJp6hKrvq1ziTeffxmkb81PVvSDxBCrrOpkxaWMo0zCXpijLYUKGjusT7L71
rFADA90Ojy4g81/VkGLCd6zevj1lvDp3dhPJKK9sKf09pr6Nc6aw88vJ7xzcoovC
CNQjngVpz4bLinLYo3syJOS955O4nytRWmf5rD2ug73vTtGIZZzFBvbldsLGJMrI
+0HtAHzFoRFGa7hfZHB+4+Qncj3s/ga28J3+QpJktrVmOKM3mutvP+R49a3QfpWW
zcSavlKcXI3mhdwZV9Zw8M7g7G46Cu6hYJZV+Q4XzITpzjPpCOtvZiCw/7ETpmiu
w0MCD9iArhcRYL8+nTkcAAM5RI0SHYDzURMklICXCL+0r635i3pJ9Bdv1oiUQCPP
nKPgi9SbJoJCc63jSYln2oopX5k760tVo4X/0x+ugFvAPbBvwEySI7bJFv9jvez/
tjlJaSWGCAXJfa+y+eXGyuFEiIrQhQb1c5VE048j5xd6zmhm5Vhl+IeILAdrRMUJ
3AndA0WA4LS7LT8+OnB2dor/OoZDezAPrpdlCY+I72xGqEoD35xL3wwEaWPM9bki
oC3uilXRj+7MoG/MH3VtqMg0IT/pByf8z7ZV9pRoag5QwkLGfZaTi9zWbUMq7AfN
9rdOV74OatrWOv3c/9L+r2T8UtvmgcNiV6V9PEusH657xaZe7mNYtU8PqSB2g7i4
y1GI5ys7dCCMVGgDv4pPkVj7ShS1ZtbYFtw3TueogJ6y35kv8aQ6ctubfB7yvUD5
2AkbLL6GIj/OQexHSOFrIuU9ra4n36z3A4vrRnBV1GPLF6EQRHBniEDBXaF67Zr1
090dRjVIzMR4SgWwYGSK3m+Kleb+Eok8sR3R0zhs+x5vsj6ka4UkeWCvaXAb878l
MPRTkRKNnVI+Mh94mO374a0Grbh8JNnC25KCC+27rJ7wwXRivLcdXimGmbl4Zi82
Hl7TgjSCKjetc6j5lJUKe/+5azOpXpjfNjy5K7y9PjRroppQDHFeF+ZNqENCfuBd
acR9GtYnLo/dsDrT00vYV1Cq413JaKp5kZopa8hgKWc3DBjCb2+lrAcKK4Y7vDT6
7KOG91UYU8/BeSG9GKdOlBQtpVo+y5A0PanPlyAFzj7QBiWzeAQVBsE7PrxRzj/f
UGdZuahaYtA+7wzRi6x88EhONvawF6wUsOuX+grwY+VQrt3VfTRZjneeYDoHkWNz
it+sSSnY9qG+CCgiUV48c13ZUTozjqqP0gs5paTbm4nuVIWKOPJbZOmUnxDkJGbL
dXPmeKMwV8jKkhOGM9O8tp5pJ0iHC3Y/qWFE6K8oJdvAb6GrMLtGjwYHxQBXoMnr
vLwwiBZo0uJQCsincumnSTp71z8LG9qvMHyO7AbrRInA2hKV99iATLJix2+fLkt0
W4Eov/1/+v39vFZA5XCLG4s7vxD9KGvOIUbWYNWy6Dv9aWqcgpbxKTsD1gBwzSHZ
qX36SiWgW8FEuxsyyvwPRFa/RnanbhSdUjQmXZKUw5YohbjMMMWqONaRo84TNHPu
hJENXZeOmLpXru2IL9ceyBzBnXtHy8bYf2ni0tPd1FYo1PmD8+S4YIETF4LsfUNq
YCzeYgLv8RIPaVgdvHsG0biP9xDZzOVZH83YxZLeqnDgj2q1bTKWg2YVzUO7yuVJ
boIKS1W1WXoHGIj/w10/bAerrDHSzVTbxIHxhCdNbnbVrLXRx1yJhHgGGhYs/cnG
6dYDo3rzP6T06qpbtZ7cZDS2L4kqOfK7vBjIPBKKPmOrB71SP+IEC5dfqu7rvgSa
0O2liEGIqhKH2rHkTznfmKoWfKYs8/waVmINPKkk/FdfimlyQTy+hpBHUAKgKyjZ
2b2ie8YQs2V0KPxK5xMvd6ptYM7kJ+xvlqNeREQNsx8YIn6fmHWivgBw1pdNV+jo
09sdSh9lGkcyb/2mG/ldkeexz2MjvIWyMw7lzDEYS+tAWPCRcK4tpngdrsrSP8ni
0JjJNlBXFVsb7w7TJCxK14fEwuJJh88Rm1cytt0Rd6+8LZl3O7WsGIOvUBldpU5T
tb/9xrFiHxshzokwp5yS2D+qpI7O0qRMghNyulIBPIuiWuALxvcS5WZJ0ZYWfL5I
eb7L7ayTbeIF/st0depXmxbr/EBc0OYKZEQndCEuSjmG8GMvXBKoxsCsFliHODFp
FW7MPwkWSFD1U54Jd7ZZefKiS5ks6StVs4aF5oHoGZ5fIA77KQa4MsmhfntK0Q7P
/nbZpwY9zLY/u2QVpY26vmaP1fjdGtEzGKI2W1sJ2SlfUn8uircmhpEXLtBSWB0q
II8KnzsAtIvq4HBG6p17Pshx+9jv8yLAaVcoiP1U3B+laoPDG82mILBEYBmZOTUj
Ic8ESwQQe6ets+EH9l/Uo+Tq+WOqcmAZBnyrH6w/wV+nIeIxr+caFEJOiCbajCvl
jDJI4/XtFupI8273Lj9DV+46lAcVlHd7RvusnGWfTDfXrZkBEEJ+73vEixpEzl4l
jf/gvaZqqaNuwCEG79E3rnzgi08+dEMH3zsFlJDw6aGiaf8/tVhAaazlrfKw22Ut
r6o6LjGVuBnui9P+4uATUFNlx4dbeM7r2/4WpbSsVB9ahcNP/43Ph2ypI/hqwYpr
KswF5XTkzU6bnTRxuV41cmt893cjbdX9qwO9z0dRPZ0gMzxyMljXUHKHf6+qEHWx
hPFo/Un3nPLHNafzGZMaAGpHMUY9HcFnT2Hx5YFmaMFsOEppi0KiqM+YaxGbR+qo
qjUQUeSbWcmCFceuhoTFY0imOH8dWJaxktvdAYC5t6CpG/k67hGSBmhKpjUvCnMx
2GI0/S7yQjFCyag+agGMCpykaJ/U8E7rNTvkblB2/EfpJCLXUmxDtYOiuiJFT8su
z+uMpY7kmeYqjFpbKZUMwrX3HkDHKVrsCJTONW6qh29kpmom0ZKGsOPBJuVR3lc7
1qPd8fxWHmh2TFgcPBLwa71Arpnxq3jVzPERYSDGvL8LqPdqCfY/O6HfBqE4HCdz
N68vvMYJPtebDCi5IiZqCYjftXwbEgqptbqtpyjF3XHoXEE2cpR5+VbU5VlLNa2H
RaLTd1H9EWA0KE78kcUfMEwe9TsbKMKEMT86nmhp+datUraWEijBwNgKLs7r0B+j
R7goBxwWednRVOmC4qd5HMo5b1lH1sUlWYu7oDHJhufh5InWBzyG9mg/2rV9rqZ7
UELBEovxUEq03qkFVTUdTPSOxQOfJEp8TaY/7WHFRfNk5eoEqWxoBf9xvL4MPlwX
TQuq0AwBlNUj5Z8lCzouj0pt7Gvf+nBGRJ7tp//11u1wmQWskCwCQO1tckp2mgXD
VPijRvGXxtBu4K99qA90s+SIEZCHwqQD7UZpYxiWURNvyPenedOlk2+3row7w0wo
gxxd56YihS7+qGOyxpUgdRF1I20v+EonwPuUicCrLYQGvtdN9BUQSjjd9O/nIG4y
OJ+enyvFpJ0n3WVpVNT2kdoreh2Tq3FFdekgQIhdt/5WaXYVzghO8OUTOAmZRlfb
nCJEYNxkP+PthbYibvhbwSYbq/jSen9TYMESTZgug+noBuNFR9RTpwkf56SI6/S4
H8cD6JKWpino9IbilU4fd+CPmxDw09uEYnElJLwxjY2NC/r19uSvF2xToIcp2PXm
LYVb7Lt2uTVIGK5N7+BsGzTc4xFHiH2IuYFZVMsIfDR+i9IzrCzNab6H5AzKjhCC
Dn8A/3QEWzbYk5dyy5d3U71aK2VX0DBTZNodVqpxj8MRWugUvH5kGlRbEnd9KWIf
Jlqp/gSUndZEQ2mqHsn+sZsaIbixCuh7a9ctxJTKWu/p8fddFuy//rypQyYnJ7Y5
nrJGqPvJjred0DCmq93iLh2UhzftAoutgVCZRH/0JBIPhPpT+4xk2RvAS77VfgiQ
0hGoj2oU7sxjwi8JPsDWSN6rzjU9oXvdKi1mT4LZheGGrV1zpgTO4VCL4KukWZ96
OX8Z2o33pjDRAWldWGsWOlW7Fsr4/VxvHgJ0OLfH4BDDwgpqnv4cE4YyZfXMglDv
HX87MnEbI6CUxUHPS62bDfCYeoMpmaEOOFNVSZnVVRqsKybkMtOO2agsDgIEsQob
z+ea8PMw01vE/+RH+OmtpACS7jAP+q0uTg9Ls8hOvSD4yiL0bs6oPdaYlX/ZDJpo
ml/bZA67YqqSPweKXgRSMtzk/w9Wxe0vFSG8KoxjdePA09Cx7vdZbRkwFBVByAQJ
fjeGwoWN7vY9HmwNYPuwLlBkxdpmKPVTnLCPbwlJjY41VZJ1RTnufUd5OtfiSshC
gTDKvHx+jZc617zLXSGCSOJiVsxKUtsLjl5yZ1xs6EyH68eJKSW0sjXz6nMVSl24
RNqnV4GNrUyIzMrrZBUxcS6MhYYTWk1+2Ki532oY+vaTnEOLnCTzHGmsuNlB+kri
3lw3ZX40JmtX+6p8grmtJvB348TSmJUfpPA+Y95yw0KqEYJ4IOwPcJt4gTR0oRDG
QbpTPWsPr3EjSqjSuPTW9YBJX5q9PTdnp75ODRgChn3sTdlrN+u59aKNMp29sN/A
wRiOSIsqK3R2xuFPWsKjuIt6dYog3Rpq9W/WQdp47Thi0DXMC5oK2mJjm0i4hNkS
hrN5WiWfjbnaoJp2WsCWOCwEF1xXApfWGEUD9rBPELcKboS/3gw3ZAzFCy5kyaRB
b/6C/Myqk8joJc+lv/+y/Pwn3Lr/fHg8CxtBGT7fWx0Gy6CYJqB6C7fkQbR3uki0
6zL5MgQeyqqTEC2FwLXtv9eAl+PjmbtC72gpETqWG73pK9giLnB36X7IUIaxapmx
htd2eglNWyfJsXg5G55QTN9Sexx/CQ9JHWY3gDf3Lefe/sVWtCxNFhVQlolvSG7S
jkn79nnO3PwMWI+GX7EXA3VNnzGHGYA+zgTAnXXGhonPnT7BfCzsCkI/7wNybR7b
cxociDk+Ry3+0evT/TIa/8AIIWn/NtkG/ae/mmAWGS3BvOXA7J42ZkMdGvnYvBXb
fWW36De3pvRrA6hJ5lzfZ3oWJ3IE6me/6ibXIc4UVMX17mUJtAgOR5rQMwVsk1N1
nvAK++GXwpq6ZjDvpKEDnGvf3v3CbygjywBEZHZbGEBOG8XKoIckbSptaB6UCkSk
6jvSYJLgLTju/1uWxuFDtxB5UOg2hcqEyb8JOq5gU1EYcdkq+hbQGO6fV0e/piH4
RaThzWFNMHpWWP0NidpfwQElpk4dXImW4m4/k9I5+ucCn3GQivmKxUPFQVbpa4j3
xSWDyjaPf5Y6MzDMNSgYABNHmzPehFXkyLYDaGohBxCHbAIf61f+on8Ig+7YMZZS
TBgPlueKpMIrzU2PYgaDqMFxnt/5MGAJOlpWnR2haaBMNxd5YcP72eAu2XVfEYEY
Yc46gob36dJldJHxdt8qIfWnEKMYktlYTYZ+daKBHTrkxh1pU71Kfuome6FiDR1+
i169iGOpypK64sYEPPZEHFn63rkOSrZ2oQjsL9Ynnphj72o/iDbVWjdDtlqsNfUu
7sjmh8wqp3+KKBmuRCdEb9ez7xUQXGBd3l82FAhdYK8XqFK1W+c/DkUB+r811snU
CZAhOpij0mkdiXeXd7MR6C752oOb6tC71i3dzpZD20uEjOdzXWF906g1hhkQv9Pf
rwTjfHMD3IquXRGDXHs48q3xtAq5OjFPr5s6MELhWsZvZCxsPnDg2NI4XKd7EcXF
TYtcRTIzYkiOe6FI7ghmpmuRUPdbYPsRpDmSjJEBDgqLvSLG1vq1FLL2NhFbroyB
PiSbH5hbWSc/NNc4YPmogBFEMxrIU1kA0H0uTd07HlstKHnynDr+ugQlrJHQLQlR
bQ9MoacfgJb48tP+FJfiXzMw6/D3nLVSf6aYgVw66Jt6D+iLGuVLlgh7iGjPlC3p
vAXrA5WUYriZgSWjFGS+Slx6BgfMkiHS7a9SKZOfd53rSVlObKnLF9Y3AxaYruv8
EtXfun8a0IQlLKPCFF3LYt6ntcHvPmdJpcQHmSbIpnzsSA+64qlXCi0mFiZKCxmc
TuoVcK21megwh/VkYpf/xAGS2PXH6N5TBAYSwG7e/jSEXfHBA8USHz3/3vVh3iEG
fT+d75HtWa73PRX+CHH1hVJ0vYhdnKOlskfvV3MxlWepUdiBpn1VL02nWs1Z013T
HXkFz2S69OTIyf6Vi4OokGbOSnBF2ZuRZCKjbeMMT0/Y+pQxZ30brRavZ7iu6fz8
bsY4sFlMYc3MhGdAVl6su916Y8t4t525ixUyyxxelJV2yCHHPIzrKwLoFOOdkdlU
smzIuupt94liLMs1Eo05a+7CjWvYF29wwv0fXnG6S6sTHVT7AewMN5xNOQVDAxK8
DPtw5hBDv20GAfGwY6CZIPyOU3zpxbXp6+Vura17cJrzMPoDbGywnS0Y5FXbLksw
kryVUcuAMvbUQhdASkjHTEEy08uyMYw2ElfYGgUNMP8tUB3IbRTChCrAe9JBPxpU
JrsJm5t8QTHdrQZtryZ5CWzokruSqdvRjpNDzYDThjAln9oYgE3ju8d4NLYjvRL0
yn2neoJAMK2hgrl2wc3m6SCXdOW65FbIAQDQ9oyqUE7X99npek4pNyUB+qFtc2nx
frQmL0ldA8QIJkRRSHW7muKpr8IHJ/g6fMc8ljcIzuSvmyAn2w4OoOFSnYkScFB6
ztkvTb2VN9r+A03JUSdZ5O1PmvOz1NFcFBi+THwWOIfnmIkkkfnPULM/v3200NBI
WXxd63YH1Sl5BqsGncWo62sop5k03rPoyKFrR8fdmVO7IanOAK0cGrZ1H2uumLnf
RlURMTha1RwsncIH6O+UDG1KzPQo+KyHJyUTs8y6r/was+fNzCBiLwVLHTfUDYol
/C7SzaNTpyap6pfAylnOpNo8sm4vBBZ6zSF0KIPDLcy0KHhZnUn8sy2LjgGG+4MG
ByRiSeuMDHOC/HfD2lBt350QEOxo/DO99Xg4/1NLx8DyuPPNj9bq2jQrrXX+pPmE
T9OdiG5lKpFt0emfb7j50CftBmECMQqRCfDeYW7KBFsBnSLeBnAphpob8GS/BP84
VcICS0uzS3o2p2xVBBliB388+SlpLQ70P3RGQmysvN9itSAcq2EBhVBoFf/bsEeh
nYDQBLMlNCYHm0rLuP1BFeipCzAzvVqfM8CV9y90FZLzGEH//q+a/cdUXhT/QaiJ
yeQ2cIuHxLWXK27UQbvwXEoYN4ro+QmAgFQjZaRJJuF3q2+zjS5ZEJ/w1IjvsmmA
KKFJNhPrnXx47p27Ha2gZdHm1xbIDGWug2Jr31saARjTNRuEtxqmFwqtPMWzUIix
vj5xAOSte6na16cI7WlXl7TH9O2BkCZOVXEJXOzPRkkAxuqkE0cokb1nXGk0NMcI
T97A5y5+7tKTl/UL6dlA4PP8AKRO9g+OZfnw4WUD7JB9vFvfAH/7Cd7jrEBUh9Tg
SJPSOFPKBzSM1t0wOBrZpaY1/1gvi2sWHtUKqdJqBops0k5sVOzLdTTRZ8HLQxqi
NFBaOaVCu6lhoyvtj7ySOE9dF4CbcWIalulHoJfD8tzIN3hg0fhPP17ItS1tVaa1
hw1vnIZb91Ube/Mt+QrkcVHRYmW+4skzFgrmOLl4WBPl2gBTHgWjPU078nhYOxGE
BDTpi8c0qmO3lIdyisd5pRetq2lFoK7cC4oWyPK09daOhtKQCPjpHFH2bz3dZKrL
irHZ29p0jb80odcoK5Gejn5SlLdRXl0xC1VYMxli/bfYLb9GltcQEpvg0xCWFKxr
WKi71DJMIoWht+zoHUfhSJGEklK4G6jLlmQwkWbuITfpQciI3pySEpgzMc/B9Q5S
F1HvC7NSvmnS/1XEVOKKu4qL9tqVn4yEm80YFQSV+2BgZgzaJFWjqsq4bI08gwAt
JqTk5sCfLf/ulqlAGNuwS+1AraQtTGWGTCsjjMexExwZm845tDd+6dhVzltQVBd1
ySX/suvrI8HdeSiexY8o99RYhH5nfn91Dyz5qEunIURx8CWMaL8nPSZFoANrBc76
EcujPltPTrq6CrrOE+MNuUIBtdciBRYVZEaKAPjuuUwdcza+nw4pfUsvumSLt+w7
Z3CYvlccGW7gzvJ66N8asg0eWyYvTZSFJpn9A7moypU37fC8Wq0mCIcxjQes+w7b
qKKgFPsg41rsb8vziuoDiFaQT95w92fQ/TrqG5xZ5n5bKroBxfvKor3Qt8SguGVy
vg7NMnYWpSCfnpHEcoHz06zeG7ZjxJviBG3Ycux03qwpeUgqTI/zJd5yHr1JjnId
tWaHfBtm4iQVR2hkJLm6ORc4sDcxNK8QDY17JbF6sHOG1+N9i7hpYuy/010hAraL
w9L+w0tZBbBDshSElXbnB20EBJAq++dn2CPKEQ2JjmE7MKfxQmkAZPaeknm6JAYt
40lxG3buf4sGs4azUM7XCZUqiphkKodviNKSoTSRBxnfJTLsOQ7BmtJhNPzy4tYB
9JoCSfQUvYqzYFybaaMnmBQQ4eZridAOdytcO15nt9F+ES7gtloJGJfhM5X8PvNT
AqIE/KN0Ijhc0FWr/Dd9rcm1QOwULaOVuk+kQcYytkep/3YJM87vSz2ZAY39GX3m
VaL4hg2uLtuJDoCF6h2cMr0frT55QM+dXGJDFsCJTLeaSHf8hMUm9521JObi+Kui
LHOmzKCITvSN6YoUv6QCriEWE7CJlv/yAMVcn4gHhA2oEAJbgC5rKm4TEXwJxiA6
WEyeuKuCK5eTMtzUGZ8lJFW+egB+Z+sx9uulq1uuQrgT19DiPuHOQpAzngxXuMaI
T/zWdoYAA+N3VtyKWNKHwKqULNivvKQSkQv5J0SYKpHP/W+vIddgNejrdPS7GIhz
P/Chl3YEh1rK2Z7hw59odg6KZOgl4EYfdCJZ5nvrpVb9KbIXAShVZUwqEhdOUkh6
A2c9q7NuZRC75p+eiwMEcWdTJIAUuQD5/mWqbpGNqiNScV7XOKhau5BkfS0ayNj4
4dOkACPpaFO4JFQhIdFU04Hlx2YEbwwiCDhIgGekEIxW3rIln4bMvOaNNJfzYRzG
YY397OKp7CP1zdGpwuXSicy50eEutE8sEuoiTryLSxd9zgZbAA5UI5472AkZvPUN
P75gGZNNTu1l70lU12nedrxfYUAjA/rRZl8aBI3ztUwJxRexdxhAIXxva6gE/yTx
zxI7RqWeOopRaQ7kDipLoaWzHVbEOPaPM7CmTB4edIl+S4nfY+/nq2UMUsmTtlCK
816S24A3kCWGXk5xIdLKYwnIILW24ZYsNJmlawjUUICv1hYwSCfFI3r9tqxOrrow
zdfGrgRP9fvDX3JJ1iTZrEwxJuHL/3bhPC6pGpuxdsG9lmL/7r3FVtgcTy8ejiKj
Ah85J8Hg6AWZHc2aC7iXPG43X+bZXUOPAhtrpH1Q37hK3DSWw6ouksI/8Q0kEGG5
Nk7OG1O1NpjD2Sw8s+rsIOvq5hGvlmnmbErn6XiNiVxTaY/8x1T+p6qSI6Fw4QXa
El+E/Ge9UwlcIjxFXnXuYqOenR7HI/jSvn3ZOWQlslQAi3KLHTJ53oDpUrTeJnE3
53ntPu3P9djaPozOl+yXHnmkYbJmw6rx15bbgGu55pHIcOpltDBr3gJSfTPMGJNu
XTQbN1Fmvg5fbcld8n6vDiqxtfGrJL7iMfU81dMsf6vkX6HN5jA+KbjcH6+9AYnj
vbrMmb1P2Z2zck4wUqENZLUdYJSTbmER0P10IzudMLuRmpqI+TqyquqU8ZdCwGec
7GIOkyQjuM/OQnJm3L48hPOMQlBAAt60LLXJnluD0FGk3KNTgU4F9/Y5SGio/WA7
yVvFBgPcnZDkP+PglQ3+pCs/Km5Ss9YcpF4+7F2DWTvOKr71vL8JqucvZYooFNYr
KC3XCbNEWz07g2U9/8c6Skgs2JvYOE4ijkPzAjMUk7GzdsPbUyoLP8PyzynjMx2v
0HTg99MtiMwKkwhZR75klC7LkdIbmCXPrP6Ei81HN25m5FA2rxUznB+g8EfOjed2
uB/pIiDeOD0sx+l8e7xfLwhP8Q4JCOF80P2orf9tbfr8wDR8ZVLAEy10Je8GPB+J
7CeR4+maRDK6spYfdVnMEHBTp/UkiMETfp6fs67vl0jyfvCw7plyMHVTo+qm/SR0
23+zrK7qlfYQUUwmOnkA1KV5ek7WGF4JDPRpBkeTCZg4G18Oph81j7gyMOcDUgHI
E3zT3vHElMTF19TTS6JAAjslSU0OT5UMJFiC5GVdf+Osrk2HAblKzjzOT31iObs1
GoEBXkuptLb0PA38Rd6PlwGNntIYuzaZoa2B67l47RLzHGWGre6BSIdLwSyQukDL
iKuU0u7oLEeYqPNOGdy9ne3IGhMBnzre9EP7nFeruJOWE/lLKsY3NPPMTVj4HvAY
3eYpTWl0KBhv5wtbs3RvH1OZ9sK9nhydTpqXzReskZcAgqdJFGFJdCURQgViGq3Y
JmpaGfF1ycMhl19jEMZxoiYxgGnr6ErgSygB6AtK1/+CYc37FY/2U9QuUU6kBefe
5yoZ0S8TqExu2jA7qZy6QmQzLogIJC6/zQ/wpwLTnZo/Q4ATWyvb5Eum/XRhgfvy
uHmgh2mc6Q9C9trAUqouMJdyMYZBiW6b7d//0BLsjbv6vCotm9X3MvqOh6TM8+zC
uKe79tkH2e8rKyw7QtsNxTXpNJRTlJGNjPpqGy8fmwPK9IHhD+/RDW8WH35eyKka
lpxpaeWEMoSUIeO6lQxTs/W/Z6NaN3k0uALKWgH32B6BZK+a26L4FfC7Qi1mB7A/
q1t4WVvkp9kLDeIeXE4Fg2JZMHfZ7zCFJlREEDqzD3kFQ/Xa1dzMhxQbolxg9pQi
9/RBgzTyzJQ+mV3aTzo6nFUnC0r63BKGxdtPQu0d8RGRZLZbrtlRRhF03xNeSnIf
sYSZmq/xTr06bPNbgRRbdvBX1XCqXodIPW8XpMnoZIAHJoWgAfRBvCtCusMjUcnb
zAyOMdALcVEVKjasCAXmddq+0wcuFh3bjNMiTZEDWFblP7Wfoui2+CzfUvhZslTY
RsQfMm/v8iLd/3pKBx5G+xZhqOQy9McSkEpUDM9zEwqo029S10RtL0kGqmgweqo4
M18zOsUSDSnk7gb1FlgAHDNQGzfd9dVbJtdrvgRsJbuVdkexsdRlVoZ1cSkjTMqd
KJSZS3/5VQMBGsoujtlJPWzbhOWN1CZe3ZFDos4aHxp9SmDdkCeUPQj9Jwwwnq0Z
Olq4jiYOKWJMIh3wUwWFnBZr1rYIE1DxgAXzknK3Oj8RUm0dNEvI9DvdSz/xoIoa
sTp24KRaJNMlhrI8a7wlWpDGydIW2+Ooz1ttgzme7rzshExORVS2bHVnWFLzY6u8
YCPKqqfTQvPO735qZy25zNxzx9P551ty4RHWP1npHt1vbbTwQlN0fO7P3UC5fwvt
J3EkuqfjOVJ0kohsO1duI53D3GEZ8sJu0krTJkv7DxkaBh7XDdmOFbK/KX1Md3fj
4MNb5TMG10KjN5zkSdDtJ/CfKoM++b0PA8CK+UTFmz2ZeiuahC08NBq3XRIMe/Y+
R610eBGfJYjBAHDvCfp85B5ICNKD6vf6KP0+A61HR6oQT7neOZ/BOZH65q8z1ezk
FSnawpYWPZ7HVBf5Sd9SLsWnx48+9Vd69P773zQSiCD+6aqhFyQjYCcG+2sJIw44
OUKlkPpzXD6wdaenlGzYLc8b9aOqUKn12/hGoxfv9reLhJ+ZyT9dipp6tVaHkocE
R8ohgKmGar5YVvFQwXov4OQteayFRFCzdFiZDLAL5H0YE9q7VCV3thUXQ/qPt11k
s4V/IfW8bRnoy16Me0IBHBVfthKthPO3yxqHksg+7LA83gzpBVwXRhlichh/Z/mK
dgkM2aylZxBOpNilwUdyEXhNgWuO7jkcQyLJ9jzKnaNZ7YjihL2RloXLoVUmmBOG
qAgDC/vN8EXZ7v7A1DNZtb6uHPCY63HD8nw6mCa+hJ9G9l5UyhyqsRRXoxUhnjng
jcdWj5Gd2AXOj6Fu4Se1waiTc1/hK6WgEIIX5VPDRVe2F2XtNeGUeu5ZI7tg2dtR
QQowIG1vF6Noi4qVmVv3gPGe8mWq9WLFVy+S0L5e42e7zo6WMGgD27GlFQw0I7gr
Ri1hgvD1JzfHbuMkZHEnHhYS7sJ908nZQeVBetWAj+6rVdhHG4UuvlK9v6e/a8eT
FWCzYGQl34O3oT9yOhIDUz0j3I6GfRgQCDKafns63RPaViL6etwCQxFySGDZQnI0
maTnuF3J+ebWHZgZ7ZHv9sLO8rqv9IPOWOanyjeysmxTElzX2LR4R/NzmhLgF6nW
yu0vOuKPDb+yTJsTra8Uc5od+6tqY1qh5dzgqly4bkeVeHtP+1LpAtM2A0dXpZWM
P5DbYj/L53OuzachWcXLSHLm8QJaRi4kRSFjOXBffEkuDiZHECKSCZf7C+gWkDfb
KCGkjrgwYEgdJl1kTQrONOnwhUvH4JSLXdV44s9md0Lz6+Bv/AlUSNplJ3UVAu+C
dv3kl5jSfA56p2n8EcIEiqZqLje9db4Z4O/mbJ5uNgaQ5lMD6Sys+VXsUFN3kgiP
/N8O5gjEB5CHmpwXSvbgWD0PYg2x5iJh2CUFkjkSpF/1csLdV2OSEqS3FAEEFwAE
RnXi68l/n3wbEIdOskm37JaBEfuL6YXzWRyrYxmQp12OB6c612moU719hw1TjIZ0
HEnOD4CVIuni6vpqJleclYFBgqtwaNh00MfuFt9lMx7LEX+wdvV1tzr+YX1OlReQ
htBjn7JNG3BSNzJhQVC+3sJGkqbwORnfb1gmlVdaSNbwlf8xKYVz6KSFd5vZy9YV
Pm+7R40BXo2DF4d1LwDJAny5Qsbz9wrcIr0sww04xTzkaoAVBWRlAD6s4bs+7KoM
t0QMT8kQ7cAveRWAmj1Z6se2HOF6p81eKMDRVHFo4k5KvC+RrigvSkra2OhKgcMz
Mh5GDEAIOYAjnfb86kTO3a1XYVRKfXoSm52aB+49AUD9X2mc/yVKFtyrMI306cjT
YTGDg+twD/AEy98DhEAJ1PNWRMAk8Q/MS0erR2U3IIyu6oNsUVCube16NDskscm4
iSLdoDXMdxT3lAY04zq1zrV2p4vGoA1SFPIEn9VYQsoay6XNeLj6s6gWXPModpbX
Yb0XA6KFf3lQY1gstFzqMKOXIWMyCdH4Bb2NrNUQpdoywysUmAGEeUEASkZavki7
cyWay5emBGRyZlnOlBPVa2/oTs9lgxdwpb2Kr2fmtLMFMWOipXbLwzsiYOydKU45
2kPzvFUB7gqKlOzmRjId8XnTpogSMrAa0aZ+1a9sZis/yfstHI5QFM0nxTmk4nNC
1W7o3vrNfWO/Xvr9NGHvuXE0m/Ae8FhgfOdvGFInvfueqyOGZcubunI9LahTXb9m
MDS+2afcpL0QIWWwFtdIRhdwLoJd+9RLLUPktsR3EXUxGllIpga6UVhiWXna4rK9
V/GMXedHdof7d8hhDJF8ZDKdQ2k77YDU1QvC9y0O8aHD3Zgr+b/N5T/HyOP6+fK5
V/r7DFzvXkKHPl0jg290kmOLoR5uqJsNZgrNMzq2KCxpD6a0lQ6NerlOr05MylBD
4C5mq08sZtu3yCz//yXub/iRzMZpt4nohqQXkUUZOvOgqAFYovBhwSS98S9KmMEb
Ai5FIJ5jzqsaLbJP67WqthYwaBvgq7v3dRpMScBwua0O4KGDqWjv5v6WS7B808gk
doAzHlmyUoaelE5o3cz855pFfDv4X+bwvXqLhzeOfE2JAZJKNk0yqjFdZapOmxKn
STPxXFLEDYLFuqDc9/DqtBzjYBHlqsvQMcdZnP1Ym1zApz3dqPe8RWUwhLMDPpHE
Et9yahHP/E7BKjRWjBcTJc1TMWBMLECi0ukJruE8sYimAFnlg3E3YL6ubOqiNgjR
3+SmmH7O3hdUSgcxalWEQHdyxKaFzR+Pod4VrPhCdUZAPGDVn3IWxpTn8NNUJKB+
9oBe3VjYSb5iLs+bgUSYgM1vaQBxexqQNtkssztQf55/q2IQ65RtAPjUwfsKdqDz
UuolUuqv2ohJu1S64qEzDiZc9CWMrN88BpCnor1/FcLGPT/5RTI9cy2RBD2RZaDF
FH2D8XJiVMtxiaRiO/hLPXZkRu3RLnGUSj9hp7Lxrn1j+B8Q/zRJz8TJbZRKgM0f
Gybaym+fhgSmOB5hDetSZGPaF7aicCWPf83DeupSFBoNDTfiWjy9bqB2FKaA5In+
gXbkz3RVsEfRGatBA/Yi/5dGc+IRDUupocTVwO1R3eZLWbVia288kfdHD+SekuUJ
IBTkUJf0TJGXgzPq8FT23t/xUFIw+ErDpWTHxWRML9OIvKnzoJv+rUKj2hT/DYgZ
onMm9NQicPtXaaTw+HsAE9LBCNeOUcFdr7kBq510MNzjpScntgk2DeoVRczmSIf3
5oeBQtFVZI5731MpGtBopRTqJUR48Frk9kdGqNvwjS5TVXwopEcfQ8fXyvRuy/dI
wIYUGe5aY2yRlBQR7uqaKEd/ENnIRyFZSmLEUsA5c6tj7iprI5Zl1CoonNvSxvIW
ogy/yAGWOqOLD4ZHb0mGUWoZPBckHdP6TOBXTbfvoxr/DGPeWrxsZUeNFQbBXODP
DeD1TcqLaWkSPyiG1Q4xeD+WX0C2a1VD4rFPBZy8QoYLh9D1DNZqaAUsXQntGxFG
HYQwX+xuJVz2VOshz0cdqRtinW69clVIA3RxOTlfcSgbxVCMxjItZ9Si3QYYefxs
xCrz3471VvXtnUkGtl23r7q+PuvCq9polLNtABrewToMo+MnqCUsUAGgG/M0N8iS
YFzaKrZc+3PDwswOgANrNFtiU8fchfhifbIrArXx3RvhiclMOvT1jGGIped+T5iU
V2b7AqLYgFQnLiV7kYDtZpgXKaudoEZ1w1g1dNRCUktSx4n98aGCoPoO9UnVoO5Z
sPom71K8AbKJIE5+RT5KfHC24JIiBmNnlvSepp3zeHrE5jRkIsMHEosxgFb7dLct
8gwDZll7ClAwRFH8KHQsWWPPcJ9MPTXqAj2kIwJjac4dFMAcCvAWCvkudo0q9SiH
Kw+ZOj4Z00v8uQNCDybigs5cIFC1uvc3m/AamT/FsndwbQQ3Q9VXUWlmsQ9Me29x
HBIFFatGkvtYHHcxjGJ4wAzaDBvZcTyQ6QjqxXRzza2zyPtLKoHdLwVb3oOIm1Gy
+I1imnkhogGKJuz7RDDSZ860/jw9+FH4YZLdV3uOWbwVBkRKrRFE0/A9oDQCmyPv
FSRPDZORVUjUVOId2IhJWZuXUbJu/6LC07GrzUI5L0qjMqZco/hIVvplG4EavTCR
OQWwitjgamcJkEafuvuQXPiWcDYHjbIzegptXUGwkP66Kddakr+nZOtmW5+rmrVk
MQTJC5QbZ1PylJv5IY0tOBgQP/cKaPAo5q/DHLXcPycSowq93/u2hQkjJeZfkE6Y
Ap82HVulJKhTOi7TbJEtbL+PYFkdQwCWSWuef2XOHfUieneNB4EK0rY+1Jur2V47
Bkr0zMH3laNP2pIXOemMDjpRv8eNb8fnvwWOzs5n0IwfCjxKN4xP+tLy1JbqR1z9
9nFlAekLoYaW3gl6xqH+9at5WCYC6AaZ1Pa0FCUms9KQVoopdE3I+IwcQm22eBZ0
k/c3bgHDWxZNW7zFVWHEOBOuCWVk+g/eQsE7ehz3a3FD7Pvf3tAqf/JtLIjTHgYw
7X2Wv5I1ML6VcG0NzIW+vUSpLHc5ehHM369mtEbeX+/nxphNSVjkmj3NYz26UwQy
hH+Kpx2xUaODHBZBSfAyYBfLJxdBPd0rIZWN2BlgzCbiUA7odWTFugKfRuLXLko1
X5PktQAsGjzMcW1xs/62H0e4sBNiArG4X2kHDV9dItQ6rjvpdpxnrqT+88sRIt2c
4hdRbe3ahg0o2RF5IpQctJgFJmsSBywjdJe9MAcPkoSc8ijFHE/UyNAE3e5Yn1J+
LiF07lj2yk3L0hhiIX4X9/2h1bkjtCASH2wdRD3yDJ6XMSB/QieqzYOvIrJPKDSK
NAu5kBWSoNx6ZA0GTIhZZI95zeLHPc26S7kDkhTwcYSIQzg40Zb8i6TMwmp8n3yq
pZqv0//xaEcY2m4HO972kTOzKujKmK1lFG7tF5e270ZkpjDGPbncYsk6EUZJ/MyL
L0/ErPvvP4tRxZiToS6BNYtJFbkpwScxlXZUGRdj+6Q5/ideUm2lekvhxrhpmU6/
GvDIay910Nxwpi3twvr0Elnvw0dfQxg2bOg22uJgJtosMJguXpFNRBZP6dDvb63E
ctF+IIjDq8IIryWo/TGOlNL6JQAIVT9rKwAceRC+jagXZQXPVQ1wG8gwVdzGQAgT
rqQ0xr6BU9q3LZzvk/iH6IkyjfKFpiHDE8GrvalZc6sJ6iZnuUkqzcoEUVYPFhgZ
m/odM8LH0Chd4QE65J07PoulCm6N5/9Crk9VlDTJ1nbByiIIeZk6iXPT87PrM+oO
Tl4madL9EO3M7EVwRC3mIqDslCU8P2hUY6T72W9xdtcNGQtc8XOKpDcQh1U6dEok
2RKnQBAGF0oF52H4xocz3u++Spy3/6p1cma4fyP4B6FfDzQ9k7yMsHmOzHX8l+kc
F3OPp17KsV912Z+se345Nu3AYwf3/SKFgIq2lpYde3LF1G9EPwRm4M8OuOShbga1
1337UBI/B8vHVH0/MWaTH8wS4fU2PFEjH/EH0oceZ6M8ZB/JGwBbGZzTdMaEuWn+
53JrUsQ9C1KXp6ssTBuZpjnRTsEkoLd/KJCzq/bR03Xu3KMl3MMng1rWZpZZg6Xk
72af4nbA3w/f07XgatGvwNW+qmE3IZ5uS+qHBof+obIgDTHKygQsm/suVqBaTchW
l0nsoMgAXvIfPcb4UkxZgGp5fj4yfpvngrrpnFSaiNMs+Nldey6/FFZrkbs6kmb/
ZjjxOt9daQVLxU07QiRyZeIFlV2F4gVVOC4rqa1ZyhiacpwP4WqzOaNyhLqYTZwm
j4AdkPqOIEr+90Kzr2jGxlHAJ00/l6gysISupKiS4RSI9y8sV9NkwYEwHmfrh+1s
7BSdVdZxLWhP40S/3bfK3ZkfwJCEjrjBpzdwJujhueQ2vE8Oxfsdo2xq2dkvXumT
sRfRhvzvt5oFk/+vbIEHEDlQCzWkEzF4OhjGpPiDWcU3Z8Oyzj4rLNvgyepxOFiV
GMiUHXMq4v+9d1fhoYuZ/d0+DIoAlA0Ds4bPgQnohrsrWYCyKHL2rAV+kOCnFWB9
WMgfNqP+vKo6FUqN+VSQAvszhgTp4Pj9utORNHPsN1wqr+M+HO3xRxkNNjfIa1Yr
NUIuSboUOEBffjg8DPxqhUvTAFl4xEJNn/4U7oxrP39Ozh9/J56hRWnYnE5yJYWT
vHDFN8LXytQBUNRjCM5U4rqh/ngsRgmFNZzD3MokKrzy0MB1hg0mm3LO3rhSyQo7
hSg+eAs7g09/Ke2VXQZdeTrUY6toNKygCYvAfvU4sMeRa0AikC/w11BoJ/jmnx8W
pj39x0wNGFuc+gt/8Jhdk754RMPCYTJJQGYeY3vFUtmeWA45dk6xFEfBebxCoVsZ
L2I15aNE3UIzMghKVIlOHxACotpBuBkWG+PLj46uTw98HXDfEDtAb2pCkOLt7aHi
+NqGpqjuRxDsFCv9Ep+FXssGefpEM8ORG1UotJ0zRvM+7lVZ2/e/J0XS5qTT7zx4
q6RWjkpOjNfeYI60FtINQDuGjl4qN6deI63og79vR1cAXdMaQcGwKNnNUgb8suW9
7d6QAKzKP1mwR9nMo2tKnoBwhTEZ2vjgHhmfb7L9PBlcyrTGWqSS96sb/3tNW3LB
5e3a4vC/xdCCNbJWQ+/m2p6zm7TOi9s6XQWl543FKy8GTwmGqfIwjmiwa+38SWnF
GGba9Bk6u/MjSHvOf82u/8N6pve40SIG2b/u521wSYeRSxNz8S7ssm3cPtC1LXW+
+xyiboe8FarbeH7qag36CxbotGQZhVy/KQCRIzABzZP2sOegBQqJO0RN0yFXJ5mQ
VBhbrnL/XybB+x4lQqcsAFWSb/pqA+k8bLf1bJ3x5vgt8p2N9SkquXo1ooi1WCrM
IWE4hvCw6kjgHRFLyXs5VpkY+EvgtYgBMjF4Cf1bY4eeeJfLG9+CTSb9WkCzgccg
g1hJC2AhxdT+t6uHkuaJscdJoIWMTTi51QXCHFAMvCm+Xf5Z1vhjcWHNaCXkIpdz
s9Mh8dmXWSh0T2OAtnixc2jMh3xriYpPCxFFu3tq+azN+G9qfMQFQi2uIR6YMNGI
U0aVqB6q4kARWV+l11wOF1MAMeWf5TFBPRdRBrZDZpAdYy9t2EoJSpxOWhqrXTkB
vSkSfL2NjoW2DLrB4UDmgpyau8uzmxLIsUKV/tj2/T9AXV0BCrCTkejt35jsqBQH
ztJufrPcy9o4uqcGnwo0eof982Vx5fbDQpovO7Ib+Uiw0LvhbotWC2whK8PY4SjZ
8Z1jWApiRiuMSxZSvbwodBAvOh9V1iKogrjieIEsxJRkfVv5GGn5iLK6cb83/1M3
XrTedELXo0Ji1+LTlgI2Nzi2PUcLUiltMtQI49LhLyCI4/UCqJg5yF0K/ETENFfa
QQFuS6rv4AQhCv5vjud2b+JKPrqwhPbvdGuc4qB5tXOWOeyk0TGutQesGG8NLPih
h6ds+Yzb2RGsK/DhnVWORw0+S8AGypBsnYHBvwXQZyZmU8H+7GhqdTV8kxXFq55Z
vhTO5xhDc7uBKZ+cHXaCGyLQbmiimhkxeGwjx0Z4rfkhqc/zRxRXGIaOomcTTrR+
B2LpNTcLO+UHFjeNweAXZi5fLus3H1TrDvw1ekYvQqcweukgedC+L1d5lLgoZ2ho
92KoGuAN9chdSLcfpn0dbDeIohwYRcivs9HYqSuO8JXiwPIhqywstxJabYlZtSnx
7Y+ZzrukMKvLRj5xctEv1i6v/UQR4WQ8NRaJJrrk7ABV8UoMCz5RZSttoi3yqr9T
LaiNvyD7vkOXyqrIh5Fxf+isn5ARx8y2hlS/ZtgYCb0z+bZRVkNfK4vkC55o8q1w
RaINT3aTmYvyPyCIawhszoz4eWWVl9BYq7GuwoewF5Zzeda1hW2Ha23PX3Bhmlvt
qpRtV1iyMgw/Rf7qRjkBO4u//k3+4+pZqiF21qeeIFj16Eup7pabVHFOjyMo47Aa
FrB3eeVDDkhR8i2Mq+HBPdKFagDJqitV3qj9K7iMKjNa7ZzNEZ/vNvgA3AVUO1Gj
DQJnKms2lQOZTOo6yPrEiTCFNa2r4NBwQhR+bE53m39Q99jo3tvg4FoKt3oEA6I7
A+OKa98pnxugKnhBg/Sna3FqfWaptR0KRDqcW3Gk2e/qckPxJo6wbS0F9u4BGrFZ
06U5daiBw/16rM1yrKg/FgQVdYHZn59kPt/SdNKqotx6LksrCAdRUrFwKuUkRwq9
YbfCEED5AXDupbS8S92u+rJWf5zMhNmEzE1kfo4RG5zAtBU9480E9EA2d152R1lz
AEzJlE8Rvsnqni/kFhp4ysPIyCURchzXeabZjjDk4ChvVwyqB2tRJ+nrHGMUzlbI
pLbxhQsIDJTIjUvl6+UNJ8n2i0eboUZAoSKqBF41AkiasiKqi0WvRqakKsxeZaZh
RWrZ5vsfT7vhcbpGvWIF6mw7el2mMotK8nef8iyskb7Vkzch8DAtiALfetnqQDWM
nyadEOBsdxPj87TzPztnVYH03v6yJT8cfhRo7/2Ppvs2MKl7Nf2O3myy2L1mIV+L
Rt3n+3GmyLIN87d2bT6ZM84fWgiAlj29vgrVTUNCscPJCnauzwFTSWz4x2Wrg1yF
3B23FlS4cmotlTz3EEehkoTVbHv/7/svoKZgPMjn3ACHV23seM1TAW1udUWmJEti
9r3qWJXkckfKKUpa4Tm9sZEes4hZF1fUbbINC9d9iwpboYmmCyUL1+4IHde5NeNo
VriSbZpDq385sN8QBcQ55G+dR1K8v2QysjwpjQMprVbae5yj9Ahmkla3rpS97DgO
RdSHMPCBK+WwU/lx8IWtfzrVmrdADeKCFhgUyp+fGlsFpczM4yjnXpxBeb1V97yb
VAF8fciOTK5oKzeTVUwwm4PRoEymKYtMNgUmiF8hC64ykbW7p20UJzlHFj9RYOQ8
Ogb2Dls4AriEGOJIr23E2Fob6T7xYjqcaGRoLFWUnkpce+DC8PSIf6ZicG0R56MV
H5Bv6/ZGZwyfRs1VAwy9RDR5m/gnI5OnqkZaxXZIIh/aImY+8I4ZnB1f4uiQBxR+
vdKilqCyK6SkrTR3+LzNrAOw7mxT4Rev+42D2qTCkxdkxGfQjT/hu7qPb8NR6ynr
cY4nOnnulnK70VqOdpNeB9XU0UxfQmeezq3WfYDclp7shKejq/G6BLfZL+HEuMmM
sXyqRaIP8qL4/rVqb+qy4aq3wWjI43rjhfxJv13mT8IkrhjZ8bGN7EodCk2sfae/
nj7AaV63gIblpHKwTPlNKP9jA9zPOXmobfg4bm/L6NAnR2vEPZLWSc5u+l+OGgRh
+s4gEjZsAx38z3Ytj+tU7uFeUuk0e5lVVXC1R9WQgXX4bYjLQx31Hl8cbYX1Nb/R
2pNA+I8znLz8xG1Fvc+AymkXgOeUWVai16IUjpCevu7rhhBfwKZgsC32/ChP1tG0
hq/MlHtmeNqxXoQFGRWIFji10wYYLCROzefe0TZkZMRTdYg+raKiy7fa6p4g4gN6
FUrdzHLNgaMoJE0Qg76vvCIJEPUYQZXYwTRIiQkUAD5PXT76SbBsYJ9eTKjlTr55
RDYwJlcmJSsePAoqXcvre1XQv2f2Yf4YcHLkmYAudmPNmr15fzeJ0d35xVFP295V
CMmcixUirZuOyn0bnYvOGWOALdLDJi4dMvlYAAJf+oM6Fd1wygxTnjd/PgA+ndM3
mWiSpT350wQo626dgN/N+ThGTPYE+PsNfUD2G3srbqnSFD+6Z4AU3haVwp0v8T9M
t7tu8gUMHZMEzpUiVljNEU9BWALeSjTn4ZTApZJoKUwgqOSVF8thVAUpokYWL1F1
p9CZRXFRfQk7nDkALX37ebXh6yQdcjkgqbg1bDIiorRreXKjvSAmdxE/XS4tu7pq
YaR5xd/UNuadbc4jL3VnNgjV2VqHkb86CxgmDNkptV1jfxpVIcunrl5Kt/iySyR9
H2h8pELqzyehkumB3RrP+EqSbXzJSJbUyhlOyaIawFsBxub6+iEX91/TZQUUtPo1
ZdgJJsxfXkVbOwCq8dMKNu4Yjztieo1iadSQGn1BPoCN6yy82xxDYwEyEj7ey4yB
0RN0CfMYIwUg7vZrTY1dCFyifIJ0G5XPkViiK2qHr4/HeGflYD/ms8KyrZP3uuVF
ZXwK65D+r+tcC3zgnWbXWSP7vfQ1bk9Kzi2P3pUN8Ut/q0mU9S3hwTzuae1LIqrg
Pq8IvjjaqK2UrXK6Hiv3azLuF2JzR3pqyO3K5pCAodaj6Ii0I6TRvrC/LMG8fE02
j8k75uHwkksGpZlC/RZuG/EwbjaUwOBjq8W/+EQJDicu5KI6tY0fiUujyMFMfh4E
jyGujGtyZrwFQvtSHF9BjLqi3b9K4fj2ewGbSt7fmop3BYDULQZoUy8sVl+JQ+v8
yRq4Q2mvPcArlKEV+rAbEF2fUDGRl+NIrPqgR5CxZ96QuPOxCitLx47COVZ6Z6C7
jRGJhrPhSuo/e8NfncJ1qxAe/ms/lkSkgNxtj+hRDwSy5j09PniilZDlD7pX62b9
VOLTKVMSZKF/7Hlip8nD11Sqr8a8ZC/3zcvMlFeXz9zU6JDhF8Z6KEiPetiz839x
TnCMLfyJqfP5vwOkXCpzyK7Q4LX5uk/g5KPExuBqlxdNrZ3e109ofdJ6FproxNHt
EVLyvn4tCzmFVFyDBrDJba+dl2OA5MElJHZZPHou/zOj8Wk7ZLTzYIeGVAlUqMWB
Zn+6Hf5RmL0mzkEMhVpn3YEMmisF2mFOfO1DDHotblz2Y4M7lldhYRDVmWk7VrgE
2sxnp5LGRlZAp5gV+ZpAW4jaTZZR6H73CBWFQ9LFjJWv7L061jIkknY1PLMtudKK
jPAa+VTC4AXIWl2OPyFw6XlF5j6Ycrzy8OHJAg6bZXaS/Wep78uTLGNio1c4gitD
9Ogy+hw/S0qMtWrvAoIo2NIgFalOvGEqh4Joq00+dPnogAYElKRGfaPZEub9yJEv
V7L65TLJKXBBfNsfdGkn2rZKdDB0pmbLMUtvSRXZ27nL4eblyQGrDlsxSGcO3ja+
B1CniGjHLaPkjl0Fc2UWT9EqxeJtM1VgPxjdE1d3TMJ1Lqo6/3NK6jYfZWd7COgd
KhBET37v0kjpWrMvWZCqcaH+AbCgCDf2cz1voFYJxH7YTV3VCLMFWaMx36D6UkS+
k1RUWhtX/6O/dAzFskDyCZ/oVCAuLgNw7RLs5t5v40JnTG0yl0p16prJ78GcL3MA
dpPpaxx/3F43z0gtg5Y5yds70a9NiqLeGlCJsUVbfFNO1JbI0ep0x+/Z7NdBS+ta
pHWRQyTWIj9IFbcf63SbUfkSkqy4qlGokFaD2rOMAUodeeRyhB44YAg8pgRXUtIi
IWHKOJg+AqNyZ92IOKeOwJa2QZmo4L5gMbmQfDauyWn0pQqHRkE2yup6WeqAHPou
Qba7nML9hvzyT1J4I6RQbZQZP3AYRFpU+EGtvD3r6sO1SEvOo42JpWx784l8LkgD
jriOyHHAw7PuPDTXHbRcXosAAvKtreY7jIiHenprHcQ7zGFZmZYSemq8jCd9W0xY
VNKEirP9w7lq+a6ngM0e5WJfrYEZX7Xo6B3q3FDEc/GCga78h6rh8A2JPdLjAihK
rUsWWMB9ipdXv4DTt3Y1E+PPsBUjfQgxqkyHrvlj9U6J3f3ocSqpgcvGU6nlGZR1
LbDhu1m28/tgx1UoQcz2fMjutdUjlwS8qAE83RgSaH36gVR8X8+eaxkTLtjNFv9y
T34m/oTa6OWdcaELifTU9THOt0GK1q9SJYww90vDP+idjPrTY9hntcrE9t+zOJro
mq2/mEukhOFC836e6pRLmPutWtj9Nsj7E6wvO34W66tdmH2+538JKoUkXa8xx1uF
Kq12SxsrQGfc0kjVDU0Pw/tttG0VyCY1Z+RVOra66n7Lkx7Bo8WCUqo/sJPf667L
lWnB0o8VvBoP2ISbemSZYkqGdeRLFMCbMebuuS8OLzazad8sDeEDsk4/I8qCNj4j
+mCV81J6brs5aCPX3kPXsWtVJxVsQGQUYvt8tB4fzkSYcuDV/YLqDcAFwRh3JN9t
cNHVAJT7sg1JuvxrR3TNx4oMxbwkwCEK9cg2douJBAqJI3289UzRjCrWebA7Sonv
EqdWki9ruI7Wmm+9V/6zV3RhkebohX+hE2hwjygs3v6wcyLOcSfpak5kzrJQ/4Rf
hSmggBxzjQcW+p6uZhLO1XvxOes5z58PU27RvHBPpdUHr06E09D0ZU65wYmB8Yfe
geFQHMjiD0iG8zWmjaa05l/zdY079/gcw3C+OqcYwtNtRXr171rRdqP0VGh6Oapl
CjVLMKEbMENZIXF/T3BVmkDiqP8b0IB4uqqvNAZcCRne4Ckn3GW3x+Hhler2HIq2
PasChtD4bt97TufJ5+6cPwZoSfAbRJ32wUdbACtczun+m6b+GKVXEAfJTCkOGxRl
SqN7weLu2p9bM12TXkaT7YAR7VoDvueLnyLhuulaxFR22XVVjJzfl/qvMm+ySVER
sEKgq+m5s6U9kBKmrSm35i7VRETSyOynz6FE7G/YWBo5vzR9F/XGlJgfD1Z4RCko
SELYqfugtmbbjoJo85icIBK0Zo56LcFvw+gpgXSu35A0DfaveLeU6PhRXOgsxl1j
KAGFCxDJSuLn6RScqCHFHQYTSr8XxLgMjK7Ct+R2wK/Yho73+k3H7sifY8bAWrRb
un+B4hsD5yw2Q3XeMkPAZdvPhE4uEzkagn+sVAiW7nb+SqsIBhZgQ/lsuL4qBfNx
P8qiHLDs1NjgbmbpSCKD0zESI3GE13aInY99mT5EcPPKHWx1NsIx3/xWSO+zoMQY
z3n6EisBiBVZXaawWQEP9fozvzBWSLqhzPHQLB7WneXs0UGVNl6PaedAUFT2MHEp
juuoPQH/uWUaX4lAu0Bu/LqufsRtV5S7jYV8MZDJugpc8ObBqCTH2eMwIgaIdgeF
XIc2c2MmapB+0uhP53YQyL5LBvS16RhhVMY4TKXn6PPvsBnAa223Ts6qXCPxM49s
GVlXic7H/Vo80PEoQAUIPZqg+/KAuExTUqN82DQLfkm1RyItwXyA7B1LfIZXsjLR
sa55X4SPBD4+9YhmRl5R5aYyGyXublBTzDOOHf068O+sa4Emzdi15K+Yt1kSftcd
ILFLB7jg2vCfCcHv2HUHzzNtx70Dvno2PFhWXhTt+YS87hBxgjxZu6spnGkj+3Ly
cf1CvTvPFEDbtDUG4HI6ulXJNySDc6cCWoguZlyAJV+J8pXrXTN8+eI0tBHMNflY
pnqFnmUEd96E/H0zvF9qZ6+/a5SCfM4mdzDfwpFUUdoJw6CkJo4ir0WmgEi8OfUO
aNAJDiPGTMRWruo4DylkIaoLAcBAKl4OUURW97m59iJAsQnvgLKvunRo+dNQHd08
8sv2URLLH1VY1TPacJWVZXQrAtBn8DEacIvV486dgzO6oUFXxwa6h/lxbtaU0NPs
RWw8B6upqjXrsZ5UNDEAI3sfCBg9GV7MvUe0E1FiWJItbZa693w2t64/HOXbnR7j
F+pKtGaZcqvdDFowtVZG/D5jODNSp7RtSFR/y7OW2QmIXy+jde45U4f/5KbndPPy
KC6dAgp1KzhhICheForNM3VTjeDbjwV6Bb64fxyDGNRq3Ek/a/y78uuR8Hz5Ravs
bn0H0lOmsjF3Qibr6X/Upw9ue1RTelyBQMN0efiMfgEUI+2Ga2jO/1Dry5R1Rc0v
g7fo6/f+iGWe+DP3tWS5xOp3TaajIAqnLIVVe9GqowzzkS/Gv3Q4c1+0Kx02miSY
7qr8hUJQzxx2nIoVU+p1wXpCtakJoco5Ns7NdfYGApZxBnY5riP/QjxwQ4BsmNPh
fM7WR9q9yKS6RR/yO0B8Xu8goKxS82h4r5Lvu4Ct2CF4dfOZ++Q6ZtH64t+5wXlJ
zgPesjYaDo6NC/WcOtrnKhWUksesna576hfrKqvy3npo6k3dtegp6fG98cKpJDCp
5H8YPj1oaGpf4E7cod3bLslrg55E4a9vff0iswY38FuVmW4+KIKaV79Mjp8IyMT6
qzNbDXSLiVVREo2EWv/e/rCf3s6oWAP9Mic88bYqHARxcvItO54Dzhp3TOa8zArS
9cRrWXZTbVfj2A6QeXAykh+GxuIwxAJarcy6xlUzTcQKYOZ6Rhnw5y0GGWHK5lLF
ORZpo2I5zRje4PJ8zAd0BBiRHCzKJFU4UsgZ0C7U/J4pUfKmfKwX35YfmBRFHcn6
+lsw6A4qeHEL36Jxza8wBI/oiKZqqaZuYQHHro8uRCH7Eb8dONAXqANRrTP9bv7/
KLxMflujJE7sd28rrN3+02l8kNKZ9GA7P18C2HuchKkgUxRaweM+c15sOUpjLOZC
QwrxOTdXR3p9bmw1/RGiGOsWA/e6Cf4I07hj78gRS+KhEXuIiCqAhqgZ4H9iZ30O
Xdwo0JQ4AFDk69DV6vHZltYp9ZQUXMcB/WnMgq2vaO2ystIl5yz5lIulDaFVo4K9
dW68BIh8CxUhsWVvYJ5xEmFU1v+UkjDZQGwuuZiN1Y56uo+RV8fTC1xgdeFBsv2o
H5fLOd30YsAy0hCu35VrQ6YXilQXujgs5OLRQeGbsV23tQ1y+z6Dr0gZ57d6KWqZ
Ez1sLfr1jfuVh5d//Pht7wH9V40kXoq1kQmSfpYWz+pu1wuC9poIVuhlsz7IwgVg
jEza5ObXO7hDW3j0PXKET1yUSV4hef1qUGFBd0VbjD4OaH1IDmXiXNkevxJQ9C0U
sGTH6g0rnOmiSFEx20HqpSP2BLct8FxubFSWVVvVIfFsvcOrtlDj/E2kQq9V8Bet
EbOb+VwzjzCXIZbtkURVbJZ5eWIU8GpApInAo2QMsm+ta5IzG/nqAWWmoe0Jbv9+
o/TY4/xYaoxGVCLlxLbu1AfBh81EdyONuEo/0MROH18poaawyDVYnywXz5arACSP
9eZF4XZh0xbh+5sDXeFsWQvAFLxzWlBbJTp53AWSrxgNufCo40NIT13fvoY7WFLY
2kZFxXFqbkRhlnjl0PV6HfPf0U80SjA1ygc04rDZdTLcBmrpBZ58hcTTu1H1fNTD
8EEEJxHx8mwS5CUnYChit3OGm/6iK1DNp4eB8N4y5k5QALS3QLEp1+s/zhX+4zwY
KqOSobiWsy4+/ldugEnwrNQXRS2rqklfTZNGp0y+BuKUg9CwUYL5zDDiD44x80iv
j7oNbJgzEnDXn3h2qdVuOAhOnRwIYItF4sCcbD9M9nJIE44MKr45XrkMKRJ9LGk/
09nYKlaCbxACMuuz3juf+agu40YWLlH/F3NupaCl187dB2mJPgg6ymt3RyMB6olu
UasNdOB0kRqteLfCw6URQOywBQB8u/0Oa4grkQzdPKZEwdZWOzkVtolxQ/dK7y4l
Nh7gMdnLNomt0LZ12xGnLJoIUCS+B7MDw+WmbYrff4TdDIu3vcqHjqDrnrgShjBC
sIXc5BpHi35mX9DqvDFxbr0iYMvI/yzl7yP8D0xn0nLceC/BdhW/dEW8q1uspu2s
pbPUPS+08ZSkcOEsk0egRiBzFsU9+uH0tUKYpVlsz0lmgI1HoTUWB0vZB/yj0Sko
3J+4UbWJjp24icwfk/vwChGDUAAYAb/P63t71N0xYTCEbDqiX5e3eO1aTQ8WlEAw
kUz9qwvIVWjx6eabmplmGilfFmDLCYgxIM+br/BLYFU24e5PaPsQGtx0w+zOa9jB
2zAfUNx/KCFfUI+fhn42yzKB3Q5PgMZa11DKIQYU2Fr7c4EqOKoodfdKNoNpKb0L
z3SqLxcPtiKq6PhLMcbkh4YI0GafSPIHtuapE3DFCDLsm0lktZKYPE6sWwU3KnHu
+uvzIVUEdmS8On/E1babl5hn48xL+/iNmPwepvd2x0AZDHbIJQPbPtM7/lS0AX2x
a4PTcRv6JqyPI9dA7BevCfG6bQDpXESzMZdDqvw2O3GOwqmSFnTwhbMLe3sZmjc0
2g1V3d1CiP0LhUp0FADaJPMuaqAyI2NB5giDL7GRGRY9eA0LqlM5JqxUkrF02i+Z
aMXWCMI1Y/QYHu5bKHklznjYbmhq/KOEBXnKbHpmgEpCQ5t+qCwyDhtORO6xlsZS
4Oyv0ZQV1JAfEEbfx+l1nvtVmod4IsA6QUnlnYYwAk8SsxqSudZd9hvYqrgcCXS3
06ieC1rYNmP4ZgRGWZOyYwTIePtM1TccklIIWjDhv8/aBVLMcdWr0uR40H8y/Irp
SG9Vdt7V7a+pGk/K+H0fY3ZDu4zjT4daSWUbs7RB1OPGw5jLTjd06vzd9efZB3lw
sA6LcrFno/CwRx1uuddYqqDREruxC/gRzZyFTf9pwTg5VVow+81Vd5kL2s6ns4p9
3uVRNSBGl3Yw9L/jN2oG91iVyiGpIW7ES+fp6A/p/3gTpbKzbuM+uMuO8pq8IHEU
TdpFqNkw+gkAeoz9oILsR0aL0eE2n2HZh/Zctu+F+WCH4IpwakV6C1UJqwogyiv0
CLBq1MCOS76BMmtEv8t06zmA6p/Af5s9w5D82jD6qBKhqVD3ZtFQzKgpGQUI43yu
LWsUIarIBMHbk6pp/g+Nj2NMqmQALHoGrRh8G7S7CrIqkXDxeKaZCT1pVnsgCN2E
OopXM820N9GQdaw6S8EUwJn8MILZjIUj9ObMj8mSlHWS8rpDX5LPukAXr6RL5t+P
i/BDDHhZOykX6w47Bl1Riukw/qTJB87fi4oZ/8RefOmRNSA2SzSHCAUNDID6KlV6
BbX2DHHyooqYsYSkCqOtDZG/18GT04gsc50HpIaflQguS3JnBTi5eq1a330e6+vd
BTndrExfs/2YUTaUkCgdlHsO3IrnIYk5LNdocC01lwxnE4zZsUw+XxF6Ar8Rr+L7
E1CZiKD45h8quCAoIIT87NLc/w1KyKlXW6mjxF/gYRZi7Le4dPFCCW2dwHf7vZFa
w/ID+yeNbPrJ41kSrEqplfCNsmRfrHv9QZQgyEnrXrEAsZh4aykaaTszjMycgvFj
iSm+sLWckyTn2RvixMWm1vImu0NsH/hpNe7ps4aN8dX0dTBQc424X5ep6waYH/DW
9c37CeQJqAEQYCKrwKkvaWCP4agMTnRvl0D6RW/tC1Axl8uqLcNZ88eSMRaUmpj3
8jX7j5NDnUkF2nwX1qxdHBP2vbdW6cIkytJmtjGs9NnXITH2P8L33L5bf6dBBwx1
UH+uP0+h2FKTXGkSoVtZfhxH2vPuphoCkKl+Olp9Uj/PBuLuF1acnFS23Q13R47W
2BzZgzBNchGJC8BVE3hoJd7anAIUAUcJ+zhz1tlF45HmX83/S4H1yTG1+gA15z3C
2qq5PmJBABUJL2DgckEoCbg911h/TTU36cZ+JMQ3Wlaexgy2YsDGnPhtSU6Yv7mp
wsRyJcGslvOH42oi8GH30b4PGFLkS8GkK9HOjAEyzFNrfqjXSKTKESHTJjL7wddC
Sydmfyo5PfCeyUHGmPtHIJoFw/7UK/CU12GgHauPTABzCv+API5+npc+445gJYSH
ByK87k5XRpfSOG23lsqoeKuD1v5tvImqckLplXZ6Dj136FLx4O96dGBpEqwPnebe
XY6pDkXveIjh5Ux1NIHzFkQ7oLnK/JTui1mqkv6z/sSYZM0JswSNpzALu0k+QpsW
nKk2Fj0Z+ZLoUiy+f//KI3kceFitpi/zwuuqD7aOHOt2qpKb2PTsIbs3eJuAnVT9
m7rg+k8TKmxY1hVXd2/zU5+sohuZwFCKtDItrq2tsn4WM0Sjcuikd6dW4TvPhvZS
yWc4cRuFHtKY4feDVr5dX6ZCmvd2UCuCOglJmPyK0AMWA8+Xd/KXrB66ekxyUiyK
sdxXYzT3sQWCmZOu7EFf6QjlqE7uw4s+VgGAL6tdXmrlMmCjKpmXkKui40CoC0W+
2UzZgxLiVuL7KUnrmEOze44W8k68BgVw5Aw7KwFYHtfjaE5lLhnHTG99vb5hlkv1
NjNdHeHYR3uIB20bPDMi1vh9TfoMhu7qP3D3VKpTkkUi6sGGEqn3FoHYRH6tOHiX
tLUmq3o4D/4KAmJvbv3/FK/pgtICEr1h0Kvd4c+kIJol40ponuuIYl4V5m3nFcUS
9gNpwOHBOYnM2lwBEkhq59m5zAypmX5XjjqKOWzECS58/BIoRSCUE6sk33En6Pg7
wESPuDI9Q6fH1zkJgZRXoGxWCQ2snkcWsXY2rJMU1IHascaIG5nWVOC/qUx/yubH
EjJoU+/5rK/ifnZKDefsFtovuhosNtr3qUBYGjZNnaNpsIl/YC7ClBeefq2n9voL
72YI9Hl6NsEV0AfeGO8YYcctQTIuLln0er+iEoarKuR2Ciy0kbPFyIVRsCRRt4hr
PiR06BMFOC4VILFONp7/OCtR4AQsnaQgfeonwyBqtXpdQcCeByPwRIVAEX7QFJrR
IrUuXIQNTv5rMZ8L9nJ6V3GJw0sjoND6vBjAYH7eFciliqwJBOOIafO+ZJakCJbu
8E9flEnyYmSHHsW38auNhk0AuqWnA16zbuI6dv7sYc2iFRT0xSNvUEyAsFzhylqY
0JxzvxpgmiywA6dSShlwYFYrE9d/j5QYqKk/NpNLdBqZ8Nlmf6n8AgQlySO0Rsa2
RywrWaal1RVQoEN+wuO1w6t8poRt1MaS6SHtWsMWk8JcwRnG8ipLy0/W4pZVs2LP
QXsR+Gp1rxMjCfUpzl8UWnMP5gsKG/UHc/1h+4C+pFpH5zPSiangPN9KrhX4UfRs
B67zttnMTx2D+H63yeXvez3potVxi0M6ssB3YJCtCCKd9O550SsRyp3PV5yx/NKW
9LQ5aE0dl6WK3BR0OXuw+rlrNjBrjbVRxgTrwZftRj8fpIyUge2LjgRCmhwGoVk9
HzWqI2GdRzzmu4JKG2WUdNFlvPnd4K3YMGU97W6q+8RTdAtDVzZpMwQMPius6E6P
gXwM4eyfxRHSnQBwR0J73pJOmpjx9XqOT54cOZyIntKPNI55CugRo+YKy7GYnbts
q+0UZjD43g5zHgNOJUvElp929OCk4H5zNF/KHmji3/gzPE6g87OeowVgUYKiSa41
HKaz0uvu7Zo9LD1Tj1UHlfQjgmAnJT4n30r5CVK4ANdtUTRjulNxSkmXIFZoXQBy
t1pEmdPvK4RF1meVQ8AdNlKZ79tINTkti4i/lB2Wwsrc+kPu7+ZTCMonTk6uPe5/
Od1GtWZZ08ryj9sBAp/IalFgQfphom5DUXXn3MMDrgevlTJBEtu1UvwI549Flns+
4hJ0/wAnd2A8J65AkLTW/ShA2HICf3hSabafdNOzYDAKxT+NBFnTK2Edb9GHVrSC
1UeuO0vt5HXVBO+yLpv6fiClWxZgH07fs9n2IrF34AcWYrMmLwV8+CBKhIHCYdOE
aOrk6DaS/XTM7gowcOZh7hQfGbddFd6ZPpykh+XmkMjpNJs3gBH6DUbL14hh++Bb
3uYuqyiUWA8PVUHogkuEx2FnvAnENG4GceUv0wGr4Bjbk2NmLTNhKiCtjTIEhNWy
uoFGWvg3TFXUunCo+GaOjS6ZrneVuRrWJn4hcgxqoCeDrAjznhGtvOQXJqWu+U85
ZcrokvJz7T+QPB38C38gFstmAKXemF2mO4R4WFXVuVxMLqJKv7VyojqBAWSCMk/B
lxLFCIHOTfHNHZXrxjGMgtBkfHpBL1jC831V1E19ji9SWMEPw0YcnV+IkPRhx+gp
y6VOI1gFhOQc2gUIGARKxrHBFF7xkMmOOSdtuSbSrEMDxk8RaEu8OICbQbPmO4hk
J7I4DcKqzQnvK5vumbIWpMIPKFyLoXLm0dKug7ZrkXH+0m8vWU9sFRyW3/27t8Xa
aMwPtqenCl0yVoXqbIvcTLM0lHpO0Rjf5UkaSwmJAKd28Eybjk24Y9cfognSF5og
oa/2MAlr08JvJxCg5d4+rUPphJ+sIVE+whtWUh3aXJ1TpmPWjdh/qr9hACUS8VOx
1NmaNwSV7VgD31/SqM4sI4JYEpxJbdHrVEfLM3aNQpXLf9KsFNgkOIZxIzERx8pu
2AXLfmg9oSxhzAqFjruDRrOEUzYIHWECPjsfMAEr1UB2krARoowwX4HZXbfztPWJ
+l8K4RUEz6MnWn/EpwtUqBJx3uarlXpSwJEd8p+1/csvs7bIf+3Sp1RU2fKnSnUw
q2FTsTIOcUVg8lCIDfaALHWhPxM3EUUoOki77JVcUOsbm0jVeBwRWUKW9b28rhVe
6TZQ1vyS/2okjDQ/uMaQR3aGeUyh1cuk2x0LS7XKpVT2E5CnBGGs1L1WVxvAYx0t
8/pGERdjeYe37xS2FvscwflX/hu8w8jpZKksGqjNhSMkIuWBv3Upmr6f+56yqArP
6uv6LrGwlVrOj0S+MuPzSDBtJiokFuJb5tb9qSkthZSUm3XNrzCq17gKmxYtaM35
hBEiEx8HOcH7qXzlDZaohYFZnCHSoS26QdCj095qfe1BfvtrrtLxSgelaa55eG6R
xp/v8DSmm086xGKpOGHBsvC4SuzH8lbUhDpP1I7V+8WuYwg1a1tN5dv2JgUOEwAs
GJCSgd+eoVPd0/4/AlouwbkJ4vObSvq3qUmXWaQ03XKs8BsAU2FTN2yNhwVPbQzq
nxIdpEvTiJvcspf9Ka3f5LOisa2ZzDro7hjoB4WFWyRKKnG8Zff9bpQMHoMSU/oC
t1OdR7JaPGRxkzwEt7Q61mk0EdDzH913BfeE/yd/ZSXV22UsM1bIr/sbE05xR+WG
EBmY8HDVV9DGtRbgile8+Akv2WKJMNqnjIxyOOVOYygb4cvimrtDQuIKDandPXoZ
O2KJNAhYxgs1w0KWNEVmP7ofksTn5cM588teCX6wXRFmPDTMTJNxLwgWyGDnu0A3
wXR7OD1KMq7cx1IxocMq3dWv8UZZXKiVkwjP+i6v380HDkm2jpC8/msN5gDpVUAq
Hr0W6fsbRxSKG0I8BzESaQ2ViJrMKdvJaxKT6ggmoHWVFsxnrP9J5LHkoqA16UTh
h821CjoZNnEhqyyVpRfly64YhuCaP+l+BoP6R/wr+NqLWjImIlZW5cNdZ1FhlcVr
UI8XhyXRow8/g8zrqx8+Lb1SyoRfGhgbH10p9DNgurER/HmVuImzusfqqlZIMuFx
bBXKcLr71h5Az6rAqj79iO0m81JpYE8THxtCsx33YBNNPEHwNFH8V0KRb1/r7uCe
EvSfn1EryGp5dKD5YvhvU6KMzErW6gAyFNmHpTSwBV+K+QHOZ2SbjgAnHa30DH9O
y+dhQG7uPn0TJCHgyuHDbqDXuoxfrxgc2ohQ2QXJaTBkkvEKIwo9siMKC4fOUq1z
Jah04UGVnXYt+bnJwFruTwrNjwHJlxXnXsCfZuqmhUbraxJuFAjNyfQtBPqMgbg9
hP2nj+2PadYQnKcIknl0ti6p17WdxGTKMOCyGjw7QVls+wwJ2+0LGdyPowhxSRcR
byMbO0oyg77360PSDWP7QS3+pd7yd/5z/slZ/+j8k/haWLOpopyCHpAdYPLM9RSR
OTc/3yUVXjfZzdlvGcUafrMAuV4aOripi+UMnucP885sjV88nCMqLTvBdDBUa3qg
dDpsbVCNan3+VzxtFxoFpZvaLxxZ7u39I4kJGzNM1oQJkOVcpHUZ8a8BPbqmlAt2
wJKXH2rqV8V8cH8xNlJx3f/c/mEWX9yzxbKUUDKvbeD90L8UNvAf/K98eHDQk2+r
5wxgkJ/40qbfs/pm4N36AkGAXOD4dPgOhlBb9PJx5MXuE+267r/2vpYZATRww7Yf
Utz0Nyc8ALnLdn6iIfx9ONBlIcsryendI6Qld04tjbHOC7BRiWROCLUmOebSpDY+
nf0L0pEvKcV0hiIUP1i1OBhnfflcbDe6QVl2bEeWR13U9gtf607jTMX1DJc2bn+J
Rj+WdfRy1YBo+CvIIPLXvjXAZ1fYrbzASoYZvqmnL/lA+JNZCV747xTQHeqCSKKu
llqzLo30qCecvoH22+54W3rS4VtMQA25GoFQslwraU6V3uzNQP7ioFk4DLExRsex
xl6oBNsmblpjv83wLB01u+RYjXgnuv3+sj9e8spAYw9j5lnNmIZdYRhY+ep/k3Yt
TSGWqp4Um0shAbuufnN73n2wZiT3qnPl6slkmmTekdGQwSC7Sj7bLkA8XcNkWrRa
Fj8wVQe5jbxwSAEnXitwZil67Bsej2yPHKSq/lmwXnCWm1V5fMBxK7ycJ6XsQQWX
2vKwj8W/P1gI3ZSYJjTmtA3u72PrqR/Xy5AONhlpNCLeB3SX+pdjgmYHrRrqq4Ya
8Dnlt1zzEmDeTqgc5Wv7g51Y25Dixy+Mv4ioxr95TWG0g06NU1k6Fx4CxDEv73OS
F9tz8UGRh39vTZx20psbWjCLq/kbfAR4OfIb5kl0qrhvVIcJFPPywTc5IlMYkqzT
xy0UVkbWod7P0MMU6MZ7rXhPgRLrYxMuLyG3H1qGW7rcv4j8za3jsCrzKQvH/7su
/22F6UMTIMVFbwtR3fYwCv+fqtbyXIh0tbrfwlplBt0MNpjI2bVziaET+8T13KF2
w9tEQYpNgfZ20OvqL0Udxp3R2Abk1H73Nq96BpPkA4QOB9wg5jVDf1HmGuF5Jq7e
uKvU/jJl4UtRxVjX+qa5YnFkLvUF0lqbbxdE+qF+3zrWXzQtB5woWyION9KTXKu7
XZ2xZ1G56mVR7VLTJLyEBf6052SqMjD0ZGJxP2N3gc6177D+6F+EgZ6D39JIpWDC
px8dcyBOKxVc7+9DADtRCtzcqexqYt9qha8SCy2KuDWhY6U/+0E3uJ4gAXy/RoG3
zjINEf8Cb/FtR3cxzqRQsLIW5axuKpQj555GJOELnRmgwVqn2mGrgJVqtLnk04wc
xUrwMMuPIPWeclZamJUbRkHTGm7if9wf2L+iPpr5LPGPVdlNKTDvLyQDLXiiHrzk
Kcufw5wwqu6U8WyRSmR1dUPoVhbCNJC/bDGep5z27VFPz08CbdP63mH1hrx8Q3rM
BNNmIMhPmg3R698lCK+YGqovr5HlXyvQMqmhSeprtBNQK4F8YMblajmluytTZ+8D
ql0F9BRklUcpII2s3ptiHr8HBk1Qut85sffJN2aCEE09esBaZ4iNqzj3kZveBv4g
1UhDY+/Ih/DFM68YUsqBehRIpbJjVpdJcRt8NbNYOhDtXEOySBke5XcgAKsYrHuC
cm6j97fHAjEo8HnI1pPN+rzuZSP/B59c4nDhPSlLm5fX5W/s51sotls1RLjx74Yy
oWfAYQ/oEdgMjPyEqk/m4x8XcgYNmg7NWtwiVkRx4dYJmXoLqnztOCIzDkee6TgB
9oBB4ZKuymZksif/CO6vf+pg3Mfx4gxVM+8Hf6HH0YxuHWQfZSYnnSwKaGCS/WG4
3MA2bw2FOYGKgsMlt4Haj7Qdzh22fkHrp7hKiIMJdKD9XhQS2Y9rGXlW2eblOB9/
RdPHnUX1PLWyMvYX7PJj6t7xTvxW0SPh7QU4R+pGxx4LNugRqQ4g5dlHoeT+pD5n
AFS5PrsfUZXGLNVIqxJ8xKyRxNuWhTZjumojzh5jS1YljvHp9GZsajY6Uyd/qhMl
vCRKqEv2bBNS+dUo/IoJajnu0AA6hDypJHL7ba2PnYq2ByBy3hTvXKzWeGPC+aGV
01C3vtht8T2ob5wlzwbNQkvsqGZA6wLntDs0FS5l/XkLLxRDHfcMJwK0Ka0cjHfA
AYpFRNTtVGF4JmkTI4ii+6J26YSE7AeB3BDYU1cx5V2/YEzFuj0HaWlz7Il7jv/A
MrPs7LouxmGrADb/a/2ILx+etCWAHFBqCgYOU7ztZ7+RRoT42f3A4pphMm0OEfBD
4KhgQw7S3Zg4bYxIGqED4Shdq/7iRn8O82M69eIFDsoO91lBCF1oy9Ksc//rWdpL
+JQyKAFSsel5ChvGsNHBx94MEZfNgQw7b+5IIFRFFKLW7HuvuD4vZvlfXkfTJPVr
5Su65XbqjlHALxjg22Hwm9GLf1m19gzdJc0wPAkm+pVW5aKIqryakjQaWtR8D86k
Q4dA3+NxMt1uvxCDWVsNn2be1UAVH+rECy+zJK5nZ/oruId5Bof5WINGULdhMWx+
b3rgrXUFxlx+irdy/EyqVflJDth1EmueFhlMnaqt0HAd8fMmnteLsoj45SePC6xJ
IRdizjgHd2GSCSxxz6NFXQ87AGRng2fS7VasLAjQVeKY4no7mbzzJedmLQ60gc0f
aXiJbaMH+5PQ5omuCgis6kU7oz299jVmHU40ZjAkVoIv8sY/upVrULpP4mhjUu/6
Wxl/TIk6zqAQ2KSzZKuUqh73u8+wgo08c3kew6ZgwZb08YZkkZcp+1lQFjsw6GUM
gFy/mKFB8w3yS5ZINYIOwOLAqfi4GodYJdSbHYSEhBRCePpy+H0atItUeAKVORjT
cDUcpTvmSozom5CQOvBjwAGVhWkwaC7ngrrG79HCPwV50F+A8j7SPrAI9Nx+hGlM
Uaq3AJtfHyNdEIo59n6P1TjVunXlpna6aHOxaWHQc9Lh2ZNkQVNY7yyFdo4LbR6B
BNR8hfDySRqD6hcGZBERfwFJ/Ikf/Bu1w0ZxmHWbyVqx90TZLLWZSqdp449oAH6P
20dc8ehBUwm/V+kLrgL3+ibr6gLQ4je/gaDX6drK41JTlvxoARTCbrsBDXriGVqO
sWRTBnMY7W2TuNYBmfop9OfobpzmpKDC9CXu8eCtdjbUoIwJ+3q7cdkWmvOCMEFz
+Xx8jd2f4JVpCOg22bQb1oxTD+WvfVvY+7VJ7Tb5wD1gY6x63DiFf6/7Bx4+V9v0
+0LOrwDIz/k7uDw6mYFTY7z4l/Wv9MiSbudyS/sOqffnGqgFBq2UWcU9u6tBz5/t
LJWn0oW7I+vLbI/TzgCX3AKT81OzIaEewQabtDemFmB6YdSt+OifjwbPOcWkigdD
vTHHiKGGw22RB5PBU1lccsXElxJ8qrbjuNZZQ2oC0Iz+dXwBFc57Lxxa6fs7nX6y
NQJW/tzzHkgFGS+CdPuf2FUuecmF9hmgMu2l5QHqb0A/CmnVpB2Isrsnj6i0nxkB
eXTt5hkSrZ6U1xHYQ3qMW99lOSqk389ZPIWXdhIM+MKj4uUY0ASMj964A5wshFh2
/0KU4kn7fUiligA8pHqIIyENckEI1TNWg7lEtyrMjA2B4ysCC6WfsQ8MoHWeBJk6
VLKxXBZCl249StsxIsqpToMThXRfGbwOq+LR0VuR94GicJRmSQi2d+ZT6C8tBdKc
PNIa/9DH20/oyyIfdhlCXfSj8tu5/5Xzy9hP50hXTCJOsTSKHffI1QWK00hz0/SX
vtrU4BjeeMXjzLYMIx8fAS62m+1elW4+eLccRBc0PT6CsJO+gZWjqBiyxlx3m9bQ
aIKOAMd/w0x8Hm9/YjVHSJUfv6Z/O7CVE7TXjD372xOm9vHGjlkvUId5lOYGCoDR
zg/GsfqASC7EPJO8NyS7mHikybv62cMzZnaybRQPk2aj+inM/dbfEUutN17oXiE7
G7T6he0nPVt81AIJ5RIX4xN1V5YvrvMAyw+RmMKRdmQINt30MSHeIy8gO0XmRwpq
+NGL3Hykwr6aEHaUo/eiPDnGZiAdAua/C8geOeiw44p5R0JpB7qU5N1CMQkg2k3q
S9pCocBi+GIYd7mpHvj4yIlQgdTmGAzQ50AegK3tIY7/BHYSpCCm6kUCiBQWQfha
Vc4TT0Q2xsuXdnQVLpwk39FKyJmFmubOXnPGPHFwQM8fik0vQrINo91ln6DlhYOu
fU+FkpyLMgDFtgCuKurJVSpE+t4iGUpLlskXTku9FmR7IhUkEZSGcGt9VejeXIMp
u2g9SjSBOW+SF2Ursd7TnFo8l5EZQtBt9S9OYv3HWPn0rWdBnAVSyWzn+XrxriR+
oye5ddTqtfBlSe7x3AKAvr2yWPJrHIWzAZrlN7Vz7Z2pfwTBszB5dKXbvYyEMOco
COoTOeQBBPDzCS80QtBaFlklsRTcLZfZrX1/TCRdfxQ4iXZs2AE2F4A1BDU7CkHb
A22u/BURCj5AFJ473+DEI7l/1P7m2i55o6qaPjqzk/n4hxQnt0wKMyreWBqWrDvD
Oxf/fAMBld0iXVeddQDEc5s6yvjC4wgXW9s6r0+OdJA3kcCzkKIjV6fDa7p01ZM9
lv2GgVbjGPoh2M7D/tsGzZkzrEjjTROteF1EXHk/TaPWQGDS/i8uGw+W+yv+kijD
Ra4leDJkSjG2ZzQkWnHk6imf274wUiOvXb3wmh9/yRSkXDAgOTfztQFke9vdakB+
La4Gz2Do+6sNj0vhGeNaUidUVF4owMVoWt9pPAahIpWNwTE8miOZsnc8sd1xxeji
n71QaP/jyjEyzoGnu/nLAgORruJdClBhLc0wTWZ+YWBJBiNk5Ja2ToFNFBBmPgNq
jZnODJRiDHmTLlOM2j+UyAFW52egYZtfbB/LskKZmSy7ml8GQIGwphy2jMNtUmJx
RD6nvFmjABZuTvJOxvGRsCZqSfhl7vM+8PwLqmCzkwNURjUjvId2w5IbZjE37zky
jdW6/0+ppDM9/bJDhfg+evwllsHfqBls5Q/tRvmAXSoXBGv2umhkH54lt3wfKXMk
lpuuCFgqeQO+1l4z0roeVmwYW9ZBpz5UORrrVo2Lqlb+iXNYtE9uLNsvMTSq8RdS
ZvwcID1bjMFMwegwPf0PY1z+WFBH7CKDmzqjMUcGuBA8xAwfZga7yUTu50hC1sDG
1Ar//jUp7w8eundKEWXhwP8RbqkYQcr2kG0JYjogrr7r+LXEpNV6U71yX78QFm13
fjP0eEswIzL/A7SFAAB03PWEZV67BWUWDP/Eryru/qj2VFzqvHzu0k3IvZAeqPRL
QBUvKoRsro8pToKU2aXBTW8UPWVzf9YpRm4PQMcbJWoSe7V5wDTXYCkrzNZFh//V
c3hPESyu30x94s5h8plvXX23RxqubmZhVaGxz0adfu2zmf23nEv+a7CEs7a8tg0n
N0WnL35YkUj2+imQHzbSsJKmABkUowfD/JhRh9COxRK6vYSuW2KkJNI/UzwKz+EA
mkeRS+tRbLZww0yXXQy5W8pk2/jOhVQZMPHhj12Ig2bLOG75O44D338jz4LNua2I
HYtB81TJXdnrj9554zJxeaKXWtZxJOzwYv9FYmBm9dsdVzCrmL5FV8wkS1dJwUh+
38cHAaelKsVFOyzPQTkw7vUKFH3QjqfynqT+PstpbhCAB3ahl8WqgqsN6Cj8QHM4
YztcGwm3PAPaHdjO3I4oD7AImCbfMOkcaKYoK5Dp2wHwpHEEEz4XkFz0wEMMxeb/
Ft26IpsB9QifDPgOrZXZ/Tes+2w4NiaaGFOqkd4+PwOk+I0ReDZwvRWZmCB8L0NP
52Oxl758LssL6umLm5nWlnOOjLADfBXQc7hRk1CrKn+X08P/nEixiENLSacpA8dE
XqQwaBxD1z7l9Ootfsxw7MSNnNrMQmaVYcgF8RQ8C6aVpJ7LFEQVvE8ePSN1AHbi
GrOYgiEDD8Fi6Sc2yvw/YMafR0JqJVjp8Tx8xHgzrinhwX4h1IIXn6GwWrhMtsrA
HlE7TPbq08WNMPAiNarWiq6W4v/B+lH8sg3an2CNkaT7E0QDvwpjRvZyVgsZJsIt
yg7K+xJtdwmEgbQ48LftfzEOK52/um1qba1IF1cdCl4XpsAE14wZ4yz+3ncL7xG+
+kklR0ZR+5iLUHptoR9eDVnHtB4vmb/IDWzfM3dySnAW6FTl0kUjD++rLEvO3v37
lEn9rcWHKsj8khWeLMVc9FhStQ63DueV/XbeQ8LMAtkVb/Rw1s8daU8HP9liypSR
SHMfKiSTr/5APIMhVUjgy2gLmvw0hzKbjQfUa76G1k1SWaMs4AHVghTMPSE2HW1n
MFuPCRPbKZO9rD+eEOu3KAq5rK2pAFeS/OIjDuXIPTJterKRShrRljC+zxa9ywne
QLvCUCIdJafW7QAsFLbboBRyPeRZIbbp2OLzlRi7UA32Qxd7+wG6BqRV07mN4JrD
t2sV2wjzuuj6RuhYkUvLuskUeDGPelI4zj7PH2v3CaXGqZ50IzA98qWNjLQGXomX
EFtKDqwjnyqytK+k19REXKJjZPV92Hph14bbopm7ZOPOMCHBDbIuk2ZlMiH4OQ4o
3fwXynxHO4A/LgKGLBB/T9q3X1dhKWLwSodvknVLIK1uGp5VC27p38dJHvDItWy3
B5sdeMx9WzAZQagsIQ8EP6qTiwyxsiMXvpWuWhJR41d8+9tKly6yN8A0XGDTQy78
0YRkYTVKxVS8uqdJ+QfVJ/gGO+/+JTOXmcJBYQAFlOfY7Wh+iE1ulWtPfiygOJtB
UDo05uRcZTFExY7FF+oWq+KQk+YVaNA7u4VRofdaF66Yufs9JgrSenEUSU2A5cMh
FNwo2epENRwcud0+ySixRIFmUThRUXt1qTWwu8vj64i1YYhFUHQZTkjghOdLm5rB
JYStANQsB4oBr3iuoqLigT4f4oGto1sE3vZnfGm9w8XeVrwklNkxf61HT1UEUyad
oiTGJLgAESP9bzcKbOs3vWHK76ykoJA1GG8hw1HElI9EQr08lJXn19eD9Cdbrj81
DiLb0AU3PpPZO/NU5WpdvpOWsiNlFRWP4Zm3O9HxoFROxvbpswvEJ1V5CHUagubD
V8NIirQh5j98VJF2ua0XMkJ0jOiLM8s1aAbfIvTnhoOaQ4cSKZze5d1FENy4SD9W
pI31r0eVgRa/LclyKRGGNXjKkwp05s4yd+nQhEmi0b4sg+0+mSYWGk4MEk06BytP
j4L/C4Kn+HuX970lMOct6FuOdm0BNKyCoYDSk9HJ9/D+IroMEcLSeGwl09aZIdwp
5tLR0skLnyqTMYiWpRS91ImdMUM4TNgfgAL2d0+wsZ9VpIC6fPFZ2k0YmI9XLTzv
pEbAQETpRsFtcWrxucHl6j0P42UJ7ntMBD6XNQq2X6qsojAPzrrE6JqsLJCkAcER
scUzedlwZl2cWvN5vsKPULm+V+6u38Vd10pexwxPzdMJFzIGY+tkncnTj3/VcESl
c8fy4ps9v61YGjk1YRo+3d9GyJEDMS6prFrlWgHf5/K8kgMIYKrTxMGitVtIGPxh
Neu3dsPJ826kT5XumtBjbmOhA52TWLwkpfUwL3/TUp7bvzxJyy3aWvUH1Ks4m5Xi
fHrL5PzCt080DbBurBa21ZzY2GFcXoAJBzUDvTqDok+LXtDLvO8towFQuT09f6nW
NWdj9Hf7f9xSLVKZIbzgiDQskWJK3SojmPMnYD8wAxmUNbtfBol77DRWvGDV+llv
eeSLP/kHAd/uLMjR2QgqJja1AT1wtxc8/CI3NUG6SiTfjA9/M5TDNEgOiODslRMj
wIe6aYpjmuCV9gEBsleK7xNTmdhHSzvK4MUyZ750jHYNB3kHH3rw7A3xhIsRcbkG
2PZiADDBJe5BPbbzPe31yjszweTxyaIjvOlfUmqEKctYmtzjETY7vTF4D2N0Qmca
W+mwMD+ehWn3l1/dt9PIpwzLEDgIeTfSI+hVXNFaGRApG8sFVGamWuD46RS5RoEx
Z5CAAepsiXRIfBCuY+MGZGWuTmApbaGId2oPnzwfh1zIFgWmmics9VrT5WriLszi
itqkZxJE2nyma1e6If1RGUgYBWTi3lezIqG7IAdbQxwX5K6h1N4zjKw4hC+E9BJr
w5P5XdaGguu7i6TAs8kqwdORBd7G7NUl3tCSWVOniwsh9m3efLSdpPUCa4GCv0EF
x590WiFU10p/10xcCkuKuX39qUkRSWJSBcZfP5K8PUWvbL3nCz31og5RF5tKCUQN
5TANYpUv0fUbwzt/e3ONDuStnp8y4Rg7ynjiwzzchE/FBWvcnRo8EfDEkF3OIxDm
To02qUmor5Ras4GKiNDKQ+CL5STQOyUQ+kvvP6lan0JSWNJFnlXyr4IxpO6aTF+i
MVLlNXuvpn7zGf7lHpgOGTSXMZTyik+IxaX8cyQuvKWGdeytXXbD5YaXRKuQT6q/
6JU5ay5f5fg/PhhQ9PB7xp6YD3jRov/JunEsk0+XQ0HUyjl/HQnabYQ/NgrntH71
uYCenAK8GjrQL00bb1Kv9nVD1yCclpNdHwC1vs0siSzDuMVNOlnpSHyrHJzNee5a
RY7mbcDjFLo/ksW8a0YAL+EhyTDW5ur9g4aItyTiXVngZjaRW33EeH+p1mlREJwb
m98YQDYbN9EFJ+sKKeVVGiPqVttsI5IeJq+cO0QcbfIXtcsKBu3YQ6lROE90N9eo
6lGiliZw2CKNm8U+06bA++SZeYVrcHxIlgsVi8KGoEtsGr9tKHecj1hr1WYvEIqb
/Npp3rZxFs4N+NM37xGsa7QQKwAfExySXque05NUsFpTYmsoMKLMnSUKTMRNZUUl
ayUnDFVw+YqKRS8k2AM5SjLWWIoPGYIwlFq/BigjSJvjPwpnhrJ+XaQKaMmwmTof
TsLuzkzI/aHHeXjap58l7mTsgZAF96ZXQ5qkoEZO9W2s5aOi/Si3Zm7R0vEd3bHd
86HAXDA9785/wvE7BZqUErf4m3SYgFptL4wOucUemMaYR6Inp07+ZuFHM7vdoX2u
cmGTCeqIiXRKd/ERJqOax2gV9BB7DIqwEg4fCRQQLw+V7uaFIQR4Bz4xzW2imPl/
Mo7DOyllLhsutWvT+LBckPr5acd5nBXX0/ATfMCAebOgekLpneUpOm7tAKMJ9cLb
JQTBZ2Sp49i5dgh3qgp83b9W9bMfgz1NuvpzDykxMtu26YBxhs0QBQRsl4aR71EQ
EeFeGFlUl0Al3d5NuidsUUq4TWiGIBiU/0ei1JEVVBhGRL5HELdwk5Hz56wrxmjl
VbD3yDxx3AP/xvNuNesfwwJsOdygEX7iygYIPhAz+hFlEoI7rTGt+B3oVFceNVW7
SOx9me7GXEEq1z3NhEe2WBXlL1E4pXaCg0vi5EUoXk8Lb5uAAqwvFQn6IRJQXzBV
7S2eXlCp75LSMlCQpgFGdA4pBWK6xuHSInkdNjaA4VqokZPAnJI9D6iYmbRIlpgm
oJmzA73usVaReFWRoWjw0+4IWcnZVjif8o2XWz8QHBx9fNENz/3bBKzewg393MSV
yWQFx4i04eIo3cPZvQepsCkNJnoWdY/pY8RIyK581IVXBH83V1Fr47MpjO//Kq3S
PoJw0pb+bUWdstcVqa7fljFAerbdfo+1uY8OBYduOJ8AJeN96Ra1Oqinfd6gy47S
nKTw/jEf6Olkc0TdQ7bE9+d/yUoNRL5T5/fckmQ09LAWlbewANyRU7bKpwCSW3Bf
P0IL7n1Xeop/DIeOo4jNmX0HBJShA0b8QcxcmP5HwqzlB2Mbu01K6E/BofzV05lV
ekjmjPsVLPz3cKOa9ILUDoaBQA38FZkdGy+3otaIg/tw7rDIOaBsFTMj5yFB5mey
wsex8xzOVc6PdQVaROLIkYpYCpro7g2HOP6I1QSutOpt8mZnlYJXk9ULt+dqNWCW
2Sct0H9JQM0f1xVdnme8G7+ljU4hDnTCIkyGt/mcpjTlJ6oIVSAvNDDltc9uUIQX
U3EGzRa4/vkHOHBSu065i1WD4s6igRgNSTKHXoLdWh5eLD2vv1F73G5/n5k3FS6z
i0mR+u8z2p1OkkFYZ/ahTTx61qnLYEXeLGZd2jEmzOWoqIPZB49yDV9BEyc5ims1
upZGP+eb0mvtngOslNJFTfdazhwRGQ+cTLel/Zyc6YG1ulv5tN8/Co8TvTsi1AEc
sBmbO7uSh80zZ7PwkvRGrCRJCCximCotvY1ZjM9D64VG48uD2uj0a9o20azO3f6s
zZSSD7+M9IZgnFG2FyS2vLeP5O+eYXQpk8wGQgbeoOpiknZOJr+/q8b3vgaa5Vo1
J0eZjXz8Rl0uTXTMUZhTNLKScCGyKO4H4r5oMlbdn8b6L0PZtFFd9gwUbQDyCkdo
I3bshhKbX9Kvn3SSpzsmluuCqzxu2tvA6uiT8F744B8ss3wC4YmqLVrLjOfr/Kjp
QvKxyBJPiWf4jTAtNT8t01CUzeLODCayPePjjLT/WH9CCDihdwaA6Uvkq5aBjGHd
2x5h/7eqm5ETskRMeV/B+dmELORjIlPPQWIOXgHhS7OgZHNLD/NDIxvMI/Mzkq9O
PzGik15ri3flojwmdrnR1hSxw0+jkb8vpw2ffkujbEVCg1VADG5aafGRxir+RI71
G2/PLQDfeXj/FkjVkWLcrj+eX5Dg7KxjUSQ2meIA6Vpt2DZpz0KOC3et0EdeiDZ4
x0pR5Fgw5GDW4NSkmfcxT94ot9hedPtvCUMPoHm6dHQccFZktdFFU3JOfIbbyDbx
AAxtgHye5/8IB4YTTIdkvkPdz8w1QwAtpFXDFWO+WHR+gYl5wND7QwP2yI/REttc
BpDfIon7jUotr3tebRu0rq8LG9rRr6LF6tuchohRFeW0BoIshwpgfMRfO3V8WK0F
hXBt9ut0P6Pt4xrDLQiGHLGNLNAntXUH6BwfCS8G68jmVymEurMcGFWyp71zmqfy
Z/qfoUPhPi8OJEM1hIbXTLxKx4qKZ71BSa+qGP+K/th/tvxzUtAm2TgHI2TR0HaX
KaHTo0TzFmDF2eJoyO6aQ76KQznZUGPsKP+VHPExWazz4lZQlqezvBa3YKBwls+i
nvRrwl2Kh0HthW9Q/mfdtQo+lgI4F68Io7sxnzDZnqtoSNLZtoJw16C8ygOLvTvG
07Shu6m4+3/7yF+PARVdzrdQfj0F7gKxUPuvKQZeZWXkowRacU96AERaa648hHyD
BoCXCZZIehgaLriDQS8x+d16gW2xR08VghHp7Uz5ckHPizWtHcirk24wOAfRLL/g
eVUML6/AUssk1Cp7QUzCjzehn2WjmqLp/78iIektosrFoyeL8ppO+r4BBDYz2+qH
2phvdsjBqkg/4XVQwlhDFemdRMCrATAtUEObIO0vnJXn4AwcB5meb0VO25ZHxgtv
MvAKfzYtedU68k02XNgUArHwWraHF7/YCufP0T/z2GE3tiWy/piyXNKw2RirN0W/
U5oWIRHMqc9uov3X7nu/FTwwDrc2/ILhmlRaD44xqYcwJlbFgJ0Uwt52CBu9uPO4
bDicT+P6EaiTC1qSA4j00m4JszSCUixic8gpzPvuaXq4jzYNi/uwFYXHirSWdUOq
AQvPCtA7Ke3k0fmHz6zBWz44k4Te/jaPXKkgYUcBq3Wrnm7qRlsJiG1W5FQ56UTn
v7Mrl24krylzPb8gcnYpuvcOJeVXMzRJMO8rY/LL5sOJ4oZ7xeyBzssGtjh+aMP9
NPT6FytAjTKPXkTFH1Jsr5KhUFzBtSFG9Qx1er8E19CUBky/xWXJbfnaz5jrjj6r
c9C47LIJTci/mpB/0Ut1n+xLFxmyj65bqmsWSizCFUs5sxUhhbtZe5f8BLDhtb/l
VBik6TIURZKm554xGfuN5MMjAKshoGQhrQCGlyh9cUywv72kPnZ7NlIHFvWPC9t5
+W5wVB6HVjs/+XMqA01FdhnM6igt8wLEpu1dJ8halnobtIYOnhojPCxNqWwQzE3w
Cjj5io06eDh63/kUvFRgkE2X8+CdcL37ti3eIWxBDDKR8ytcP1sXeoIdu+6Slk0r
ConkuTkeogsYwvt0z7Nb5icLyvXygD9mSc2ruw4zKtHWA/UwfB6AR9TP8KCRL+bv
jJ4oWLbfxAJbegDb3WtfD0jldYmmb7IGh+oOIIil8uilJMD9wk1e+2JH8Plxm3v2
8uQJYz0rSmcnn+28OX5aU6Qc5RBfKDIKeX1Pn7iNr9kVy9V1ep8zOaAP6int0O9I
3jsG2aZ6g0dLLXLRFW6Zuj82A1zceIhjrsDGcd6WkqnXLOZNbv4Do5u4j2lrGcg5
Fu4noh3bZ5VUSR93fm3+h9zKP05BszWXMnYVfHhAMZHllHu+LAw4AsMVksx3XOlP
SE+VotICnyeYZJvfzkei8QTu5VNibWxANl7dL7hBRTDpU0ay4wE6rXPm86ZT1udw
o6BztmOALl9UxtfSinRMgReG4VeYIXmvtetBWSykszBWbCXw2ODRi21pPJ0d4g1O
jiQQutRmCKoIryVZL02H0FRFwztyBsAHHLdEHrNlgyRu4yZEcS2ATpsVI/CPDH6m
cVgD/OGRsc91RmfbZEPyCEDcdW7UBlmxjGwuEGAO6a/Sz0n4c3DZrd7d3Cg1l6Pc
p4F6sxrcQ/dM0n4IxkrcnjpIIFsDpWOGhLwJcZUZucxvUjcRgcidrrFX8eWLpqLe
FY9MCQk5e+zq8uQYGn8DXbCoAdEz0KmQv0+vaV9ykqZvBbffP54ru8Kqi130EWZ7
jHJmQBIl3BTz3u63vTeq/gvylG5h82e4FIWUMiMILsbk2LBKnOks4/HatoCkyXKa
oKtigDZ5fzXoXVas7SVxT94kLEM1thV70sA5OmmKQERZV9+aPka2d9EAusYMOz8u
Tj8K41v8l5VJ+B9jexmvGPjs0oALCqwDY1iw1sP1JEDv0bwLPOnGK+7H+ybHO4dJ
yL/UQfrPIWwfaluAy95oS8OGCRTOKBWTzcKSqS5B9Lv3wRU3Geq0+bsoxNRGkopF
oI6UeXwgYbq8sIuFTo6AceXMUNnu4Frmikh4/eyljoOyFrwxNo+lMXTv1gwIq2X7
1Dog9bU+vF+/+MtYXeTAu61zhkZ+bRoX1Dprd1+Juptm6vKG1yFX70AeuBnDiWfk
mcDpZEPHIhIozItF3xZNB8fjvibSWxI+mHRRR+dajhT1KJsfhzCnwBxt6NeCbkq2
d2QtvNMoEhOB04mKNrAPUYQ+D7MUfkGpKCsSxEBcaLSmjhzg/3rkInQSfHp5tOoH
G+35aVix3kD4/MVtVlQrteHZjoc6+ntlSQO54MH6q5QP0T8dCfuQKuX0piqWg+Nc
XkyVKi2Q2gLOsBrXQyfDt9TOPJQ89ihy79Q3UfPL3jgskSyZtuVhDXxmcb0ZcyUO
d7021edv9SCTDgNWQnsjyzEf1QXlTycZIIslcdNlkgUJKxEDjX5b6CNLJp261md7
6yeSR6fSll21eoq3v0kedvhB1YvJQeppDxyhbn9/qbKkvfNNr7xcoC8VF0/0CAz3
mJj4WCls2+HCMzDHF7FRhFkLjlwLvDbNnnch8/7PtLzCHOZ73HHlCH/P/d4v5HI6
vjQ3rVmsTw5Sqp7qvL25i50ZpOWsJls39xpOWMBX3sbBiSniBUGtZRP8p10YcPxr
dm3ti4o4y/DtnIKEpzkCXn4NXgxXOgKoBNOXreZ8z6PEXBpJ225kMaWWNG+qhBkc
evcZj2q/6f3I91I7+eCmKoveywS1OdN+Ir1glyleaMlSXHUyBO965wPJjFde/cIq
9nBIxiUPV8YB0rM9Zpd+81anATDoKdg7fpyDhbC9gSCQHNuDCEuy1OoPY9Xuidlk
+66zR6T+1T6ngIWnS/mUPcDYS/H9OlQM3U0QsGnbDnTKVBuYGYYMv8BQmtnABsXg
vG69lxSiax//pktKi4pPZ1BJi0yJgd1zET9424NZkiPD7zgaFI+PmI/htVRwAhud
nKDdXfO2vJgKZqLN3Ku6f0hsJxdin7ot1qiUGmSsbSatyVfITB5AZkBPUT79oqnU
S3T7PEno4MDFOdArOPlRvb/R9glKgHbu1TVyvMEZxI3sRkG1m4o+wzAEuq9ZrTf7
4pseIzzW6fScrrj2t7ANLe4b4IPZd0YUtcrtR+rgpHZPhIAuXWhizCaoJiJL/fAy
QmC6G/nubjKMxSnNI/CsL+21j5W/RDPV0P3gM99OdKi2J7S4Nur+8AGNM5UjTOQ5
OJe7+7IbIjbDB6kpDo0FkEfD4entmfx35XOGAkuSzWFRJHUtwqS21wm2I6+Wz1+6
9v0/hebXbDCPDw4HfPqm6/ecNd3ufQsXtzjehXkXfZmAIttOc6Ca6j8Fdl12mg5t
IQaof55eCkfgGQjW1yLuo0NplpKgmUnatulzlvANzgAi+vpkEdQNix1gMvzSZaf2
f7upyE6Cv/+RHH/viV987XIfp/gMnrZmQMYl3vDnHIfF5SEnh2ezo7vVRLk4Q2Cr
txmkWzEBBWnJ5mIjz8/MT47xfv1R20u361xguxoP39i5zu/Xvnln42B7FX+xll4E
4uQjw5h8BLntwX8mF5na1SyS4UyUhEZdWt9bP8j/4TzygSDyZjyRIkSKIzeQpj74
u+V+ItyP99qEkogYpYYJTvW1+N1RoSFWon44FReghdEix5yZY+KarXP+CZhyxxwr
Qf8TTOtKKNKbqje5Nn94IfQ774WOtJaYhmRfwzk3ussaLaTQ/dJrnJiPosgRhLi1
jFx3qz2TLDfqhhC8QqStVcRZpLGBgy1eM+I8zfahjRDcDoE7wvPOm/BtGvoY/Pa4
68u5TSFvnj3AWE9WRl3vN3ueeN/SZuDc3x1Svn76ucTipfUxTX4EC8ACcML+mm3L
vABMk4M63d/aV9OEwczThmcgCk+AHjlHx7Qn5aQuqcr8c9cKzVHr0RypiX7/o+GS
zNuKtx7VdY6qWQ9gESXjs3ommIa1sO4a1JUCG8gXv+PA7ZsaQuyPIaBkDI1EdBt+
ITMMrdGbUQ5xpyOtfgFpi51DsJxhxEWHsCJ8KHBWM/QKz7yHWBZITGe3BqEnXMuc
HTaj8BXTQHQCgdoX8eUeAae8DUHPMGNc+UU30Jcs93bJnaggsWfDzBOm777MYb+8
5z1RckzcKRMo5TXSv5IwKdlmZhvA8GyRRJbt7wN2TtYftLiNgoYsZR9K/ClDEk91
JIxURnDpAjkNDxSX4/DHh21zG29SLFtZ4rHdJmaRIR/cYdEyHsLSzfMqorKolD4D
ygYpHz5a/ZrIBgrg1xFN2zHdsh67gvJ/8T8PAIwB0lr3WvaGpMMPHKNV+VP3B+XW
SLB9Rqr8M1PlxzOigYyqjm8tai7n/O9sGvDCzkNes9DMx7xqBy2243AP6jzzyGUP
nOLWoJkRCNFpat88jM1aBY9HCp3QYDlO4YbZAtF+r02NYP/Qr+/I1opvv5SC2XLs
kHSmJf8ylFaloP3FS93gefr5LDrGj0ydglPtn9ncKAbnkXJYylPu4v287gYS6BNS
zB3w98bCd92BJFCXgWdoOjTfrnmRxE8lY8oBqSTx0chKljVWmr7cEOrBfbxWc77f
0HbbmupRqh8lRqCh1AVSWF6CjvkGDSjIi15DbuzejsRplHPua+ghXYjrx+nGv5T6
7IBpJ9uQvB7eV6DgpN5kxHLQ+0fqnocRXxdEX5R5ZldRVzOEpqiPihN2HmmiDCWx
RPwceQ3JcQ7hfM3gWjJGLEw/rIGZUioBFf9HoIh5chjF5cAlCpNHis8X71/52lgv
hlzurpdKDyvUAj2Ybr5EB8cbaXKPLncqbGijfaGlR7LGHPC4xtoX7EIxtN+jjyR+
j/zUDGYnozo41m7nBWVIWm0fQJnT0zbZSfYmRrW4GMRKuC7RKERiRs86vUTDWTcf
Q/UPBRZxI29e3e8IthWxU9TYNGmSAF/c43aIisAMDyz1UvWxKC2zxHEltfPebFxV
msKy0yftlRuuCucgja4FL6uo8diswoPvZjJKPz/Bp5vZuxLjsedovhZ52WfUnRNP
l3YTea88merQbLHqREAAVEvnQVUl9T4onBHYHAXoDViYDUiozfF6TaK9whizJeu+
4UNtzr0O/7xx6wIQkTu/WHHEniQdqASsF+d8B/QOuUGB0ZKcpGE7/b6wJ6fcyfEt
jbOd6uz/XrxgYL2Rq8ia2wtxUpN+B498dtgq0xDul/PxiqKnF4C7XYq5o8Bw1YaB
XohK8F8Fs9OqRVs/T2V2syjGsbQj7ueOBiYu9d4xC/85HRZLpwMkUTeSuEjs1Bjx
y+JB+9WfjfjLKgmtrLqFhbILs/B03EZ0wsxg5ulyBSQExNQ0q9H6on7YGYIeptw8
LfewyKK+mTWDRg6mh2wWiT/erE6heRuVjw7CABOw7QP0Nv1uDdJPbDeRqRyL/D7g
YsfsWezQe9Czj2NlOFcXkO4SEP1AvFFCI/pugjpyTj/NF2p18T8YcmnKgoQKyAVY
6P0Hj0ZZJWsJkle5loQRdrUNrU/uV6phlxO4eUNw84YIwSJi2TwsA6jE5t3rLIIt
RoQ7do0UMwodBEb4QvfXqe0SYlMv5eLgHJH4atLLUhDN7fr2e+mceF0U2JrP7qVp
V6GylqglKiIXregxoditR9LTRvVT+0zEdDZWwa0kj7ZEDB5Jv8t7oJEbuz1LpR86
SHDwqOT7I9+YiDwLBH7X1iq7n3l6rgCcY9A7qb3FvnZZyJvB0RofkzNqJSAgxF4g
hrP9e1T9Co8KOFF1mbVJwbJn2FH54WLxcyydwfOMAYfwPHMKlkZhUW4Kh8h8i1gV
J3v2koTlCZt4qEM0a8hdm/Da6l2a+yp8SqpQlvk7tNwiGgL587vUN0WRnGgt6LCy
6saAikgKMxsjZ2xIdT6gkFpdJQsNDkMilb23TncYASZ3kD2wzolnj1QYF+ARMk7g
UxWTj6wGPMaOlqMYDweT77kUoOf1LkiYgIEz3Jz+fjXhgKB04ib5BO70wRLZLXEq
4GIwlF9TNaqoAdxwV2lLcXGUZMCwZLwEgxhSuTQTPuC2EUJcNEfhpe8akQ1XY0VJ
gA9FZ1vpT0L3uAmv7sYDLKwKKQUVuhARyArBvv3d2ydr2eRbo3lVW7c83u4tCoPV
/aGZseHF3pCB+K9t0cWdkiU/o1E2wYYFzTgTf2z0Vvtsp9vJZgMS3q7IwG9SbpDU
NuWOoqcaa145/qlr4JwBHvjhrogcRnppzrD6Z0OQ6rEu4jo5sA16CO0e7GUyJyp1
/LFQ5tHBrTR1AJjxBpeZaLAxTMkg++I6h2REOhmq0nD7HiNkOK1Yq7rq4QLq1gOj
FGMpuhm28nGsvESgWbD4qeGmS0eFb6KwwotmzkFfNIOO8r+VbEejRnhJPYMUTssV
X76Hu/7KH8XLbqHcFsNUUxr7ldh3hVtccZs+t07c1EZHdrX9hIJ4gQlw40BdGvD+
g5uiIqrAdgyqmveixOeRNooHWFXhxyTqstrOEDmDEKus5Bzi6UxYFPgE5Bl1oLhf
QISfoIxoN/aCrRL1dMmiYCaKCeKtFzAxXipHoeUlNgIjJRq32NYyf4BNxIx+R8cP
Nphc3gEXSPQzogM5m27tpqCJVRWsxGkU4UUsT4L4+6yAaL5gD48SycAeFExFR9YG
V6ZsprIi1idc7SCk7IAmNBv64egAhN5QUm9rdeEWoezpTL15FiKn32yWpjeED3Wq
SOnQeC/7Ao9a6Wj0T/8PlEgyfIvaMPMIKscapw/GNFhJXDwn+z05z3G7hibFn0+O
fuxE/BYvAzVe/Y17zE+uU3hcOBVcOzFRtaRbZVlFoj2wH75qkj9bsI+NWA/3eWGM
1zYmGfOSc3isi5SCJCdTUWoc1CZKBbomKIHkdIXQYqI3ZvJVQq34Lq9Llc6si2eC
4capvbysxxUlO/sfap8Sb2oyymWuc9nRzc342YqWmsZEOyBA3MP1KSTQGkcBJAoA
H/R8wqnfe/Ik+NXrE70kFrEQ5ENQyj0navkP5JJV2lfP+ag3mfkPE7idJscaoPcF
Cfuu+h9GyDnuGSiUC67QyvgRQ3iXAXq0Hz021w9Ci6bKefpqLVKhV+IF9iwGgfoQ
KUNVbPDwRt+8YSy0ePczzV87aJn7iqILhoQv5HjVDI9m2DzGv++dWspG/MFebaNl
/PCuh4huGCVY1JIvU+9wI4FZbdF5Ps+hcjrbn8AGkwnXfXkL8o0zSR6gk6CbUoDX
sQ1cMsIkvSF9+LhEFdWDj111Wq1GZJrjPflQLzYAEpdhGvLB+C+Per7Q6pat1luC
27KacPLKZMr1/2oSXDe0QDxD5iLZ7FUT9HublRaYcJumw8l6GVjwAdGyw6SHnMeh
Iyg9q6FxMuVKDxD87PBKVTRFugC8+uZyQmBsSbQ9WROX9vxmL3BUtdbEyddt/M3q
zq7kL0iCELHqUzWdWeg1L1O3210LnxO11FQfZTklXxF5UxVDVtJqO3e4EXnWJPCc
HEx53CrZOKmH9F6OhtmDeXJIYGAKMoCzvC+kBbYknk2Fzer21g/P8STfhFfaz404
eL9EzMeeCz09RlB2JZx/iya4io7ueU4YRXH/XTfjpF7cGGPb7bZXMfCQE8tMv/6j
WLkMBO7Qu83U9a3IjiiA7r27tIP5Ux3Q7D53YsL55lkj+TbDsXj9jvXcits836y2
sBgq6yMokmOGXJsix0KOjBnrGaTekDuOr8Eh+08rwKBKAGz5Tpo8s7L4Ndk+o0L5
Hm3RwZIsujRik4dMM2UhCKegFE965GFH9eJZgR2VZZKhNy8yT1nTV8UM08U3meeA
Uuyg5i8HryMjJrzgZL7bc6dFlMBF5mVDttGG1TTdWN8ynb6ry0g6MXb08Q5Z+nLX
3gLVmFDXbQbQW3J18UseG+jUA6KW+0+cF/oNgh9q+XH+uZGCYKOet7MwsnKc7Voz
MnHdkV1D+/E1isKSlt0ADYtSCnzOSXuJOPDViWaQSHoJNZ30wApiGiRewKG56796
Ue9IlKZE7Z4/3n/qD1wyuCqIePmQyoiv/AOgGiUSsH46qNtuDLed4aMGvJDinYsY
3EVBIpRitVcVkw8ENxnpTb5O/9AyGFfqECGW7BxLYP0EQTnOa92QLi2pHI6elNRb
Grbw49GyR2nLKTcpDgaGWmW8qjppm/EKxilYm7Mk+Mn5i3kbm7zrJSywsDXX/OfC
dwTvtojGdM5a3OMs96OQKjHRVBCKeZcQyyiL/kow5XTfNnGA46cf9rOPHPEb+xDg
YQpR/Vwsiall/u8RhpP9ho6XyyeQqK2kBdxxdaVICv/xMA8O2Pq6/B1hiOCqOn+V
rq+WJEd0tCMu2ur3c9LmqTGjmlrzLcn/3j54KuP/uwQ/a2i3m0nnKyBA29s9L87t
fkOjKLmxpQIZKRw8Ff/5gEoZiY7jYW//eWFEkbl3I1vgrbOWSnVKDUiX521eCH9B
Z4UndZ/4II9scCwJs+F04HTUAo1CDQoGoH/n3CwpLq2RF5YM0YHdEki8aI9EPrsu
cCS+4P3IoyCqEta0U+jltojmBZMkmYlZjk12tzfsLEKQUfVayI7DBIHFLxxqGJ+j
yTETmL0xGrqfvP/OiWOq6/1pbCyQccS43XR6ze5tatEYfAsquHcqPExe/lRtk0ke
w3TOEp+G5rL41Cq1xCHGDFCKCQlL1P2OIR5ciieHL7/hbHyBbhHGHWJNaPdch0ow
uCAScbVuxlN7OZtTfAJ/kaH71qiJ2EtysyOXv71dDvM5xlGrHUC3FYpM9S0OaU+U
XTTExpm5fbAU5H4FZ7q22hXcof/x6GjFo436q0FIZlgSNqKYrbhGWlmLBAbSKV4Y
zoho1PjDPyiv8VnTjlAjUWbi9UfCetURIT5PoBDLNml4FfgCcGqFazyX4CAcvrXy
6xFV4XC9sS3E4VjDczWkFRQnFaIERaKKBdUGtBcazqdduWmyLF0ywVmWTQq2k/BS
4ZaRasBAO9VMo6UPjQBe/Y1jzw3XPpbt58nBpk07Y2FO2WLF5eR//T/Kh9rVO8ef
Yte6lOYZ+6Ct/F2GrbcZDw2hrCCjkapXT3LcFrHdSs1D8eNshA89CWHAH0KVFjxY
T2PCgxBOpTOqS1xoxhZnJIVltD3p/0Sohb4q4bQ3soY9wlOolRDsKlTrIwSj1Ho/
sguio8jTiSQFtF5CwxYbkR2cP/A58mU3ARGOqnWNKyqzBKIxUBvevHUszc5Mdoqd
tV4dLiTyrelq+TkqUdx3rvCX1sInpjEFsvjX54knavgRMX9xLU1eqj2ufY37oULw
opJhVvIUdBDzSQZAU/0Ijry50flsDRq2XQQe/YjFZ9Mw4lGgqBPyxxLgaHGpGIAW
bVzSZ0f+wbacc9c44VTjI0tTbzYTrD1a0rZYlx//KTHJDdETbqAjdg+A64CW6h+H
hBWrhCdrOxJ40elmNF87HuZZWrsh6H+ASCvV1m1+Ale47uqq0X6ikQAzFQwzcFXO
fHgm42/tQ6Dw024amvEovVpNg2V1aF8iAsZSl+CrubKH+H7TE0oSAgK3ghwNlGP6
oT/mw5u1SqaTRcSY77lOddWWLROOVlRty1ksSV2AocbYV34MTw4X7ADI4D6C/IKn
5RRM/roVVXRKvE1btgxSC0aLtunkCpYLJUoaA9zawww0dE9QMDDq3egPV9E4m09v
XGSpHAFy9faAADl+qsJKiIA/BCug3yX5RkTh+xZwDtXO0tTIyJFyc/pYfHd5Lo4R
gk1RbaHMhpHUj958rG9qgeEqqfkPBYVtec0s4rS+snlazLEHsLzAPLmRBp0bF6qb
XKW+L/uDptOJD/CAXKqzEUN7MAJJ7+ULGpk3k4OxcA5aMaLu64qqfg0m0IwVbHhC
iEJju8+yQiiVRsy7yrLd8NYCQfm6gn6+/QHpliisieSucyoielREzT2IcJ+8mQIw
rUYvLgjehyS4MlX5Nreb4326Ulebh26rIxaft1utffIYdLUQVNr8k8zw+gjiTxGg
Ql6hJV1bO//kkZ67q6OPOKsxUmCVWCz9K67jGYlnkvZnPzbRRdVyhjmS1eVWPWKY
74LlXQMb7TAruU4xHTFgw7XuF+rizqdiWXg60rpEg1sz/1+ttU+SUpTOWiWjw/f3
Vrr5wwXr+8LuVji4lJttx1pZ9W4j2YrY9tpabnDwYOYEnDVa0JpfCBUkLT8p8hHQ
aB7GrhJ0GZ+tl7XcPc1eiks8ywiUuhR4ge+82Q4AaHTOpYhBfc4AXdUUfLrEytts
4kez81ePfqLilziXpE+v50wmKzPaG70WROWK2Nf1mxrrDxV20/sieBYX+8klCv/K
kzVqcJknNFQCwU9KKGqjJJ2VRLuRgE8lqjvu7ScpqdUY1IeXUoMZgJFypCv0RXCj
wgjDwa44Mvniq1oaWKIH/WZQXPXxO2Z3lo2ojqFxGgI9JuQcfpKtYuGDQKPLnWbU
ic842oQQtZjSmIKJgNj+EHg2iXHsAVgtSWZT2yXoozCeEyRyTCSaECYaZN2SR/oV
BX5pdrkouZj+E69wqK6/eKQk8cliBD71j8Vy6ThCLHXYN+vqaXaiypDOTK/gDywe
oDuoCS5fhhPeJIPR885kEBEoYSSD2dNTh5Fqa05tDBE3NaZ/SAN3HWsJ6RecOqWh
dupyFEpQ2UrxgISc2ZeqqkPFzBfFfjCtoIYVjNXSgQ0jExj0ZRW7jcloNyGHsjAg
fTiOGlSqz5i1KbygCQ5JwWVgpbJf0niLCP47dcaFdAWCv6RhsGZwUqIBU+g/rmgP
HC9KQH7pL4tHT/L8lenUI/b9cXO/HJ4qiTGrGW96sYFNhAbhqzKymWfCV9EIYIsW
w3LvWzNZF1SVobUDkUef7Viw1ys1+OnGee6iGIp+dh3nCw6v+zDMbBAKUbvSsuyw
You/ofilzUvg13bf+G2nZBpuYefs1ZA5qmBn0RL8U8lBwzXnz6OkdRGzbqGlm7CI
Jww7pnd3LRASrKas5dTrbj8YbbfHE7CA3dG/2YSYD2+EhnIgnP7hILS7D0jZSDF+
dnrix68XLYXYprbIHkUX3xDbdDdl0gLPvEtD+Drrr8V72ZGWTyaIsL1Dfz8G/HZf
Heiz68uZWrjMhwM5Ps6U+siVkkQFW0PN4PH/L1HBFftVRp+rptJNCJ3kM4vuWO5t
BmPwM8vnXHElXxfNW/Nhys+NvglVEfg5k6yY4MkBRCSwYJSqbHpIVHGW52aC1SLa
bbgpVzt03/Jl1Jct7szjlmX6tatAtFDqlNuiGkoTKCHV80DjDwXK4nGDPv6jDWdv
ibHjyytTu5kQ7ZYIpQ9cfXyX7obaWPLI9T8r4wS0NIDHewdbqIKUAalHaqRJ6ne/
nvYYNY1lcbhYTZA+m5F3NqO8FpfgbjqJkg8hf+qXavLI1HGg4YpJM9neZADJgbkv
xiynBrZvv82lkT72KWXQtJR+yhboeZtfEcLy5F+N05uZwniSzRjID/68tuebk1+X
YxUNFKBCRRx7JNnrnAiStl3pNKQbI346loJdcVmfYu09l6oXsnON2bft2halTJVZ
xFd/42Az7h1/qBa5ciSbWLZ9UG9UGfK/A9iqoXWPOvTjxZvGrsSRBUVFR8ga4kbg
8cZzqlyWQKT13pnXDXPT0xKBHzXEAOe4e0zj/uNm2k2YOFRfTcq6UAFeId2FmWyE
MIyGAiP2xMyi3mIh28oPzlrvataTvlvzVGO5jP0Ws5aeUWXpDjIGTrs5FTJGuRTm
DiQouoPiJWI889SZXj/HafQA3URNNksggnym2oXAN0Qq5cgmc+bMIJz2Bq1ueGsn
+Ig3mVU3tmSJYb0MAwijHibHyLd+2626bg8wT7pIMCKGitSw0S+zsuBQxhle36ck
ZuGsuXjrQvyjwFrYTRT70Hr8NPjj1MuLXjbLF7YbZK7yAe13THL60oUSiKVaoQGP
BY1z5qm3jGQCbb9mwY7MRwE/n/qGM+Y+DsbI7pGtrdnuEjVlqpeMigb8TRAyrL0p
4uWH0lA+yj+BqOnbULKDU1tsP0t1Zrgy6YbmhKyZclDOa+AxYXmBRKfCbYn3we6u
IgxlLuLpESfvDO39SzKvNCP6RPGnGgVUh0yupXORbmRrYmGnRLSPauebDdiDU9+o
zHwwtMGBY4oqsJXUGqQC9NaqJbToHGUupAZoK/VDd3liUibjjdBESfxanCoSh08+
Jdmsjoz1dj0G2KQc9d3DGxP7XjULaRRGzrMszcvL1SdQN8PNTswLMiLA1BPd4mHk
jcxFnfpvvMWn+qUALL5Bxg0P2kzLq2tr8nr9YHDfaSt2t/HwtjFQsv/g20nR7K6c
SMdNIbgCeuvGhaKpZsIOrluAChUtlwpH4Ov40IJOXzuUQd5yhmFpcM8ltjy0EqQr
PhhzRafj5tkYyQkS05W3uFvjopj/gKQJKkkZHHAupVCvlamPObE83+htw+KnuxJD
xEV1pdSsvzZtGGUBOrvzHLgOlteetQRseZlDtsDb5ZGpD/nDKKlEw5IUwmaq5b0G
svpdxNgWmeqFG+nzk2Hx637NhNjUjXQvkLVj8b1TsJf5aOc+WuTGVP64qUcUj4EM
IOKNcsvEUmqfMr4B4BowK36i3lHv4/mM7PHaH9pcTCAK8vZ+02Wz4xQIuosUoySB
8Nu/BqLGYHCI8JNgKWMcqtSW0aWHW8qyVJyZpX/K9U69bcF7cG12FlwdRVbAjoRA
YcQ1eu+8cHoym9+3hxXUj+eElTAQK/lahTkcQFbbT/Da43V9spJaMIlOA/2hHLKo
z7sqAN9liS+t31Jji5s2QvEQjgMYUE1S1MJX3F0VczT9AmLGOpHw6M/K9P/4W+lP
V/hpixMUWzUE+FgI33S4I3HFiwouyT++d0qHlP49WIYVq/zP1v1Twp90hDnzDG3H
6AEZE+fcrAYTiklmKSX14GomYSWE4p2OtuNmI1et9LQRlctubYLJ3h94SBMHVt5l
9kWINEEYCGokPUNETWPt9CYXQnGG5ItBe5Pqn8qQUuiTKBdMTYNpUWIqtGoZ7FrP
juDzOSgQIeg755qO1LqSIZZbH/dCGT2U+SCGsOwYpuvSJENXcT/DbNN2c9fGs1jV
YRUSpW4LJisn1w3eSWI/SvnPVnAtT8YSEWkp9ulADiTJELefqnBoMxfVsZxWJouI
xnOjj6N7sfK437wq0Q9ZddAgdW/mSENsvyoISG/eJ4D1Ax1Xfj0gMJn9fdWXLDd3
PXL4iK606JqkRKPqUGTfu59MN/fHrh5pckhW+21WxXcN4cfz0dPfShNGWUMiHu9e
RZGXObzfygcBMqpKbSAkrDqCpa9o/alWsGMhWvj670+AQoZFJ/pb9piUEaSn1+fD
vUp4zkXxji/MuSmPF7GOGXPIDKIUqDAGbP3ucdM7CHBx71tJYRWGyczQNuE9eMry
f/L7uXR7b2hkKnDhWc+SJXovFTBMlm+g/MPpJwV3IhnWknKqAZCqbzsOmAngEhHp
gJNi+/joxq+q8fdx/Ie2jNs+puuy48gJIfyKLWVeYFUJFknvelkPoeEfe9UzejBd
+DxNrMkrd8fNbsZYZ6n55PmZGjG0pUvfZtn25WMhJGZ+2eXHe4QnpkJEJtLBMJKT
1ZA6U15+PfsM9/e17FDzE5ZcHBe7uvJHxjc0U5x7wFdOtzJ/wo2/X4smWIElUq7G
Z0Ofl/841mzL/hohEgrqzCgN8vRg+rBA6GBOltmHTc+ZM2VXzvv/shbeQk+NoAWY
WfYIkeRU+93mO9YUeTpfBNw9jbOjnGSldWcPSELnaapNTeIgWr4Ge8q7LcVtgWxa
6CAy4XwZriwHnEv5G03EMbzF8159yFI5Hw1IeDR7UbFgKrS/39CNduWgHZb4ey1g
UN2/g5MYoHMsa6DQun5fn1rzzGxXA0Q2kDt5kVMBSEos8SNw62a1hsd+dm5sdW/+
s4uFbSiKW5uD6K5aTKKU9Blx1tafMdfpDrgV1/+QwhxurEqPMr2BtQ3kXul/62+m
SVU+2WX9W/VPMUU4jYIFtinS/A5KP7Zk4SF50+tlSqZIZ6EAaEPE0tL/+ufojqgR
Gso5BL42Up89Y3daBpGgcRa/kXsCpMpVjJmOn+ziydiYpOw/t33fdJHPbfr2lzck
X8TOz4leJc3Br+AHrqdav1G+I2X76ql9LTFXjbNNvJmKQutZ2QaBZhrRy4+t3rhz
3R/Sb3HdYPg8XoNQ9yXdn1zy4dGSAjN9RfqEJ5BBYXA+HwN39TId+drwed+Zsuf3
8kLB6uhkKbrhqYZh2cbDW+Ggb03/KoBKzC7sgI4KvKUiEhbSG8N5sGTa4HzGL75U
9+ODJEyzMVgj2ckt7/NVlWuL0uWu2A56G+DLmMfwxN8l3LODT0Ai5WKT1C1/FXKK
EEkEuGP12itehYM/o35GtUnAiLJCOZ56aXPCTJkVqKtrRIzHDAaI8HrmDwNF4Sla
c+iSjwWvLIb5xnjMZ3ixNzf1iqgt0u5S41Prq1qyz/iBFofgYqM5l+42jOfy7Mid
mAPViuYeAQQ/pOF52UTjTJMAWr1s9SDhWwlSZJwK1wh73gVHfte1ephm40IcXzWH
VR3kWB+9iDaeuUvIzzhxupBVm11pDgF7f4W1GnfSVJmdycVZbTHhhdC0g8JA16Cv
Yx2ZwEhXynFllk/yAwWIJUVQAzpiNkH0tH7HDou6IWV3EC/f0Mmtl4WMXujWfv8n
aAr8jPKyb1FHeroHKUgvve2COGwHbALDbFJlBjNASL7ijoG9VWRWfqvWgSdKXLUz
S3Ra/oTqrqu0a4X5+Ovcsx3Y8g3ZS8s4/ZukMFwlIkCz34ySzVpb7U8BcDZxYz2h
/0N0wNsDIuDHnPujstrkTTUQ2VnmBopwMBkSabKkELtLEWqVtNXFCNlvDTsUDj6A
6duA4puyGSPqwvpvItWxOLSr6SZp3YYDJq4D2cu4+NGA4xcI2W2+xzFnkAUMtXFK
zZqr0fBkUtUcjxRNdhE2oBEr9SVH7NV5MnlAbcR5KkhD0YAif5ILRIHpCJlUX82F
XB/F7vBsfXEdqDUiJDCsKsftgdwZ5EK48j980g/4KCw9cQnoWCAF+r1tZVkwxKOJ
gosiWd3GqU9jQpkfhLitHddaDS4O7QO+ryLj9yGTSobXvj8vD4UuFNgVTZjIEOwd
aXVs8f858o2udocsD2De1pyLtFAn46stQTpA59wjsDXuWTQcWngaRx5RyYdppSlF
5Ek8uEvFZEByZUWalF4A8A9FTyI2STMca4S0AgE5GMK4eNnGUlac4yO0bVAdUJRi
sfI8GQ01skL0M9PXGFbZhKhsQrEnQGELLNJeo8i5UYi69+vndz0MFwwfngVMT2zD
nlO87xWkH8443VIXjJDktUnnaygRVdUKnUHzpY0S54aQJnPnUbeouPc4Muguv+Mm
7Yh9wskoNTvnl2Or5aqYiTBbWGlO6GS5Y2S5uxMy6W/5bp3i266PtdY1JdHMiZoX
/WOY/sGJM8K/vrJalMvt9lZHLOFQXxvoGIA/j0D3IoE+86WByfVXlwJV7ueT430Y
4Qwos90b0ww3lWNCVM6xaH++6oxgys48sAsi6t7IMYwXinaWPrH9yBoBdeyB1rY3
ARnpL4zSJLhBwrdydbAMq4vqiYoXEJQ/SqNn4jzfnMOZbAwf8Hfhc3VVWkn4VamX
WsR2SivlUs/+RbNN8RBiQruOaOnB8TzNEgEVgorCDtORK0TbrnCmhK8kjvbIXVGx
EHVVW8DTaSpLMT18Wc1NWigsJs8AGSrQtExLRmjN/gh+k+Who6Sz/8+7/8/GJm8o
p+FovevRN+OM5+Nbmlk/SeLXjpo8ZTtBlMUOR/Q9HVNQan6V4yDV2n6OLhNmxuPY
fUFJgPeN2sHOxtcJwI/uRObhqOlnk/ODXGVT/23mUvZRYD57OIfL2nFRqdGg/NI2
FqQs/LwrhKsR2k+m7x3A9PkV00eh8bm1hQewAtKDp6mnA8UnH2prO8p4QxHVIbfh
3CreVBJVnXUxlL+54365AQ3fPTyTVW4bjgLCYU2ZmlpmEsvqjQCmwtCakqDQ6Qwf
azfUKst/QluJjmvFnT+h7NWjitCZeTiNdry0MDbLjzB7V9cdapzBRZFuf/0LTpF+
m8Q/2+HwxbRlHJDlmZMGJBVSNznZrG0n5mT9/j9ZQ2y2suuGqh67zqJT63ls2JdN
XSm+8YB9QtABWHo/3ZoEK6L01/thydTN5lKDGYOzB5QUOsOMrcf23+as1pKCiikN
qB+Cm4KzGMil8abBEBAkBYINmj6zwVsTJSYgIDxf7ODfUXBea+4/ZXhnzm7VP6/f
C2HXwu2nhP2Jkh7LXjumQ1v/ziCGrWstdKjn6IyNrMGqbmns4gjQbftZQxqcJRzy
yngGUjzJnqzNlSmG2eOHJw4hJ3zVep9RabCjGSiAl+XOuId9jCWgmmG04qk5lYer
h0YQ+MY1UxA+PWSHQTItn4NXn0Dg05WBlPNPhOf6EqF2szTz5Z0UGaHnwu7FbZPc
oyVJCeIwoK9yNF9zQsH5zcNBsNmoC5EJ+fJzWj/rCPwU5SGqiQKrZzr8KlidhpXy
Mn9TcxtbDzxe9YEoEQ++D6MGBhPbmrnAXtHcb+60ghwTy808olw5LtmW6zbhuFI7
1UjQ1zp9wy5p2tTI/+gtrkvIlrF0pNRdHF7H5CqIdSB8sZyoo0lUvWkYkKYC1CiG
pdgycdA4BptenBJVhQ1vCQJoGF8aW5ShDzr05nx8UxRVSfQBooJ5t/LTC6ltcGkJ
g1R69Ej1F/P1OEZ0UtnvFiWN7Ai1J9R1iLoiMUcqAhUOlblbOFvszCFJrpRU/dXp
OC0bJd1ceHlAiVmIlABBLWIaM4RoBCIXY9+isenW+ghYi3z7NjYj37YKpFibe/Rx
ThjkbgUUbFcBhl0AymceKQKsopHV2SCGVH4yt8WK5kNsxsyFicnaKONYQU9MAY5B
1CvCxGFHlEUPALVQG4fzVFf44ZMVpPMwk1XpoH0N1VDXJa68FVsJ7Uy3nIP120iB
3iZE/Kx0nJZAXYhBVevR+NKnw5zRXwJrVqBUUB3iTQ2moUJv5huBovKc+EyxFC6x
ginN9aKNFpILAJAwRvE1XJEAELcXrh8LDmdwrh3k2O9RW89k8+zxmbFPiCngSFnx
NEJX4FB0n4vB7C9VUX6B7UdbNg/CzfkbOBFfCyX9YKExkfSP52oaiN34jgI49TO5
4Xt3vCCUwSl4tvIw5SUFOnDwgyE1vud3Ger0uesRg+1pGHo6Srm7AzxCGJvz1szU
yTCEDG+HBMYjugVvH5wRuyE1F+rgEac6snZ7G6r4QVV5cH3Wp8neCkfZ8YaMivDF
6Et/6imUWSYxqKijTQdzCIFb6ySqKh+zvE/ktFaKcQgc0maW8t5UOn9n6z8glHO9
oLIVDPSVhTDBKNK69RButpODQZG2P1nRu8bTnp0b+uME7h+bwB4uOm7oiyv4rzF7
WcvizD8HjzU5C2h9Ef8ivX/4bN5ZUa7Yd3Gfpf/caIGso1QSdy8hyidagAXkbPoG
yaSDyW9CkWgq+6Hdb7FmhcbO/9Pb20bnklBiWjDfyorC8eXnMaD1O9CYaIJ/8stP
AOgkshEkPVKSN3oQBdMb3t+GllRC1vdAgEglanVnUcoPrDvR3dJuowPc75S1girU
IKTJMGnnu7QW0Iro737OtoGe/jFd76k6kvxt3FxKw1anckJjOPc5IHz3Ub935iAY
3w7LeH82NpiYM7nuRywtn3kL5Z2OgvEI+u5eUpNbK7eze2Ov+kjk7ejyOSFQJ5mR
3wD9ITUKKGLvELQkQGcemU0HJJvb/riSjSFoJutrwGAhNFBdqmUkymHM7rei0b2i
ywfaaPBPMQ1NkjOg3ZfjzpBMovk2NROXBUBfUqCim6sksbgHta8iZ3ZgLJtBSDo1
cEJ/RKP4I9TIfAcY6uSTHGRw+7hsDPJLi1IAG/LdCm+wUSasL16Pbf2QhWZpxOtO
tMVK3QoGEsK4+jJLWsIs62IZIlR68j09hDLpifisl8gT3Nf8LGZwCLAgDfmGq+I8
FtysAwpRC1bvP1VuIFzaNML0ERl9qJjini/VAwF6B4sPFMDaY3v8YaYKa1eREFgk
HKh0sosv6nd975wDq9z8SGpbs6gpj20KXNlIg6rSgU10eqTL7IjqNcVZdSKxAIXZ
5ctKAbgqakbwXqPrjKoFeUfzDaJWDHTteALYZ1OD+HtYFtOcxNI3sYMfi1Q5rvdN
pE0EDrDfzzV9NuljPw/0odcUlxHzFppxR+X67N9Xs+YfeKPTEf1mdTmDaj/C8JN2
Cm0uF6a5R3ub4tO5VCUqeqTXLSzPKQZPKe3eH2R4wajrIQldPcbCuljAy6VhkxaK
SXKpxxvvj/HIsXJeXSgRHNdbf7TB1PmUgTnTK63SSfZuN2q6nupvi2xP13RLpl2Q
Xm/mmhQ/Q1e27lw7SIr5/AmCkG8uw3i4tKWvb60LgbZCgTAfT+ox6Zl+pgshaaRK
z/vtU/YTrua0RSQirGIn3VDVIYVFkW64aCplpxuCCTGk8S15oVxRLqXkA1nzDN13
XzTbqq0lQxc7tJalmdAkYK+MxDM2UkleifU2N6WsGH+lEEJnuvn4x2kg//SEeFGn
b2KB1NFZnFG6I2yj1LCnAAADUN38gY4FjQGr9lutQdyJUcv4FncsDFNj/vQx47q6
B88th9xC7htT4co1Qk6XBEmSO0Zi090BmmmY380N8SlHEC23NQ+R3nKgsyZIYhXQ
D/1/czHzt7830h0dLapNcdHSJapzFo5RHMQMwPxyaXWE2bWL20DRfcT6m1lKtzks
i/zEJOHL9LBBdeITKk0N3mwlIxXJpUk/da3Y8cFHyiv4g2+d4t/wq2Me3rHMsQvq
BWrewyMG8J1m0BGKd7ciT2w8LRNrsTPC6hLdhyE76CkSWEd3yBF6/SJ55pfpzhYH
6QuMpTm2uMxudBNCpH8oKAsouPI+5NB/dmXcqfUcJyYi/QuciP2GYkGiugrt4099
JXkM17WDcCncO3SiZ/G0ryE1ydHPZsNLKP2icScBanv+6itpZuR8o8HEjPz1/09a
CetMXmyAK/la2aHMuEgkcW8vqO+xo4HlolECSvLy9MG0ODO6D/YXxrGwwe/NXvKm
t/3nl5u5De83+B/hHAAtFxEOFC4/snmquN3SzToCtExS7lTTG/2IpWFNyQVwGnZk
d4UNF1c2mG7xN6KMnXMrMR3GYFq+oxGXfwew3MqSyo91836QRoj308nYVUsKH8UK
MgRFupl4kMqzN18UDBKod0QjwqgG/Y8KC3B2wYMpdQI4YEsAbFvDQGzfXYaKBv7y
tCIv5/tWbLXgGOrsIJR4ieTn99SzatfpZOerOM57aEJu0686edjE25peZHwOLatj
dLYVoyWjAh2S67pcv4iKLbxHitGe2tIZlSv47Fs670Il9nMxCPDnIRLU4XmGeEC9
8nB5URnoYqXD+tNVvtAHUUdrtxdic0VvVAdGAzvI/vPd2Z+tjRF0sKANebaYb0tO
H8Noepu+e6p8cV+gzzIHy+T5LwZTyh41qG3Ex5tzhYElZZLQUOX4YOTIo4389F3o
KkONEkCE0mUUU9JyF1q42i3QDzDnYAcLC4fgpNnioQ1A0fJrGBhrhE/ON8v6I6MT
0l4i11Gxs/c591lmCniZc3fOyipCS/0fTUKywOG3LfxznwH6y1k0U4b4f7rzwP1p
qb/8JCShX0CXKQv9xkbLEMD8doRo370vlcNsf/FKn3e0yvckGWKJyPipZIFdEF0o
povKMgV6P8nZBqoZ8JVFKeGCbzkwMMfu2BPZ7c6tBZPWAFQsRY9zdIh7T1ZOEZ49
7dfgjS1FnmiNuj3GNRu6KBsSnhT+rVmX2gdv7w9gFLwvJgegTvdZfMvc4Tc3guC1
W6WTCvNhCfCx71KcTuRICdxDY47HV3Q1vaPWbKlJ/w+V2zArnpb8iLLLVGVir+B8
5Lq8fj4TcQoHffFX+Js/OsaO/z5qda89SZoJiFxb3CBKBTxYr9KarbDsq4aYQB7/
iczDfxfNKLtezgg00jgbgCYSIFnQk7y4eysl34XIK3hiuLHyo1mSRMtroQQhAPUr
ppLKrv9YSTtwCSIXS6b5AGaSnUTmE/r+/1Yemp9hokVXEKq5FkXt5EOv3xv/SJf/
/BsjWHPGPe9WIqBlGtXrmMvBfTeYzikkLCJkqCm/Yf+JkeoEOEqewI7ASkfxSxxa
jrg/YAzPI4IuCiMS8oyRgGr0eBjfGrUcyBRudhKOcxRiNuN0cT8fkCzF1i4/RCqz
pBnO5arRMa9bny1G9qXHe3GD1qgel4K7/ack/Mj1l3ICJGfApo266azMycTf/dix
Xw71wcbfd2hoJqUWF2ukqCse8xoPrpsA7+pFEHE65YEUygYQD9w0ZGnQzrKMcOkt
ZS9lPwJzQEfmkMeDeaaaSOqVhV3qrolaxDDVi8bY5Xtt24CPDjapjfPebjuAAcWM
HAIRR73U2dOnvAMqkZ4CRP5LCfRi5fqkBUFeCq9DZFallipdco0eo4F5e2OwaZ4l
CtW0oqdclwtoDqS3WbOZqQdWvjWN5ngYMO5nSo2m+y7Lha8Nqyix6+PF+pw6Mlpv
dlLCadyE8g6EWnGXb4y4ShZSu04V8UZ5FsXhetaTHu7HK5uGSp0RqrA6linn5kDN
jBlGeGoJOZ3m3iRUrOz/cBcbZFU2v4+H67HcF7I9pJ+6T/0Fgzr37F0VHSCbgxR9
mIp3v5e950Syr2FgQdzLG5Knl1/VcBOlhXez9laRcxNRIQLB3oqOsolsSM5E8LrX
vVfOtgCqYHzP78zp9OmSGcfdu4L3t3a/WU99jkfKc8lC/qTgXizrbXkrdtT/LntZ
KKtlDTtrDfUkRfcVYG1nOuWLbx45Tj3ksc+wPWwHevZQ9ZMx4oyjIiUJKgnTt5kU
gEAJZOGhjCZLGgoA+QdOmaao8IML+s3rTf6F/Z0ORzRa+EBhHlO+f6kLF9fH8tRZ
rwrdStnTFiWrMYIL1SLV+O3C+BtVQtXC/MkBh46igbieYxfbbzXmLXGlR1/w1zQB
n4CW6xb7iyZeavjVa1M5Mon+csUdqttVPu2CXkx/Gu7EuCI8LWIWyJ4bVkoKqsNV
IOHmWK+875J6vYy5MO69vbrd0w+7jydPqsZiTCzlH/BV1WzteL0ZxK03HuCKQEBG
kpFyvhlj4CuakR1NlT1XnTGbfQVj331bPJ6HfSm3Tua1UkKrSbSjQmwCqcthrmsm
CTIy+L2JlTH5FXeKH4p9wMppNLKdYQlUYehmgsZy4gS9ojA/KeQJyLBx/XAg8DLw
GwUndien9KE2g6b9vnoktqpyctFZjylw90bfOIsSCJ3gLJzZ2+smfFUcpmiSn3ep
D07bORFZWzIuGtHMysjd+MITpkey0cDFGAwDI8AfVGriAAnebZXJY1kupbErlTjm
0sTsk/GUUiYqZ45co6p/eeUTu7IK7EGI7cx/pu0+RFJTpdkceE17pkqyK1wtmHZK
Xg3TTwznnrwgqKY1skpBwMaJ1YThJDrcX3mGLej0VaAqUyk9G+4j6iUZiZ4DslZp
EWry4DMW/7HOrFBBgLIo2WOdVO2CuLkDmpGdAVUDosY1GRnBtjI4gxTIDji48w1n
dwddLuMO9Vy8wfPLKMWOa3+4+1gipL4V1QVBfjjikRdk8TYCu27lBKSv9UxJBk+4
Wdzj3tCITLLA3R6e3mig5Zmo5ypeDYNpI4JlDnAj3pAXBjJLSL4vx5qRHmj5Mlmj
mafTRhrwxXgqHfjV9PICw7qHqLeAk8dOkhPXprcy2Tk25ZfBerIVtPC5ktFr8oFG
ijAcjdZJ/VnSjSFF806D8efAqzjUN6JK6pQe2szXWE71qrfkOic2QZDQ7aMhBGH0
2CV7ob4NVjiR8itICclLLIWtYmy6l8Ow/kLIliMBmbiP/sznQwKrhzsIk05rAM7o
FRkHkjUcLqPfVfwSGe69BzoFr2BGo+0gyQuiGfuaDxC+721X7Ji+ETi5HhP+R7CM
OJXkUZdyvEedAycXfTMjDpCL1jDN3qdz0+frlSZEIz+DBBFBMPlaqfp/weSqoU2d
upjBkJA0LrMnQ9FV5kY1zZ/fLnH6ld97dHcySYShqXBr+JhOgZakp2ppPXMdkcqB
MCc+GaZrmriA+d0UHz/fQWf+W17g3kpYI1EqNaDQBw5yHjzmEzIcc03bgIFYAjjA
/jXenSbVpxEt8Q3x8SL4+5MAfy1Ih+b9OV32XpNSPlR5NrP0DfHQTQgT3G7zfD9J
BmC5TSJAxR9OqLeH9jpHC5bSP7P1cIM1ZSX4ij84o2aVDX0sq0oh1Fxf7MVbpfX8
CEwcXV7XxFBB26Ct84U9U+9yU8b3x5GMfXLRltk+3vtmZk1HZopn+W6fxc74JMpj
utlHVpI+oF3dKXhhpYwhqo1xPi8Q3YhEhKiDl9Xx8cHXMixmSoHwFRxDvOaxshcT
d23GQxid6279ZxSnXP63seWuiIvfqXh/eQbXE7VJJA9oUlpzFRwlgXSZaGhmunOL
HPf7iIYRh4WOK1eg4iB3AG9KtgD8FdrPvTZpN/XsLqSMLhhie6pEPvzmDJfCEvxV
HtqEyoIuVFjvknugJs8KlqzhUS2Qzw3qGmFKvTaLWNgbfkPgfB11FVsJusYYk5mC
23CLlqPQb5QW2he4E5dzG92gFr3ar9vSICyUijIX5yA0XMK116acRPHBkCuRpqQP
4ZoJPNB4PUaEYgYZeAv51zjfGuUasJIOdD/97KcqmnAb6nceVOxUSyJlCOcae2rV
+OxWF4C3p287P6ztFfyBOpKKJzG3rteiWsNO5NObg4lvU35C51Cn5jvr4rPZje0T
Q7mddPvJNBJVSpQOhZ1JxUYnN4dVtEG8By50b4l56MB7X0nanoA6YAGlmz/VQKk8
TXrO0Xaz//IvuCAu0k8Vvgc25hamHIO9/HUKjP2yH9Xpjo2TmbuzXFv4gl+7hNh4
2EMQRleEsuQzOCTxD9f8yeZHs7ymgm/q84hVwkNzPi0baQ2uU+Pe+m425GGduYSd
sbbf67WvXvKFCndDee2nSgualxSW86YCuWUFBwBhxrv4CW4tVLYbYZidd23ammS/
XGoVZ+6W9Kiv0t/CRlkauv4Vedgbh0Se7gJ8+FLC2SxtEKdZcxeYYEP4DG4p/19n
GYDzxOX6r+Fbh946mNFH1VvMuIFdxwghCzrSDjtni+UoIZ2Fi67Lgz+/JGgeh9i5
JWnS6T7k8vkOAFkxCr2QPETZ2B6wSnXvux18nM22ykMnq2jBzEe4FXYH+e71QUic
qdXkyuVz0LBpAEzLx2DEztS6j0bBRScyWrI+HvhSMtyq1VjQIx1yQmuais0q9CJS
GgefFsv6eWCrrIBHjX8JibwshTz6pdZlzTimkkwEHCLY0/i0r4NZ5H3OQk7xHhKP
bha6kqXsWXb+X3XLefoS09r8s4dPacGahbgjqcep7YWqgetTpvKLEaykjTxQJRYJ
+TE/xd9zItoXvHWvpdxUxc+n8AXZ9NKAbmsx1ixXihPrFD+KRO5s5madHeoNgTUy
KZR4Bchq3rb4V+Lcr10ay+z2bTUX5+YFtYt2fFKjY/kP9WdKbGiLW8kf7gf/tQ1z
tCjlDE2o7luzfwW0eji/iU2a+4BmfXarmmP/+Nu/MLZ/qqRWk6egMLk+ge5RydVv
jvHXe2yzsTg/a+dNIeWt419ee3DV0yN7JPZwGtioJIvgb/NYaPcRPPvznxYXmp/m
QxNb7AM5U/uwoL+EvLUuWI/10SACqOFooFTT+yf8D4BuFOYrahUfa7cjLB6ndeE6
RF7jSuRfSRp1e2aGHF5+NPe7s6R2U7C1VZ1e3bTY0Ufh0zEyZn2X4UUGmfAL4k+h
KSKt6SkYTgL2Q2QOjTUE2BhGCVR9u0DRE0FXwDgj58V6AfiPwI/B4Ixl+3r59TQb
Y03EpNsZyfSwLH4ySu627cGfLQgNdRqf8Ib3gktUvNIsPWYqCtwmRulLMRHNUYNR
8Cv5rQjkwfg+5dp/ARd6W2gPw/1Z7SnDxIquwyRuxVuCE5WYa9VxuJwu7l5EdCX5
Vq0OXZ+oeAz19dHzTZLl6xYNN+IQfS8j99sKch0s4byEE0QNlTpdXAxibBKou0ZC
nMs0v90R5ZbxsXX12MYdh422ZGSPKhvq0ap1IMsfmDqGF3q46TpDT/joxEiRRs6p
F6/1LuNwld5r7FlCtoAgCMsawgawoDaaCHx13mVLOvwjp3PtZ/Ml/5IddlpimEqF
0TfLU4WMU2WlF/zFViDURFLEVXgBWwdfMawCFQ0EbU80Fl5zypENN1u5I6Scj6qV
9jaSyXjQmoq2nmMR+5tDyXSXKjgqpSz4NHSwUZUh8FJuKEpNejcACvcvhGj9Ugj+
6HIzL6siYusda7c3FLjxvS9UvYKaX3hi2hvk1fSn5m95PDjQY/CCLo8km9qmR8Q8
ntKMiHYa9kxbLZPjHu8EtqbtZdFdaWBQniJ6S1s0Fi809rzqZ9L+G4DMDqobnz4C
tNryYBUQ3+bCK0PqRzgY/RauSRLkKQWDL7Fte8IY0qCUnvZCA1YE4kSMnnLXmHN4
oahIWlHgtkY6M69TxvwdnF2kB5h+G0eRLLSWASyHbGDDTprLxzBdGXTb/vSysgS8
NewZ6s3vaPMsALcgRr2G4o9f2pMJZKD5LyAQIdEPxpmYOj885aZHQ1789f+wqaOC
2uYP/rsLuB9eGZQX+i2np+NVoHwq4FQ/acRb02xI76d04Fc+kAXGw5xua9sTM9D/
7ltJ5+42R7yDDpiJ9YtseoXSYbeJpHaTUapf2/w8SYKllm5iIl8Oyv0eDsWHUd/6
jG50tH2KOofl/9KsyxtVRLVxSMaJcjbYqdxOBX6Q3z/57QdbmsG30fv321D2/lQQ
9V3gkJahhkSGcZFGPtGd/snhHWQLKkFnE/5BOSiEg3Tgm83LpFHjMOcZ+DRTt+uj
XFraWrk7Eol+CmowXTva9cQPtw/qBBFXTGfAm2cOGkJa8u3w7rEbeajdX/o2nUIG
IshXV0Dl3dCdBdxgV1Q5h9wyS9/i7CfmxgrxijOsboJX69jHU6w+gIJfWZsbpAuO
YBjNVWamC1aaaCjKfPeybpBrOcv9mjLWP5Cag3dS3rLA9WSvZ1eApJI9Acuckl30
nD7lMTbU2STAbr/WbA3s7/moPCdo9ti7ajWx4T/M1C5lDHdtQq93dVvtS6J0W2uR
IUHB9OAgILcc/GmBj0f/t5MWl3FxgsgVwdryTlSs+Ft6thzE+AGR0jDo3i0Xz1Ym
fn6k3eLSi2/huLU+SRIgsohd7XTU7v8OY9G71MqIborN1qjLbGLSkDRtVS5soqgr
K4cWKScJWLOcLlRvuqwRb+47rTpEWXnfbilTuxZ0X9XR7xe46mjlhOncCkD6NS+E
YH134cpdvnanhRqvI6R2ThAim3NXsxPyNO/P9ov5+iFXlSGoya8TtlwDAHiG+jG0
3hQyMTm8Q02hkLpVXwG6khr3pAsY+PbVQpHOZrhWFlPMReh1jsq4Dc568R3ev7Mn
3fpfzZmEZKq+jxWrCypsTZTxc4vWeEiGnjrn1ymCy6i0iJP0PWY+ROHLZ5DnLd66
D0bj+qbpG/MM9TT/41SEfau0R8dIQIlY73NNNwNHyxqCRHCHyb2uK5wd4TWw4AmB
UrSnJPvnI93pJEhM3lI//RbOHKaB/LmHVXaykt8h7iTOACf91LBJNfD3h+7oj0va
1cItixqJxRU2jMrgGO8a0vnA4ua0ImDdEsOfHCS3oR5fvtgOIzRiR+3bpVm8eXEN
YvOXzfJV798/DJgPqqdhx+46G/D/2KXYyOoj0xANmV9G2MophifthqwrCy1GHboh
NsnKvuFfyx/KgBs2cIs3Ls7QzfA+51fEB0rc7gw9T/CDjucgOYgK8A/5ebcja6zi
R8p2F2Z2Hp5XGYxRtlUV+NQsFZOm2L77vAdNrWDDHEaBCOC2wmU7JhwITVU9hzrd
zV9AbZECu2SzTiF60k8jggKKd5mEqYm0fMXZJBEqOPONW2KGVLsMuUkIjwVRB83V
kaMpMz9AxhKlLbeb1awE9+vDDWHVAklGXFoOJOF+VjomRlq2b7SKcYoRzB5J6DI9
TKMOcnf89x9Cl29cMkzjmAJSvpBshAPHhh2uqwVAHBLlBlpsAVlh3G4k+HBbglUn
FQGPSPqoHNWjpoxB2K3Vd3aaltknMi8NO8Cmp+CGvYNOgWqRDbVmLU3faWNHajFZ
DHzeqpb6r7Y3KYoH9rwQtLAhOsr8zq8VruDFeuC8ABBu8sbGspdXsZPK2rO+nu5R
Wdex+dlnTe6WlKMS4dfhF1nbwK1FZtGVtxjvoO8bfoYbrAsGwW2R5TU0qo7GkU5e
tdYPk1gMirtzzseJsS34E53RpJM62CRAdEpXlBnPPmdrfosKqMQyU0ch2atBP63v
us7Q6AVDDlXCIhR9qA8GIR9hKX+RkcPtfeVzjRiVXDySB/lIuWJS52eahEESiaS7
3JGhaFHlEznCIFrpT8nZ0+I7WZb24O4UTUhF6W5BUUHTkWevRPtBtzSvW6/aAI6Z
9EI+8SzUqo/2svQvT5VJ69LPBCr7x0RhmI7/3KhSyXAa4OkhVYOglzArVxQd+Ah7
V4c2sH34IVu5WVyRjxvwbsCLs8y8ig1TAvM9GBwvM71QvVD+saLP7tsDvyFwHGwq
kbs10rYh8QVgLjNH32XIw9N2fQ1fWPMD4Tfn3jQ0Emn779+4sRTEo+LfULfI2Y8D
IBtf4jGMEHGKpoOsWLaqG5BBcZ1ixXoFlzmHQzebAT3RRZ/LVTYLiC0RJSfLyZmx
rZOb0jxjnvGcMOMCYY3m3jq6r7mAcOBMSJU5VviupMtHw0yOjjXkcVTkyr78VUcT
OOXIodoiQF3wUvKVoJnzsguWyYNheRcpdVLO4naETojz0ZyJg3xy0VPBV3U01VCN
pAvJpP8xOhDKB++wfgMkeQ6eZ68/HQX7rWck98dY/C0ScZLc7+h7KUKd9FwYlCho
shuFlyMnHsODkVgK1eVUwpojLFjNoi1g5GrikC8otp4JaEyAxaHSBs/7MN8RopZH
4z/p1acwm4xRyqidv9hZ6jnd3xmOAXdXsajphv9xngEGiX8DpHLebmvaQqqGU5MC
bH2/zEFuUtOP0Efl5Nw8cX/wVqy/i8hfPsGIPkbnHmnMvnqSHtr23wHbfEnU9qIg
FjtkhA1zZbSEooOhc3X9vlBCCfXBr6P6Za1T+cXRn0ZW9ApKiGOR3sCT87LjydZD
AwBYo0oQcmNWt9zUOrXn/ss6eHnVQWjH2tfDBoU9JSO12+K0hZ1C5mLqpkVJW6o0
jhn4RZpbKEWTWtE+gMzyAmC8Zo71aX/O9DNwX8XNqQ/B5WPzk+r89TwNB6cNIu0s
CNgZELcUU6NkaXBAP4Ekei3jeCvUqTN7tfc0aTsSd9ImC0Ywc2zv9xFN1tl0C33L
7RgYZ1p3fUQDaTMZkwwI3lrX2b8hys5iQc0rgvQwcDl4BtxbmWxikpN6eZ7zfbhJ
+bGU9x1F7M6q4+2jYEqJhdttWLqiA52knJ26AQArxKXdxPXrYX1ayfChNQtXBoqy
dsd9iI7fY2DYrdf7DJWQTBW2Y5zPYiFWZaKo69fhKtykyEQhOAxYEHzzqNMiNSX3
AfezK6blzuNE7xPUPfuY2L497uw+o1Y8unRmVcNM5pf9e3IQoeRPIJiYQDZtxbMu
07lmxivXfAvCIZYa6rg/Rn/o4AKZoIkJR0pV6OpSBq2yw+a20aZdowIyRAYZCXqV
SMrkUBdDYhtpjOhaRiwX8KeMjja60AMdcOoFGfbZoXbv8d+KHAXafwaBZ15i40vu
2vPpfNCRef4RlnFL8KfIrUOreKf/vC+Np6davzJrXznTy0F4OIkTGS2tyBZaXS2U
DrPcd0kBIM8MkjSOBewS+AnMC0q57HbIsdYKG3Q5ih/ryWticRA79uC+CnC488xa
SgpjVgCmOCyB/IyoZA9xQ3YICz8Tc2FRbWZUYkIJQCXP6bENrd0cyJ0O/IRwim4d
q16u2hFwODbvaIu9bHNo1bTPjEyQo7OWwmD5Z4s/bdWASW/U/WOeIX0UElUCAKFE
jF1aPox+VRNimIafCgUdRemSlhrWJUeJLYsKWrKW2X7xd4wg51D1jFCKQH+sw1b9
u+sSMjR5OXoCoIJbtW9OF/3c6JUd5nFlgTHfQh7m6qM33awNffCDRD2VSUFkbWfD
KMIcur1Gs13bU5J61gFF4iAVuh43mrU4M7R3JpfK3zVKqmDM/8LpGBi1SPG/oMFW
hcYGD3lHUoRsAd/Pof4bXoxjmQarVpg1yXZr1+8OqSAlXvdoGwW3lPqVgcTvzE58
kXODmjnp+loFhCVglyA8dJvCpFVY+lD5PH1AQwrIDnPuANhe6E/R8shdjiRJPo8H
NoQGbw90GInyyEhJ0clvnkyVYt5IGrJjOsLPy0oEjo7jOXk2rGLsDy+zSBWTHAGo
Ijktx3zbNgI0/B83MP1Oz62KjMdbckRVnYQaH2Y8dYYQsTkhzb32mlAFTQFlHRoc
nyh6QpmyqdrpQgCWsSkqtMrBxiJ8n/Xr1KtqxFo/ilQmgKqR43dA/0VODPnEs0yu
y4Rr4ylji6vZAo4VNMM6SQUWvzbEVAigrqxGpvFD40kd6aE1P4t9k6vDYS/Mi5A2
A8k+AsTt4l3HZr4jeW3NV7G82CEAcJ1LyoJ+fOMFHHRPiKBoiauwfKXXS0kP24bY
e0izkYi73krQidoggozvNpdvd9/JshpozRa8M9iV90jxQ73MUZcqq3pcfx7Lk9qk
AE6dlPVWLz1jIbgMotnq7cCzkZF7lsQrCZKg6Gxus4ctk0zmRVZvH07EZ7phTCsj
mXJp4eMBx03gAeH1gA+up4oH+2bc7nBDgj4PBXmp0Nks1R4uhqbtyyOGOt+Th3yq
6FYR3O0vZYRuqXpaiZPINZju4tsXnmYOOKF2TWilFGudKgMBKHPRUxNwCGklSHiz
Ehm8S8cB5Tfo/2LoMc7Z9UfXGvyxlidqN/zHPj+z2FXoWzj5y+qoHZN9pHb/jk5H
OQZaP7IuHrWZ03WqS+rSPrmKjHZovunF+gkQKX1SRnbGrTgaw1pMf+dYT7Ngq4DY
sdPjIgTBk4boZw8tZuKW+XW+vUVkcqlN1nj7t0phih1BAghn5zIVMQiLX26Mf5TN
eDzbnjxrCHKgPrrKWJjlKzWFQ3nndVKTi/Ednga/8yGfhyklNnC7BEGoPlBPQ/ao
2PicniIAbiCS4YAcDp+nNWiyS6MjMeR1ZiycEdlBXqpXfZDCIUkOsbM+l36MOZjs
SfO3yK7pbeQOhAstfSaZ0RUM3K3z6gCND5ROiyVkAtb4dWafra2DCK4/jo3eK+u8
O2JL+qdd0UW8yvB7bsSe4ikxZvS8GjrzVoIQgjwvYs8hjsR7knKY6XB8CNEgZlg2
VoRbveXfnDZLcL39pmmCDk+cpvIKytPRS50IRk68A0nPYy3k4/flKrSoEQGeXBBa
W0dcrHEiZIh06sbZ/VH8ZGdDzTwc5bGtdGxy4LjCm9x7Fubw7rQ0Rw+736GrwF3j
r8/gYtatDVHgxcln1M+wetIfcYEaPFVxToTXIKGpSpOVEd5uoxerzOIdbt7LqkVZ
XGXKmDwXru0FKGrWRnynzOoPwSsd31w3p5eXzZiRZTUj/GTyOUu/GfTwDg3rf/Re
HlJvVYX+g9GlRlJ5GV8te4vXYhu9AXfAxZWvZkZOd+OIgCva7Oqf/DfvZIDmXaOX
jNpgNx7bkBcgGtGuuIWg8DVblzQ+n4G5BeG3Q4NotVGWBias6K/sTRHVqG+Nj8Qc
PTDyQ7O1OguZx5plN5WCPCqttZZJ4A5Tz3f/B2K8tHE6YDmHdI7Zez5NvZWbpCE6
rdh2C6fJMYEcGvVuMDosjECr1/eowZXlWJmbrRLvASwZkwUEuip5BqoRE9N3nQz4
BkaGyfBOrn/8AX1VhYGAToABIawolCEuCs5oX53QewnHBCymsfHDO5THNg1FrOBX
wxkLrsrQk9ACBhA4GiNX6zv+2H6oeIlULrWcF6bFDUkBEFUads2fVDf0L11139xD
PuJCfl2wZsDG+sO34n/sKzCaQ34zkWe1mvtyYrssCCmVAgeWfogAYYWJUQZG6gfw
BbRRTUZCufoCqv0g3SndD0Ykg69BHBDlUwHW1JBrL+/ZROTA3vdillQDBSsF14N2
kTm5CgsaGjiBrjVzrOVDhBdgv264c2Ena694kTdeeWk7fL1aJ/4QZO5Mc62nKhRM
3vHyM1MMcINDTsHD5Bx7008BStKL9Z+i6sBxl64mzH0aE12oxVFtDufILaT7Pr6G
QrrKzm/BY2uAqeMZXyZ7WHb80dyBtjeZtbQbbYnKaX9URRP4ONKGVfdvbxVptsOv
EZdLmHyKxmCIDplfKE1pzJ/wV3lBoRTCIbXULH3pGKgsFlcAS/Z/tbhjvq+ZmDlY
S2iK/bzI+PYp9ugPAS0vNgo96KNrVvlDVtJobpbvU7//eL3aXJsBGnFkwMpPZgep
nL38MY93jvXyLHbzy5eH/LkCoD2U7Z/SCivnCuEeoI82HzqVdFE4oPwdZNxUu71e
880NEDBswAo5P8UFrb4Pqc6y0d9RjTVNblR6vewgpXW5TEXFLMthYAQG9aKgwIWF
OdqocNAZ9WZ6kgyPe8fVu1bVL+QYW6SOK6Rmdaqovg8F+v9+Y5dgnvXZt5EHqhmt
gXjLn/WD6nHujZxsMJFbcuJ07RPA/xaOVjx4LI79CutsxL0KsKEpwJBJyrQtp1W0
+XPpCjVrSvvXCiGUf/j3tp9+SIBb01WXN3LTnUfc6d253P+r7LDw+mmqJtxORi40
xtxnjsWgKwMd1wi7kK3bIlgwwh9P2luLrTHhjZ1MzvphD/07XjLWorZ/KP3OGIUk
eZRbgSyORiOsuUvBbW8l70anYj50sWTVNQU3CysQOFsQWcp0r1ddvRGUvQsP0cql
Bs9Nkwg1Ei3FPftS1muQ8v3Pt/l3pNYLYmb2Ft9pGsO9NR0qlcxa5UFQU2kJqx46
VNMS3Je2FuhrxSPLZZg8EebDaLouo+lfll7KjdM979RMgTIGsugTqo9s4qz/k/gT
PyeXQotqTqvHZ/4b4a1l1/QryrNlv4Lp4f8DWyRua/7XwzZtpXhCC+bJLDitiOa1
loGd8YQRIzl/ucDZLgPIbQQJN4E9AgWS90mBTcivtD4O654yGdYvd1zCcUv4ZBUb
VjhHQUeoynYyFy/swbODj/aqm166ohUTTpeRfUHax4LmPniCT0Rrv+aBe4J0bh4Y
I7coBfNJdRSMmaFBKMuRn6hrrIO4tfHEGqF6AWvE0xGI3Hs5qTAxZibou0Gzq+ge
cWOKUiMIwWH30Vuag9xYCJeXk7sk6XfhMI2xo0DVSCw9m9lIpB0n/5VK/pgO9dKG
1rq6m5w0d7wYPjTYMYEsHtRW4ggnORpPOxWFLez0rtp2AOt1vBQsombiv3ZmEvHi
m+meYcBDsHOV2FxjhKBbG+iQwNWSrDt/U8LBAlqfupbmt+ib/ccEau3dFBkn+Vks
kEq9io5JlM/DmVxLGe6Qxhj2wu+XkZNAIG1b+seQ8uI0sG6WyzkrsTatCJrITsQV
Udlts/MLtIICVlCBCbyu3QvkA2ZBOScZwsgReiy8KzakWApKpI/aAONjyI3sbwVL
T2RSHmnqW+zcWt5Kx3T5GfRHasZVANdEyDUEj0v3gZrmvJXBmTds51xeYBb9GYpF
0AIiGTGWZDdeMAh3l0Qtqrz1SAvlEmRJGOgglRWF37LAD3rND6ScCZt3H0HodC2L
S2MV7mdKEIdb+0NFoOtme/JgrbevAMbHG5vXK0CsacPdQJRmHzujIJGo9Ze2WHvt
fOBBzqbMWa1bCA1IVh13FyEI9/3gG/xAzJ8O3V9FUNKI6WRSr+GCUhBCWvqtC6S7
lxQ6WAOnzrPemRJ+nOjXWBr/dIe4QqKKzGhw4HhJ8XPJpmIChJ0tlXVelOMBq9sT
mYESjtvGfX8MPpTt8H9tJUlcxc4hS22JQEKYmOSQ+QKed9AMNChvGpZtwoCF60ie
rHWp78xAVh9b5ArI3l1psZ4tz4usX0+0nzTJb+I6VN8QrDAIMMZrjxFMuf+cMoz5
2ABsaYJ85gh0ss2wTYDYPWTwAqUukWbnkDzUHqnk5ZGG+INMo5ntSpc79Ti0Xxo1
SMmmOWm+zfc7Cq742oO5hHTPGdzDHFl+5YlJHnMYqynnlGgFryegk/N0q0Yp+vA0
SW4BocKBrY6iRdU4FoQGZtXDhPy6ylBznOOnA4ytwLXMccUORo96S3DunijjJyTG
rQhuMy0xF6AnvIuQLqRXweOtzW1fqfXQfExm1KhT6jgMHJ3Zgo6W/5tLwY36VEOb
MKWDUzIpTgDAUz5Z5xcYv8NE7HLUMB6BhTJ64uJbGRfmHuQNYYTc848eGIsqN5jC
9Dk/5rDP6Zc2d9kdKZajLatKIdXCSTCkyvK8TNRlrA328hVk/nzBGptI6wXmuqN5
7bM2N5+DxLiF0PO73Yks/kt9MNFTzVFxZ8V21SwBQijqKZbX/3fwFxPE84zojtRO
p16MZuR+40//O1T3PkrVsILFo6xEpIxixPJ10ayJ0jXqbLDkP/pjbaun4EUMGGec
Vc/S3th3bmhqfnlpmvxoArDH4L/F35hSd4tQDV8boV1oU/DZnKorjnOUvjHXa1dR
zeIcXPARCxIkZDl6sC3ZVTHq4q2OYH0QIaqL5oVS5EVGZywIz9asRthNfQxKVmSR
7DOjjRmdZVLGaS0wEfICIrf6Zm1HQm2AiUT8pxTaigPDSct01CRksemiyjy0LplD
zsy0BYsjsAKLJHb3h3rMwe3/K5CsQRupJ8oB3ItSA/cLIdR8nsFIFSduhKnT4xhu
AORxn5TMhoMg4ENw5BpFuUPLgPbpFyOTfw4Wymv8pnb4uAE8ZU6AS696UJ8KJaZk
qqJ8nasJERY3XsVBt6lDkYBqNtJiR7megcUfMxEoBCTScjRkcW/QWUfOeN55Atrr
63wyXfCSjqhwtXKQ14ZGSmpMafvMgjQD0I7Psa3uOaNC74v/gvyzRdO9TZCnsw3i
02KJ2hJjmydCmkFGm8JHMOI8BOgOKR/AH7AdX44npW/C47TjAXc7Oz/Xb5TirLzp
e+C0iAAuWcjSl8VLVBs0RdfxdCb/v0Ak9hyjNxHFupeH61iDdXyUXW2PB7TmCnlp
oG9LHGvrH8FGjdSNJybASa3hRxE41ZoK1UCtWyPgO2Y6563HLRMIbtbKENqAwrc6
qrZNkBkqALgu/FaZUs9VIYny9p7jB3Oeh1Yp54pYFXwFcMlpcNT3X5wD3jDtgorg
wrlvKZlPfp15jbvUWtnonlCzcmc3RMFR38frI7X3lMeatlW/TXqchQBxvGf4bLZI
oyRzredHV0vmS6CF9xWmo7iFCUtfAF4estg6QLDktyjXF4a7N0pDbWvfNk8l2RXa
yIQhbOmybhIabd3uq+CJuMuuLtsCNT/TQECiZmnumg5WiAaWRK1CC+/9YyF7EHbq
F0POfa5DVaiYGRTSUa7B+AlopDw9oaHW9jNrPLOLGlENpnk4yI/eZQdZMAmOeQdF
sEQfcv0xqj9IGMGnxqPudLP+xu0EylBANf+uIZHbS0OzudJW7ifQf79ZsWSc8S+F
EalMOdy3DLp1tT+yuntzP7AVYOtrCKgdt9usVsM2+lW3JatgMz5jTsU6dHf+yFd2
V8/bR+D2vWol/+uOTS3pGXCPZJj4n13xeUMYLMlWZiQzYt/ttZWdIaZ05vCf/0uC
jftOqo+IqZILStWju/Le7wy7k9Xn8bC1aa1YGrlXCh2O8ALGdjvj5lVYQx2+k/+6
jTSWBUdEWcOxVL2ql6rqMy0cfLQ0VoHU3FCZ01e6Orl6QQ1oDxtQrrJ+O5mFB+IW
pjCpaCgIAxILa6J1xb7OV1M7NAdZFvQk0EvdTPCk6C5qy/h0bbnbScUDJ8mNKpV1
TuhkcJ8P05KymEPhkg/rFqAqWdrkrRWDd5m3rQiVyiOWcwyDDXIZ77DxSPcFW9TL
CWFW3gZRG1i3kIh7NVERPGgM8hGMqbCj+aYXlDUF/KB0PRWr8Mm9G38pExrdCJot
MZzcRBCQbo9nSDuZRGZ8PdZ94oxwIn6vAtImCuApbwcraK5+5trwjvOeTAZsWKGu
bgymEhLDVZ/nvuLcNH8TrGvc6SpqJJxsnq37uP/EN/rFDK98I4CTbMMlAQQG+E4I
BsT66LXOKMi22+zLkOf34WYBHvZdVufr7yOj0YwIU0PG4l06WNxVqxMvJLJ4VjgY
pjxwrC4ulpkBnqh/wsGdu4PiWXs1p/qONNhDyZRr+fMpfIKWvhqa6+UhYUfSu19L
VkbBCgKD9mcwo4BquvKl6TW+xjJhgal4is5QWfpkKx8JLjs1cvhIP9js4C0XlkHS
gs0T5O106nFcMgdGlOVrO5dJaFPHdaQuUwmIhMi68sPqyRsOdmfAH64hYZyyUMuI
G/UXemjn9qjV070Tj2yurnHz2JvOC8CTmGCQlyljgXjCPzZmtK5j3Nh32CuIJggO
ZImT/zyWUAd+70HscS1v1rJd4A2cCqD2BgBglwGRdxQiuWqlmTCZZcLcoL6BdvT5
ywow3+tZ50bRIBBrBnbPySR7MXx+F1VwsrCo/8rvTK54fj+1W6IWxeI7dNpsrisG
CbH4rq0e8rgT4wIj0eMt9dba0UVm13K97FpQpbxMOb/0U8rEXZiGWfJN+6oAv99g
zJ3DsL4d9o4LfjFL16Kren6uRNDhWd2r+AyPf36VoDDC2Nqom2Omhw9qz9kCJOnX
PZ8+OGtpSKL7RjAvYW8LftkM0i1LoZgevdNSLmfDP9sXxfum5zKR530gqSYQxYdL
o3MsHTo/aZBhxQxZjoG81gVIxnvmNbW7OH5naxxkK2dmNjZjAtkYS63kGZswUIz8
sDe9mqEloDiDGganQU7ikNg/NNQotYYirgpJRo83DjxAhIOhFtVWZ7kiNyhtPlOg
IXSowboWOlYSCib3VgKEbGONPGfx2L1YBB65+cAPIE1UtPOvOzZPi/zhadNLrUuk
wOIhN3mY2E1fpA5m2Zd3ly0DhNlgw9BxhBeDYNWrWhlvFoCiEebtaUicw4JLR965
Der+Sj4r9g10P3fh2H0CrS6tuN3eOeUrJcjRRbN046nr7g4S4EjBNLU/jA0NBw3x
i97HjGhoRA6/Lw032ofrCfEWy7fgSD60PwdWtdIh3w1hvRSpGk9Ue78xM4q026YI
noGDIdFbsHT45XwXvOngrVMRNfAjKf/Ghi458XyzLadSLMAjM0MnuS8oxHYVwQC6
WA0eRSbi8e801UQvF8XYfOdNIgafpLwA0MfZD7cuVAoM8Gwv/hqvbT1IcdfUXtse
BbV8NQWZuSmFOvyDYD3dzZ9WXq6h5fRM3wYrzqEemTzFnCEE+GtLjC7YUn18KBM6
PTrs1oIBX4OKeP5N8oxu9KhZ8mtZXh9xCbDM92/8gmzJoLaeNH7RZobeMFZX53A8
x9k7A27zW7yq4s+I3b9AcSlzZmjOMP4BuzZQi4o8rSIMCkfiXsFXmY+aJFw4b3F4
ZLJDyPlOERdhB3l5ZGw2OKJnjC9vVjBf+jeXTrDhNn7YG0W6erkwCjJtap3Q2a24
hdm22PwX/8Kih3/O+ajPrYbdwpaEmHNqTGQVVzRcxL4kmGaQpTAaMVkrNMpdyLhP
i3BfCoj2UrY7dNpZJfd0Vjq3d8o+J+5GrQbKn8+xvblCV4CH1tlD/4JxUnBNiWhR
XFBt7AwCqFy8uXANs+MCDPN+60fBd+/07NFerhGutyEW0nIa12SW/MK8MM5WMe8d
1LU1QVa1WCetrRS0a7i9J9RV0RnKRHytZwcIKMd726QGnPC2ys0jgYNe6lfMqizQ
s/bSHt8+V/E5iwzoC3vtdVG5feA8BmNtRDVkPbzPmN+5f53LmfA0ocYAsus/0DaX
NiZLxgwsahkm7V4nJHlKNIo2tyZQnjIVOO0dVJDusucx+VjUKwVaggXYIAzT6WaE
4+z6A1PDKMlIPQ3cxtRUa6A5h/fqdiwBDmFRQhaUIw0okZOCBjfU8yyuvWcz99Qg
fniNpOMIP5LFzziDsLbxA0rT+bzOiLW82sX5ec6ANpdpVrTrVUGDs/vA5yYzuGfA
R/ai/lEowdvUooZFE5YuigWjn0eWYiwLINghQ3OW6KLsTo8rOIFkVVY05BKXN+l3
v9zh79Bq2JgPqzTWM2bTB3K7elwQuJa7+/H/G/jSrg6NV9hAY0dqFBTp7MLKl7ej
uEJ5agW99vEgkkVlZVNDBOMDw+PUyNeqb9y9Q+anapMJol+7us0OaKgfNhZvpvUI
QDrrcOahMqD7ihQH4Hrv0R2AlRkdjEjRDH0eio6eD7UdHbwVIeNuGUNM8j76FYTX
E2uan1hQrKWZiN49e/dF7G/J8UP0sQHpswHd7z84VBipWmFZEEiKOBTiP92PGTuB
Tag9aGeHDMJR4stl9iGhZGdZVyltWDoOnZE8Qv2HWiXu3CiPp1FF0KlLmKATaj+5
qr8cLjlzFyCJZwKvNMraOI0MHhSCHie5OjBARZAnIf+eT8DsyN7jIy4aj9j1c82z
/YzTqEzmTnaK9Htw+5JqKAfLM2u8dsm3Nc+sb9K4jLs8T5J23JSiPsAAvIidmGlN
QeYNhl9Pm0RVDFrqD2HF27/wmgDF1cnVpkYP4eIIATl6NHOHaqyq2sXzLnLnvzO3
x6BBglu43ZS2x0daojqDVxGk/i3Q0nCqs6c31e5jUdvXiRk0sa8z/qMZuMiODSqH
hExsL3Nxuo4uXZAGDDyb5+Y9G2lEOLuK8w0sW6uCe5t8N8+v8S/TpEtauSlzaBb3
di0eQ0+dgyVDkiv4nxaMZyXfBzfeaphNi6h75DEgXRJnYg+Qv6xOALmMtkNZxe3+
vRzOD1PhWwjDC2bAGUvgJI5VoLKwiZdQKPrH3TFVXj77u1yvrasrY7EQyT04C3uV
EyVJmF8r1+kXWK29XUPCfiVMVR6B7G0Fhv81t7sWV2kAxyrwbbR/0hgzFWwgG9BW
ESN3MtXQ+F2d9PRco0mPQ2jHKGNs1QUQSllDi3oowf1MMNBFy/SSyi9sBX9ZFWJX
dsbT+hREfXQOJ0yWnpvwNMN7dsyrE992ZxFYdY7GrnIm8+vZLXFujDBD4XZTtw7P
//tSY2RRIG0yRlngrFE94h+Xs+yhloYJ9HAQpBJjw7MGEJNoIBwCF5dq/hkidiGb
7I0IO+4GgWuR0UvNQaL32JXS8b8T+xkZ26mg0eR6c4V5PBvZRMbLB5tC8SRK4ITh
kkAPMBOOGlISQC5qPzyj5vl6suCBWzJPNJTXGJd9vX1u+CGWVk24FR0COMqDLCfd
XRC5Hi6+C87wLRJ/kCWOWBeN61xBsBwE6xgf2G1XUh590i6qukdr/Hf+V8GgdLLu
VzUplf4Q9PyvMHlyT8dvJHwD+iQNIfz/or9FG4pYVEXwg5P81RLzV6m5dJ6iISHX
AvAicQ0IqZmcHRKo8PD0eDIb3gDi1CFDViBrxRIXYU1udeQGoQ01L4izj1OgdtqQ
6KIOJyoI18pgrNGWcmMW70dJTbTdQvKAEV3UGiDhOAKKtxE54k0N5Xz5dn8RAn0a
eEwLVSxinoKUvBHP1U44DjNSJxih0ZhwEhPBnNt/Zqtmf96xzRFH5SmQre0GYgO8
U9ohnLf7tnOCkK2SQEMUo3xO9gFOAN0HjelaQEzItng6U4vpU5mT41hbt3FbrcBA
nGmKmLvh2iDAV2nGVSze2UVU2XPuhHuyuv3lyNaiNIYcDaxHc96Ts8Wy3zlW3Sr+
s9rpabftUG3g0dQN4c3vkEX+RzvAR2Lzi5BeTK3imzYMbodjLBZuyXMfpc1+J5Y/
ovItbUt2F/p+lJXpSMJcryPGx/nhcxMX0nsIv0OGF+SmNOOJfbSF8kSCtPk3rJiR
7W/ynDfoSvz0K/4eMjPJyHj1yJbubSq0tNxI6jjhEpTZjJZodZMr8BKUxg+VdjhT
I2qCEd5MWil84/eB0stTpCxNYiNouvk23rgSNwFU2PkFgR6uyHpt9Qm3rq4tEKlr
5YYjjet+17E3/mvM6f8/8UHZjKUBnWmVnLylieCikzjbFzcK3Vg89ZCKz1akZ2NX
eFrJnrWKPOXIbtOl5m5cxKzwhE87607MU2BhCYthK1dQ420lQ28b1yMq3+xsKa8x
nvOMCfTWQ0gvIZPD5tDex0baXtfCK3LsjDterLBjAw2fzSmMMTVrVvS8Mjrpr4xT
sP7CZyYrqL7RUEwgAi32rvlCqrlM/PYNhTIhe+ZP/mpAiiH1EFqdgxA7veu4pMY8
iru19nqXYuOXbE9fndOX4rYnxYrgVdEKlZWgdesuc2I6L+lwonz8pfY/xyV2M5MI
uK67PAjR4gKJHZZ6Gi4i/uOrV9nMrJojTYFH19RiIQuJmlYcHQ2J9iW5NUm/hReo
BLbz696O4Q8NTF3OkRpZCOIWaYMes9Pa+o2/b6It9buyg02csjND+o1sHfcnML7L
3rpu5TTKD6WqbgrgYxdGLHqUVA3UjpgRTLf5/2J+EgVfhQ+ZXkzP2XJAQWoSlad9
AaAeEFJkLzd+Zbfq4j8lOcxAhMVgSHZ4BWqEDfmQ88jURL1c/pbKAViBfr0AFn3Z
OcfOYLW0CZ91PVOT8+K+V4VoFIb+K3TetS1sQ1rOUXEYlCTE0U3KHWeZi/ZsBo4e
X3RiS9R+WjKKon5dlybFED/MZyuL4gOHIl5ccVzy5+0mpax2VUiCjF0Vm1ok63jF
MqgWAHPXNHzxA5hDRzzm1oFtzlLckUcQf/ckAHXChUdjCeKfFVltUW6ZYQCF9RA6
43wb3KtdfQoFqZYnOotVPOP10VoWSqJU1zNJJXgyuyQcso1627A04DD6WSJyntwA
hnGfuPZQCPP7RinlT8mgqNL1gSw+LyKJLPUFfkQYx7Tolyp5xkuwAumNdgJAhcwz
ZvKa/Cpx+wSKT5Jn0mcujuwK/d2vG15McQL8g+L+vgYmFWiJMJhsHClWhPoOrgfL
AWwVaEy1dNsg2qiWnmOw8n/sZxIa2AtVa7eac56Sy75BU6BGSL5YK9QPWObt6l9p
fw0WL7oEItVxikHSIVjU/u/3ti6qUZn5IdK0gBmp9bunGGM2F5dC2zJWcz67Yud3
R/cZwFfr90yikOf+9ZPqhWWGfUc7uifliZdLNLwCe5FAFH5UlvU28Pd8sZMl1fUG
gpw0MOCu3cC/+4R5W6WFKZ+JqKVvxjCYQsMG8kUlBpoh/huUKOAkj2LcSPCrHZY9
k7tXXoHftrQ/TIuhHb3D0dTjvi2rVdWjwkAOzHZVj3D+sbk2/naSkM9v1sP2zXzC
J/Pdb9dZ0H1HeswxByC1j/qv0u5cheNslOYJ6Ch4XaH/DkHJVBYw+QF+mJiCAGwx
zmuAc+mgsCKR5SB9zj4GUNbGN8ZDnXOLN4G8aSb+1Ij7xiSossC5nzSN4u/5VhPt
QHUqw2W4LvZCiD46j9ji4BPSQTa5AqF0b7vVtPDbF/nMV+bcvYmPhHKJG2pVMmA2
wz6uGDy/+c3JxOwpQwF3jOpmU7Vfc6ag8hd2aR8eRl259uaESwIVeaOou0XFK4AA
d3Am+2CYDMGP2B65ZStDoF4F8xiK2PQaQHX8WntVFcQ75QAKyg6MR1nzyvUTdbKK
MarQshINgY3cBfEnUdGzCT2mYy8gjCe4R1bypE4W12zz4rVqZzrrtvWfetKHl+WT
10pbGbtQ0Aeidb8qPpuqDfEakUKg/DE1xj4XDLBVMg0dXHN9MFVh1YA7h6qKErlK
8TY9WsvswUryxRTm45cBz9FHT3RH1IoHGxAu7YBuhd2W65HZo4IWNH4qOKagZ+VR
+1wpoKgupy6SGfCcwTtJ0/la1WINVnMYJb1ILoeLr5foqubONbNkESmkAXc/646+
IAmznrS7T/VGVo1cJpGdPIawc1MzUQRXiNQBmsbJocX/1RqQCfXd9pAEfigU+ZiK
eT1uP8XsaXkjwQSrLmezoMO30qyYXKN4gvpdfD3groAZvj+ohtWQWn8Jt8zljzwo
p2kjLtbBE17IkqEbuwI47+weoBCOk25HWzfrx2lNJITLDk4K1X3Qh/zVvmDBV2Lq
2HAWB4c43LMq4wK9bczXOjah60D8z17u30eOdlYiwEMkahyaA3gAfqwFMMFrsmCw
32OqPBe4Ju6AsEzT6pBP0NWcUlmgTQzxyFI1yjce6i6penXfQxEUCqC8XpgIiBlG
q7mxteAlA85kSBerJUep7MSJzikmC50tDji9hklpD2GKtRWaHUDe2Hf3vp5RtvbG
jWmiolU+MSjBDXOfzheOwYHTfwyKqh0emK9k5N5LeQ0+bE0o9cG29owbM6z/N29o
6Bfe8LEoSRLLgIfdv2keeMTixh525tIp1tOSsEERqjXb6wSYfdD/Xh6zOYv4H8/r
4MAGo0cJz6EAP+GhlNt5yfWPUpp9jABISnQiohljAgPl3gOpsUNCNT7RkVALCuND
VXKqiAVeDB8wgKteto0UoNAE1BXbQdWyuza2Lctf1oAHmYJodPeDdX5wpR4xwV+W
zUZ68782im0e5QOSFMBhj7sgAU/af5nlzn8orFakfgThPWHMDtheK6MTegT1KqoR
ZpMdNAWhWj9FVBhqB+QO9BcfoOko2gqF4VLfOgruzbkXuJB9UbE66Ryi3APMO/RO
yXsTnGVK/+0t5XXreBY9XQiC4ToxCkesxlvuwWX6ZwwIP5HoQ7TNKWvx3Q9NDPDL
7p+fNAggtT/cVHevAc6PPliluhFqr0qNLjCjEas0sZJhPYu4tH98O5acxhTqqG9z
eJbcUtbU/6AfDY5AXYCdt1pjX3G+f1d9LEuZHnK/BGp8g5xkjuf+U7Z+PKAAKvjS
fB6NQAyB8jzE2G+A8VLaCcPpj3vpKOgzNZeRnrNExVraDZ/a0dl1ASZCcjPXXPZH
dzkMMqwmuyIUdBsthEeSvOb3aiAwCnkrgkLgBW+GLuRsqvIqNDaFnApyB4mQEBcb
jm0rA+P5dN1wfF7GEMJZriQqn5lIVF1fE45Ab9BPhGBUjf0W+En/hjGp6VGY4XSD
w0GuW8l1y4ElEwXp0VF46yeEirypvhZwTNsQHF1cDjHksVqxphleLc/9Pa9CaG4Z
r9FN6Fv+q/Q/m2byi6o29NAPbq7aAtaZbh5XKcRd9p5AbeboGyq5V76OgnT3y+BK
90jhvlES+mYNsV4ztwI6s78GTUB73ai5Vi8h9n2vrOJAIGDGLwwTzC7DdKmZAFpi
vitncODY5vkLExoeSqaz6qMHoNjzNPe9eYJm+q+E/38jEuWIox/2hMDaYuVY6z5/
o7AuIsb+v0gx92TIFlJTlfCdVtk35Ba+8Z2auMXYzEjm6KrOcxhtGP8rCipN1JfR
ZiCQ7n8XQfPWVjdlf83u1+PKsGdi57ut/RAbg6zaqCmPqOxVs6o9Du6aJcHk67eD
TaCsAs2ps4RbxqnemjqH9IEj4y9Zej8I+R2ardhkEuMjIK4JDTIBjVn0IKbLFrIV
NqsnL6DgzvDj6qrJFff4+/7roh53/QgP2ClvuS9Ty5HV54O5pkIqYUon2vhVYYav
kCtvB0kB42Uj4Q6ycbDcn31xgvO58trPlC9Rd3ein/1Uo6RjbGxxC6vKmqoR3FIF
10NP7mWGiHf++YAJJiXeixY/CEfQ/q0JmD+ob1Vk1GWTBE5LVYJ3aK9Nnf3c9JzO
xwl4RsfMlx+veGgwHYwuufDkFh3fgLDEU7IyEQ3taqgOh0K5dSuQKynbbhHgu61T
zntyclkKg97jlwMDzf8eZx6ZPxCu2oxqoonGiOMM/dIaWzD4jMsWWhIbLnFftfkg
AE/mO2rKSJ/OLtWAz08l24UAC/mIayv1LDx3FKmsbSlVS+LMGDHh4xiWTcT/hTJu
1JUYVtV7zEbGE2FSMbBIne3CI3AZFMWjIVgrcFw5AupyQZ6rDTQf9YPaRMkdcseB
4i4q1TZAxpgWZc/EhmpvG5bnhb2PEIc5J2E3xgOTHESgObL6ETX17usacOFH1FCH
bdzX/9TuAMgek6MuSrEMdbywbdDkiEgXNuNwB2g2GIO51I2n4BQ62tKbGzNljbJS
fZQVf7w+tlQeaaMTxDxjKH/I1c4CU4JF/crBILFduy6es4YRVdVMNoN1KtyrITYk
ksj1abd1r0XIU538/171WYYQR9wt/7JMMmK569sICY7EieXbF+zXcu2iCARshM6L
CB9V2AO/nE8sgmKqnU1RsXUJ9JzLSvEEnWMFrVFV8g+cDPjBz7tmrElRo6s0phiB
CkYZl4njxkianDnIN29e0WcrEjR3Ck3uoBaPO31GIU+Qj4dqTE3AYNh8qIehuxqX
y3avkyVarIECTQ9WMtkHriuwB6gzNSg9FLM9O5kOuTC4gWWDgm7t73GT50hPwa6F
9zMdAr+4tZ4Id/cuzClOpwedwGDQcZYfwtDZN20b4w1WxxKDNQcSgY3HmIGaGcmT
qWJdHeRXte6lI9nu/F7clFYMvzjsf2R/v6Eid4zziHSGo4XF/twkSevex/vkgszf
tJhwpoc6mk3plFmgrEVzKAfvQsly84iRBtA3OkENsOcVx7I+JUm6UJ+T2y2Zozzd
ok3B9fP281ubgmDGeq1dOMCRFhQwRf2A/b2cGFJ7QGhFOJE1Jq5hL4cwTfMije4H
q7ivw2R0gHDY1LF37IYx47c0uR1axq2WuoqFigge8gghpqeHJZtWshEUVAeFhyjG
ubl0hbrAzwZlGsuvKpqUhE78FDz0VjJ0sSweFGUBdfTlR+NbbJxZO5HYix45FZGh
PxrMdDX4PVfAeoxrhT/R4LEFVQjnyt2MJDwCSf/cjAZLrlTJJAMbiDMlmJVC20t6
HDt6+F9ZhlcQqWLw/EFoF9yDy4E/CopP4uxSTH350aAem89sWMTa/Yfb3IonBqOe
icv7VOUn4gs6ghUT5ZUn0d/L9BxUCeKj6uMOU0z6J3WmKrnDa8u+FtlF7aFSN9W1
pSJLE3ycNdAk1mUmI9ane/uILPO9LrcYVmjgC7Q6wzJV5DMjflljosAjmAkQVa33
q1wnePeV9AdDvH2Ng4lmyJ3vEFqKup82LgfkdN6zq5XB1O6vuWRBJNyl/LKhVaEu
em/oFfJCLMaW74oY2u4ffcEqw6hp5sik4B3lhbUZviqk096KX14IkPDXSKjuEsNZ
EsuyFLivn0qiEt3fmS6Xi/5u4iLkMXEvQY7ZSO64NK37OeVCUBadF49JM+bwGMtO
/qGBb9UROznrs/KZKu69gzT4jjklK3qaEu2mhoKz3NtJoO6IjVFf2DFxyhGrWchN
hQEnmgAO62QbLAYbeah+h/OcLhBumhciyoaQPOAUMLhhgRR2Mx0zERzmTW4bqump
OMnzzBxnTpu4xdcQwxMHeajJ8+etknb+GWqr9hqHvVPKLhajMc7L832CpjAXUV5n
ZWaX66KSyydG5N+Hhn/A+MIvbPWMwedAty/3GoAlqlTiGn1idaROEiadl0RQsj8p
CZOeaLHSNaUs0l55NhutatyvfzRi0rYP4qOOQzirEWKPrOpoon8632XFRQn1vxb0
H2OWNI4fO3iBWqNtTW2BwX3JKlPN2SWOlebuTiqRW8zyTWonstQZ6WIWJtMmx1vM
U/tWE7BhHOGUvS3f0ADEXLFTmDdDAk0NVTVprQH2W5VRkQJ1QSfc85dpd1eefB9n
1zGXtmpK255oQrAAgUkUJYRC9juYf2PedUvxseyFN7X556kRdLDWL4jkZc3aQLgE
Jd0eIvmK0MPVHpZmAvrV29m0V//H3Ow4D6KdBYOihYrnANzhaL4pLUM35y04X0jV
FcGORFUlaEIWUAxiLCZkEWjvLEv4XQkK2WHMSBxVPtezSO7G0sP4ICogiE2USMXI
TD441gprFEGRTia+kBYigeekGdbNvZgTLhqB0MFBXxjZEPmwbHmSgfPfDuXGN5S4
XOb+gvDMHUtvaKbWbsc5trK8sL7vcWYxBPKN5xHu8gXct0FZnewAGjIMUW9K+vYX
4Og30upLQOJ/KTA9JTJMt2W4qVu9+VRAfQVmlRK5qrIcfALAlXk+F2KdTa387IGh
2slkXxpcTL1c7IL4RRXYrLAFQ+r6dsAc1lC4N7srk8QIClgGvdhCC9W86AghT2Eo
vDRuVGLm7vn7S5LmAzmYjltgKR06y4UX+vTmRTaEbr3LiLeB8MzTDvkHFVvPW4hb
4lE6oIx4OS8Y+TERQIFTxyQS/1npFGcAU/SGs2OxYrbPR4GSz59I6dqixDaZYkN0
YyhQY+EJ32tDW10zvILb5swO+xxF8AvDXAcuoZk6IURmrfZx/EYp8wZ3bANamcDP
33HnvxKyqUhOgJymlTzj+p4e+LWQ/7BaPFso0P1JVvEZzwPqFqiRKmSoj4mln72Z
++wzy9KXIK5L5jIexTbjL2qJ9luLVapwaq2r+EYshbMzuFOgIklat3TUnbf4J0/9
R2wZe04//E+6vuTtjZXag/E7vB0Jo0w2sOklx5txP3fAd18nFZP0zeeGTN7xlWg8
1rWT6lWAYb2/esUmGNg6cD6zHGUwvfwMsRZk1TzwcO84Gs/yyKLlojDx7k7fWtFk
7ARgyGoFmuvGoBrWzBXKsQ5Uc6m+ia1BCSjHkGVTXAEYe7OqnrTU35mHyEb0Gng6
dlg4VXQhuzI/XaIRy4DIW6lBGilrvqxVTgbSQaRb9jCwiP0+eRaS+p8vWVgZ9wgb
9lcAwgrRIv60YKknepLDZ5PIWLv5qOR7RpwAwuBbxPi3LRbbq8YJZzN7DO86XnH9
bWlpvqppUG2vzX/oWyUAu/UFa6/dbjFlh4vC0WCLjWF8SdHZpnEKctaW0PuLnS2G
vuxlMaoholg3aqwAaG0sC7piAbB51oylv7VehhL1+GIgT4jJ0xW0FVoO6SGocAfP
pBJKDYJX+DWXFG+3UFk+fNKPhDOutSm3zwJl8FeVxwDx7Zf/igndK3wL/zMIwUpd
ZDPQLjP3IOIhxyrpmeyRqy2zXm0lk8zjissJC2uvlHWMTtuYLMk/Y6v2JupsshsP
SurLWQz/yUK17hvdroL+1XgfP2za8JMKbJFk9faSu1OxgB1fVXFu/Q+JOj2kkmBS
XbjVhy8GyG82JPq2r5QLso4jss0BDz29mDEK/XUEWvqTZIvJgZiQP/Zi4+0EmQYn
5A2Eoov0ym72D/aR8/UGzTDj5UuwKmqGqRm9SMdzWqFbNcsaoTR575pQQl6x+BbW
nBBSPsu0SBdEs03PENH9+qWREIMmGFtUsi5Eba1mSrDaVFQaBv1omZSR6k5ShkHn
+k2RtL+GFIK5DOV/wIcCPucbK1qM5yqqdU0Kgv5oOtiNpqqRvrS75mZglekXvXZ6
fcZ0Y9QTQCGVzYfTaP3cc6MqkwG/hq/8U1ucKuDJYq4Ec01amF+r13xMAno3TZ+d
yG0cUs3GwQGlUioVOw7EV0RWdG8ruRsa/8jsrSNVZEp1qhVDTjfL1O4q8JUJEkNa
9qIfGuDO2luCc8oubV6Lsxjy8W/Zm7upHX9BlzOa/hp2iHSAknMRix3FypSPnYsv
6jtSwC4MS6mdlm3dUL3ktVpxWoXu6XtSFwAz6U5rhQGVa9DSoPr8J/MNd0PqSmCi
uM0NGsou1LmfuX0pSgLE1eMl1noobM2vzu3MxaQCNkhLFsodS4hb7TW1nzd6pPAZ
fQKNkliyUhedeq8gI2YDmSIhBeWo3NFoeShfJcDfKIzzDDWkMDfuAPL8Gfheg3S1
fe58Vq7mupvx7i8M2+dqBBaPDrKZsf7uZPszqfNRj8PZwyMpAFgyiqSD9WvNPVg5
Rt1+7zOijfwrG7LWpg4zi9sTtuxkqtV5o2/brzak+7bZ/GD+0GHbuA4M+EgyGiDY
gAtD/wMxaauA+HBkF4Jn3bM9JIxWQkks3KCvvZ2E+q88Stih+S4+02nLwkfjK5u+
unftllHgqftMDIPPB0IcFYT3emR8prlkcsP8yks8QYZNZjj7z27Oj/yiUWLHfGcm
a0c/QvPZukXlcQghqZcAYFxzgZ7nCwwRtselIAiZQMDUPJl4z9C6zpykRLAAi9m+
TsKSy3ftjOun6ytRUamR5Jyg0a6htSqZ51UEhu0DOakJkMRK2JisL39xdd0+z6CL
tEi4ct0VIoJaFN/CZr/55F+uRaY+j6JoWPbWp0A33fav8KVOhvmm1TFRXmZQhABB
KtO/Wd2zOXS+hex5c4xPo2TBL61/1TLvJehW+ITPiUOXqX8cRFp23t0GnmqwvywZ
jtqNLcNc135BSVbkbRCLGgc8nm1IkV0ogD+Z/ckIWxCGlHYa+FckSW6CfRJLT+Ix
EzX299bVy+Dz0NsYKdXqsuAaNHqnAGACsTtusIntFihIRR89yuLFsv0LYqUmhqob
mJ2MwCP0asy3jyHdWdkeW9KoQmDsizZ27On1qUsrFY6djc8n0mMRoIhGVuLbOfas
qH94I9D9jycdr+rh5ucutNEMrHz5AgIzJkRJnF/IcvZQ8z3VON865RN5LCIl7ppY
Rnh/T389PtVNbh7aJxKY67BTeM/1MhMO4EhgaxUM7kg7z05VTZ71DxBEgrhc2mZY
Wxd9rF11JVAyP1aHz8ub3rxk0x3IhyeT51vlAOGW84S9dQ917JfgDyfs8q/Dwe/g
pcpiMtruzrscSsdqeQG3ERAyQZuD9faN1kzr50FI6CaDimV2B7nCmXiQJyUnLVj/
C3Jzny+4+5KC0encisJD0T8uaZCOFZKt+0s/PsJ53jIy/yVrCTXEhL7e7jZY+Okn
DdNLSKwmJQXbnB/20YBF6bFkRYi9L/IRntq1IlHM9L7g3U0U8KRN1susH8ASSbJ5
UZFti7ZwVWLRB1VFHWqHcW7UGvbOEUtNcTVDKX2uJ2xd3ZYI/2NKlH+IUBxmwRnw
7K1IVhGa65x3UIZKdWS+KBJKkVbrnFLWoPjlCyIcLKAZrETrp5gIQBn4fAMUIpve
2KO/3MMCHroo/UbW1SN0wU0ztVbza7/XjSwxzpM/LntqWrUstiANgY1Ost1QTG9w
/tqQsUH7vtf0Oea1mg0JqmAMJIe0lqO8uTmhnXvWUDrQdE+2CWdD8CTPqGZGHEnn
dfOEDZaAGKImq0QivBzf6PN7pMupPLoVbYWqMR5ey/VbuQYZIC7xtgpNzE3tlwmL
lOygWffDVQNsR40pZO7dGZTOfmm3fcBRoCI+VBJk8qcjQGSIemfMOeAsEbJEtxDW
fDNQOM5D9xcW9ZA9dG4WxsCqwSsvjDojOyUZlXSvuOhZNvVQwjgp9j7eiohiUmO3
vKlX1y9ZkckDuGP4uEUZcXXIF0W4bMPQxj+bVbHsXiQ+dL+5ktSx9YAliYbxbKFt
zmwCdxEQdZ7KPfOMAlnyK6jIkR13/1hFk0rkxeYHeyBMGwqxpTGC0KwVOvVK1rG6
PXwpxoNtHNyDxuvaVXwzuU1D+EeO5ir9Yhd4iA73jriJbmdBV9OL62LiRNniMxbR
B8kGxTxDudc41B3pN/v6bEvWg3GAg9tnxaMxwkfpM5hGGiQr3/Nm/A6fw+i2XcxL
Wf+9l3qJaiwQjVSWAPpDVM9Dcb7Vzg00XDv4pfoNMvDYeT6//SOuMHbx+yf6xxcy
VH8jR1Gw6e1G4ica73ArUxi4HM8vY62oDQP0RQet9sn597PrSCfqfqYn7+Teco0V
flNfVj26DeUK/PyN0yF4wlxh94+nl5Kcp22e/aNO7OrFUdCOktwdZ7lwBcs4RQYE
YLvE6s/wB16vbakNK5l1f2ziDxgzwo8ONhFFNjteqsVnE7lNXAsslKUGPuBp9/ee
DQ4tweLNkTXdXp0WEh9uuwz7SRrhpFU+dranKBEurT1RelJPJ6VPIgtIlJwgxhGL
ZZlaUH99wSUlLB4o3JFnbgyEubzEmd9hZMotWLOtf54T+LpPTkwkPjpX2U1L19rW
0TQwWR6MTwbxapLyq3T1KZtYbXQ0j4VWijthockKCVM6NK2ZQk2MeYcc+Fh86il1
Ffyj3ahGsDWF2KkcFJlb2kDJrQvtKe8tAz6I6MyW2ORtSs/drDXOMYtYAFbN4tvP
ebXH27KVk/5y5fnN1ueLCi/jXKFeU7vuV4xYCDMLCkND6oSAJrS2iu6cst1UICa+
4o8Uz5q1MWFaOCSDS7XWl5hLrxq+OAy1ffxOy4vbS+3yP9FuOooI3Mzv0+9DAqFx
GWX/wB+qy0/URvMAKQT/cEE6CCunTdNWvg3uJERGQomvxtLig9ggzzGTRAQLsYw6
ilAEA7Q2JrTSW27VrophPznDmcwqSoEw4cugzQw5CrxMXLumHM36pDitiQZddIiE
876jm8A8TnqVAtZ01q85rVdtOaQlXXBvwojayPvvzt7Puf/XrBzk+ClMdqJ8649v
YgzwO3Bf1TvZJEKkZBKMndND+WpyBsCJEpYvOhJZOq5UWmmnmFQJwQrbAQByrAAu
yVsj5D26iLDhPuKm33b5K703UkyIK1jUv7bKdPK9iWNcWfMjjRYUMUHZSII3GTGG
6rwxxdLC0K+jPb0Q3EKvrO8Teb6mu/HR74uhcBI4DpHeT923h2kzNtBtTSoaXa1t
/SISgPIgMEqeDjZ9vV7jVOEPC9sHu0zuNNPfAFFUrSC4Bh0yJpkM5CquMQFbSrx6
SkJcGUquZh7YTu32Gc+u6GUOWufMb1wbvVcD0R1kh+skV0ZS5JyCgblc05rabqtS
QiPt7ZB3E6YrGVIck/FtaoQbceAuX7Jv+MxM6H5dMo/ixGfRl1+c/aQiUzS5tgJR
O6k8el/ErKUpO9Qi3wNnKbdihKDg1Szss4H5yfUys6rAs1pFxwGEdGi1q7alrb+7
VJcBoryBHAiaf/3TeeapA2hchJEQKrfFA0xOC7edEC5XcD6rO4IIHQ9yYNFVtaJ/
N0SLb8ChUP3WBg40Q32hvi3QEKRqrRADkRo1qxUSmyQ2wIn99zyv3TjbG9x+Rpwi
Unoe+xqCQ/UGRCYftnlZrA/DYeFdJbgiPQTzZXmd8FpnnMxFKIw0bvt6k7bC7Uvn
YqPrsG32plb3HVqbhYHMkJVuLtttjevJVm8oVlvXtZ1Aty0Ag6SQuid/+jrEHXS2
4dW6MohWvywy89fLewAdhQA+K/gy3HzkrP1kDphQYGcenVelfxmvsdltjrqEGk3q
AOg3rgAq4RNRLHySLKcJbA+tclQyLF0Eg333aB2jwgvaTHNUMaxRuNohmmqNqwa2
300JadFpD1VeqzdzrlUqSfeVYtSZnnLq46+odzHXfHJTdU/RqFhLzi6ftP41++8R
3Vukv4Jroye6gK0Yfk2pO8u3liVObX2J9/YILmVu7lnA8wpboEM8E8TGy9+iCPgY
Jma5b07KdpIbxQ6Erh2VKXkT2LEE9ylEOG1kzP7oDVtOvWLLY5IHjAeKAYDoB5eH
+aB7ecv6Zo32d99Q1VbJSlUr80OI6LXZ5Ic8Bm6kxCfrNvfpKS0bL2xI6pWjDvpM
h7VuCNEBX8CD33GmT4HDm+pdPLU6kheXjoUjqIO3RyggVrBc/HUKBsqr7PstH2lo
f86bvuZIvHFbIJ5KFbgTWdFsQrNrLxVaUj4pfH444VliAYuoDF+ntOaRQsCZP2gS
4kOru1PqYEpBdzRfu2Q3KQEjCpx2u+CfURXROLNqORxyC/+Sl3N4YjLpwBi+VAZK
XNJCKNn2/J6/wxXZbBlLNQFeu1lz57Kna8FeTrVOKChlBPjHJX9qEWp9ZBC9bE9G
u3VUnDYHKe25kcS07Pu6fO3/ig3dVMYfdu5w7739G1xdXQq7wDivLc0TeldiLNSY
Y0I6Wcw085FNqqfNvpTPryKptAaM+g7ts7nUS90KSYwcqghQm2v8e9wkjhcCOkM9
cvpSXeVWrjW3fzJCjIFvetb7G4noNlD5V5XbFWW9VfkEfauh9VlGPvUqx6y/56Zh
jfUhmpYXr+F4uSr0M4wyW9tFVw+8o5CfYDwCkQ8eq7FH+Oq77rllPJSOPHZkh+80
9yr3DRZgEmT9mtbRQPXfOU6x0qMZ5SrVjgngbl/9NVoxjGLTJSjlRrbNt2d7QMtd
JKYO59i6jd+Rqi1mZnpG5a7aNfS1teLRxU4Pwqcx3cQRm6gRNynODS/nJmCW0p+J
hvmyPipZYelM7iJR3fLgMy8Yha/5jqCpFlUDbVhCzCyiXIdEmZ0USMG7h9ODKeRf
vgPtalTZghYLCymKZmd5Adb7M7PJE0NCTIjmGrnglC1WxnKDViW5/hlK49hk0YCB
YYuRB5N8LGTUhIOJu4SJkq/GUdMOIvjc42cNRahokmWajVYNdHf4szy8uealtd8s
WYgvZfqA9BaIrhhcyWXpTH7pv1W9J4s+eRK99fhPA0SwYBNFaiWG/JSoKk9kMSRe
X1CbVIR6GnGo2fkSQ5dQSQ8diQ3ET4asRYSHZgpGOTi3Y7K41KbRjWardIi0S3bx
UTjxEQ4EDu+RDGrxfaxziA0LF9NWFOmxqChK/IpB3FKvuMLkw5z33X3itqr+cAKz
3Y6nTbHtxDPNY9dLGO299kbherJrAZzcZROcyosdG2uj/gipXzneYl6co0zQ5YJv
m1xO/KsmgE+q6OZEAo1Qk88UopXxsH8NnKmxA63hTtL4IjjdSaGqDigantnAArgm
fwM7NdVZsBNoDTOziy4YBv9B4AcNJT3OxeIGCVllPlKOiZsr2sD5fAdMJV6a+U5f
sRPuQcYGwB3m5a2YKrFnWHPIIz++Ff5f+fQEYfvh5Bf6Y6vLzpeQMxgLrsTkvkW0
v7IbOEnxZBFne2Ood+L1YKfa7Hh++DE3KLubCFPdSqX3/DUuY0YS9CKkPKOp+OR3
CE2sK+78cnCb054JsUM5CwSRcY0MOq7hq10xZXuI8wC5yg2A098At/RmNy4uTvl8
tbonOh7xUkMCje5cILcJoTSjhTU/SvFJCuWbe8iDy4g9IpTB32FOk1SXZmBC0era
uvE9PyGusgrN6wiALXPqsace1GVyPmw/PVEtgpePaMAFXSNVevfWfld11tgAHYyC
bwAagcS5Ry46sZCaxSZZ0nRPfOpNkYTZPPdZ9QtMQqvIuJeY1htY72/XUB45e/gz
aenn2p779aGx6f5PSrp2fpna2PnuCYtQvL7lJrgWC32JgTBsNPx1ZNTH1c5m6uMQ
jAhvzhoT31G36/0j8/o4gOAbQ/pRPTliP+zhEVJke2TQDglHcn7TJWUMHjy3Jp9I
O+11z7hbAEorMczbQPkNiE+6rEVmz05cQuSCxEyRGWv/U3+xND9oJt8G7X8cz4Pj
ljMd00PizRFJIZxacwmZy3vI4E6QeWG6llwmZMsu38//hc4V1FBMFZaLjtdaEhMo
DRVP6swDpaWcmf7PL/sDVaDCGsbQsISJuQt92VWQuO/rNmO3T6+icUc/EoG1iF6k
KJ/t6CQ6rKgpbqNE2NfN7fh8Q0TLsvFr1UfCQByTi6v/4baznQ9ujngZDGcdtUnD
HmviR9SNLEzK17pv/zO9Dh6DSchVMJ+cZgf4ht8oK6xIW7rPST3Uppe5soHtdUKi
Hm/Zz8uJ2qg2LSEVHbYgKR/ZJZabXP+xu/uky0lHjJjQCVLcbM70+ug5tiW/UpNo
HTTe/1GZJYg2Tin3jCInVO9OaMdUEqxDIBT8g6vw669qpRUTOWwFOLto8SC8A4V0
+8rDBOB5Xmd0mtjHNpoz5Dn5IAuHjQ4bQWFELwWV+cx5B/sQymWaYObs+HZZ3mvh
2tR6naxBxADS7rlX0V8UflqtE9vyX4nEYclos0FJqG+AGhUfzvFjrSDmFuv2k567
jxR6XLpKIMbeBF73zO6R9Ni4cOGagZWrzms5alzL1rl+ugI/GqMIODuGTk9jv7UP
49k9Gy+7G/zM4e2BXuZars1wpYwngRelY+PYjyxFNtTMP735+jo64K8cuSGGZy6x
/kKCZrNpqo4PL71mL7amkU8UzQPMdMzrjtkF8lhNE6hdPiDzfebxrKZzgfreayzC
iN6Fvh1wfJ2t75ip+xikHB/QFNm65BkPAkZummqfLX+68g6ReTlPG3efksRLE6Hq
Zq57quL8DT3w17TOQml5DMwW9dxtT9f3fXzAJ5cYNi155HtuTQJxBkP+qyexhUbM
aWrrybLXn7Ba0wMHhKl3uLZxQILkQLSyQ4vTBRedOR8UvpeeJmkLzslzfo7ruAxI
f4sWecfIUyxYEep2LTkASrz4sIfEJzHG2HOLXxb5nA8pKsRmX2PltjpbjODV3td0
lqdXICKfJBXcUeQwHz25l82hdO1rYsXKQuEOM7qWa8RmQKQiW1vDTQsZcoNu5uZB
Hd7JfIzLTax8PC7GasWZPyOHYbeB+Nw8NQ5RttOb32aZgkyYbFAnDQBC+MOssxvt
CjkHcWxaG64TeSxO+RlohpDDasCTWvJMZJjB2k7WRNaain+eGZ00ldjNLMsogwbX
TCiHKnkqOWPIi51r6y2LGUTZiAWPPSxW55Pa31t2WTX7Zg2WwdPtFOkdrQicb5ks
5/0NaNo3c/lapPTBBUXNX9aUHpjeCYG474C6HbMwRwJYZojcSo2USraMizEbhvAi
nS/6dtLbpfF0RaoohB+1BYoc74I+M1vT1lO+7sQh4lFKVK70u1Uk+Pza8LjjJOFI
OI3n/ijm5Bisjh6oALln+AsfsxBKb1uvuzs6yokwCScb18NDr7S73pntP65x/Nbl
uoGxVixll/9+nnofLV8UHn19xMrQ8tzZw04j2vcblGmfdtlYJvtsO+t0+yt3x3kN
1C/EwUjH859xwrtnKsnQ/aJ89owggLCy9VK7R+7aAqkzArW2sibW6Bn1H4neHL2L
NcIpRoBwhPYPZYd2jVFWYgD0xjPGvXIzDf1juarFfnt1gzIsR0AY0I93H9s6hAos
Rttasbzj8Z84NWrFC6yMMarGpp4o2CWADTwQibT7xNhwBtS77/GbtWHgwHJ1BQk1
r2pWW5QnPczgYHm7gPy5me2vAEXs3oLkHAACm3F2azrdRHTm40CXyjMRB4sOD7pJ
+iytYzWeVMHXte9mgXVXjn/9ikbZ9LnuAXTbR7Ox9sB70V5Aaiiq7ll83lGXMvf7
yjuUYn65wzgoq/Jqw3reAheSiYuJySEerfdNEGknlmUbzKJk8VLl8+Nb83I6XVw9
ypQGOHWzTNnO+vamTclbDUqaN7/4KXzubifdtFIplDgCahuhC+LBTsQQtGC4qnnd
4GE8NJDMOxFqIXEfaSjJ2XvuqXmVmGJam5VG8MF2sSbMQwCgF56pLrBw7u0EtXSe
uWQJwngySxh1GUMBdQcmUDewUwHrPRuPu69LyjUg/tMFCq+0Co5VSRjtGJOhfpwm
PYQk6xm5C5E4vdHxMgSaOGFyysUwEUSY+qJ+DXLTnpVDjeJP1Ygdyovuypcv8iJ8
rVMaw5N9O2f2mu+T4YjbpUzHlNMErOat2KwHrsCSUrOMyXCBy0I1DsMCf/erTVqY
VbQzyAV1KO8GXp8rJJDiEk0ASL2yjdFXJ+rS/Zz5UyEoXtMVS/sW2iRjj6VmPnRq
wzxROsU1072rb999b7zkf+s+oy/YIAj0eRYzzGO317lPyoozecBB/MV+mflOcVdj
X58uhFFIQFlXJTaOE8/RLGJcXzv87RyAZkUJZg6TS42VU1jdZToW4KCOSKkkL6Bc
Amsg26CD1/CpEewJ6cg2vO3Pk1GCK/Vn3Zx+ejTggn9s7oqC8pndVkPlSFrXqp93
NIUBXJ90fUOeo+ijQ0ALeKpFhnAt/O4cweL4MDL78SLyYM+xlyLdzNFR8hcwuVv3
/G6bhElhSxJfhqC9pwnx0rpko9Dpd+i5U24+kvJFPX8FpO/opxLXq0cx1E2pIozD
VuatSVnQ4BEIR/xG9FTk5Qhxpomvb+izVkejZFTFvgwHEG6uTAn2vewCXM/E2dyA
ZrcSaM/5DE9FXDPWr2TpCZhyUG4OhKNA1RLHGZusV7RPS6JBiZQ52NNi3+CkPBVA
O4Z2hGHyNBbG2Tu8s5ii2fR1IzyM9Q8iLoSz/B7aejaV4GnhmfjdBfYNEDgfrHiV
D5rJb8mlQhQJA/C0UKYNRYF4cMREMGIHEBj7fcQrDjsvj3Njf9tZ/wkc7bkVB20E
41+eqcnElnGsYk9f6yH9Q/gESIgPJLxL4q9u3/VLq7KQ4eb8LuLYNjT0vlKtjsJf
+BqIW9AFs3O6KQToVeL6YvE6ig0R6HhIPlbXevbMjOZitij+AeRIAoaxkvwKXBsO
vUA/bi2xD+Tz30/heBhTebmtRiQno0/HJRhTkuGEBFKj9T7cioAeXzIpHbmBrNIW
3oyRhx8Ob4pPGfOFOCQ4ROP5BzF26GL3NgrRXzcIJNBJRJsNOWiR81n99QjcqetE
LSLVee+fv8n/kTmmPFuVvGMQSeNZID/WWNJnDDtlwyIvvnCIjMsrQsOI6DfX9zsT
NW6xsdsjNy/azCLxL+/frR5w9XfjpzjcFexJVTHV3/CmkoHa/sTfaAeC9OEYgDI9
Gov6jLTo6s+QXd6wBxy6uO//bmEqjBqDysyad/tC2JX6aCNxNFAlkUyTn0U9WT7Y
YefPC1Am1QUvd/Tg2NGB8MQ5Ao56tmNgXz17S6HUtKDdSfIgVNckklYx6px/khkD
ubfZyi26XfwXicZbG9GWq7NGJ9ZxRDdvNeYweKcXLTnAHPhuxa3yqgovjfts7UgA
P9LQiOhmgIBFcjBVDcDPihGGSrLzO/q9XMK1LuCQtAm3HqA/7bl4Tobyc8o2K7CT
xS5VGB8pw1a324hX49B+KilDiRtX6cEgfjHQCck8Of9ZBP8FuqMinvSuDfXtcSZf
UMy2fE8g03tg/PRNZvCxARP3dZPDuR9ps5G4wZGDnPqVx+EziipsJBfB2oHluxHi
ZKrp6gVFKtjIFpkRhZcRwrGhz1uemHFdu3LMlEh9iMvdEdbeI5Ydk6eSe0baasgX
+WGY5kzQzf7bA8Iu2lGd91LJZMWHAeOvqkmc4pHn+4gf0D9Z4LTmWSG15YTITpWb
MuaVev9kEk2lOoC8FvFiKQjClLnFeUHwL3mMCPBsEK7bP7c5rSzxcE2vJV1iUD6v
8aY032J4kXi2geXhOz19PCMCuzou1QkNPjKAzrsmtbczGHikdj9xKm26QwIrUCiT
3JXHldq7C8C2Gp355UIGDrd79HjAETYmDQd1ZH4F7SKwoG9+IRwn+Alasdgv+VZb
dzP1uM+cY5BPth0i7khBMR3FPoIP0FL9esZuWeT4/dj4gj3DYyynHQQFHD2Ryhns
em79EmOVL9GyoJ5kcn3X18uXQzeor5nAY3ST80q2jOffJvlmFvUfCdoNFvnWWOrd
sEnqdFBxbSDbuNKiP1Ix8ELOmFLRXzO3ouFrdRdq+gOtZttaeCQC9Hc11XtL8+2k
nGaZoE4WfANz+VtUByE3c+q0YWbL+Ce6fDFk/63Pv+MyWNG84FHaxVmrI5UtFPvu
RJwzImlDyyKpj95Xt+YwGjx85TveMMoaVffiJmrrLj0IZQqYanM/tACsQNwdyl85
G69XHP5N8Qg/zteIZElYl1ZVXB4MUyXjP9rzBPy9dlyUsTHyLVpsGPWIz0+tghZf
8FiSytQPuOTR56TY+tTSz/KIDEE28LKXUPYIiWkJv7hj45/Z90y++ln6e57vyauA
5Nk2Urkb1/oxvBo0b7FFQFF/XRzPrvWccAVa6t+9Q6tJ3qYfe0k1NAyayEPEfILq
P3afRARTy8rk3ApX+muYdRQYt3HyyMR6pPJ9BHyTuckJzV68FnV47W5CPOoJ1MBc
D5Q3UVyoVn0l6XPO4dPoymryCrWKiKDcNDc20z6z6lgKo+E5cJyBqr2TVBtdKRu/
WNo/gGjKAZ+E/rNDZpZC7HNaT18RE5nirnbrtvbvJQEy54QAfwokUR15DGYHujot
PDXUxn0mQS7SuoMaLGfVKC0wdIzjqRCbfvVG9pzwV/u3Aqd9cnKDAdpoShGGPtMb
B4boBE5H9i0OS9LF7pE5XXaMZ/k3eXFGReSD22MZhvTx7gzlveYjvsb+SL7mbLFt
7pP6DGLJyDg6+7dlGOso1qZrCjoxp0BxcqjPeYFCxEuuOgM8sbahyh0sQPwgb36Q
ICXOxUcIQScS9XLg2oZaQS4KZoa6sm8btQoZNGcbR8fcGJzm2UjXcr8QSJ0xwaYc
YDXzgu1B1fAOEfhmeaK0ixzkxyNSXS/zE0PFhF9tpv5ukeAOs1CeWvnRdbGAMeOf
B7WNzAw0O4FBtUffohnpawkVVry4MFmVFRrYjoRGs/nNB98VULES0efYdhKinevs
wwW525D33lQWHzdPRUuKBNQSu7IFW0Kc3XwMov+RvI7ZXISJp7r6btof5Pa5Q4l8
m3md0/I6GUzfwFTrH9BDxv7t6I0uJgPs7kVX9JgGYnQZqDD7kUVm/BviYv+ls7rU
B9pLsb7zMDD3h8RHX8/wkOlDShtbXzGEHd9GyA4yA6AKN/TmsG7L2a6yBTXXcUbj
NdgEgtAxU23OibDXQ3hoSPuurNaFynlGdPw3M9aUfz4Lm0GZhW4VMJuiUOhw9Wa6
Hy0ScDU94zaWt03XsILfi+67Lue3OhxSMKEiuh3XWUzxXDilJngCYMAF7NZA+mX+
vbmUhVLa+pd7J526t33yf282dY8dcqhiE2oELhFcpWQmeZsF0vyD6pDWUfRVkZDZ
WJ6vxHatmZRwZbhnS4Oh4wCF5Gr40xVx443Jk9lr7AnN0HJ4Fq99a0H0W1HzNPWq
wfO9wgfHM44d5JwVIKcgWsd9iZPeQ2WS8zbWrY0LPvGzXSXXq6Xb5lyFPmLVVEFM
hcYCD3XZd7/SMP5PS3jBMTm0C2nNmywgT04wIOtNVwG9Z6LHLX/zEMIzQ1AHLk0F
9U8W8K42JvFvUQQ0FuoEy0eJ6FzXfjo/Q5tlod0irYw+/5scHMEh8yZG71U/cDtn
orysvsM95VyihL3XCybXNkk/drqAJVuhMOl5CCsK64GXX/7ARy6M+Y4I1PuEMQu0
NtSKGl4D7/NkA++I+c4TN1V5SIL8ZXYeaZ2Szc2cvVuX43x7Ruu25V6FL6corOqU
E4QS0nrLKX8h4TtZFu4LR3Z2c4vKg9xGOXRDgkAL0FnvuphUiNtKFH/nuDHdd4Ti
6tqdnroES+KN7hgHgWW/YsBB3wzVdG6YmGhy4MivDiXYeTp+7br97PLviaLbV3Os
LX12CTQYHURZdawhx5NPvrWf4CjERHtpzo/AkFaX++ti3N0Xt2z1FTLv6SzVolUp
NnFY9a7AEN8758HMiQmJ/QtZjDH3+DUNfugKPvjEsEuS3gaEqibn+YeItpesjTp/
mkCq8pAjqsy0LCXT3tncGand/OdTCXTqex5FEbfAEglNRRmxeKjPbX1LARBSzSMg
Rs1sdepSg2uOL9NxByLYPA5qJ5KrVIOX1CIqDpayg+Sj0dP/UM2Qr+VDzunpBEKU
oNQUsRNQwBgiCTk81+QKXYfzNLc4jhfFBjfPUDOQOG5wdl5VDbYCrhdQIfQXO7k4
rEEBVD0NybF0hj7RPh3q2wIFL9vTq0sGK3EM7/s7bb6rpJb2ysd5gCh9O2+11cmj
EBXsoA/Vyt980ilPd7QH0GpP9DDSgMZwnnnMLFjZ9lJrx8sAg5SkzwIP/UwDx/OH
+KTMoNbO4O9GpzilMRIKCldBI4L8Ute258TNDHXxVlraGGQtIJ8+Ox8h+CZLr1rM
VB5HEUuKcowh+WChJhQHgrQCkON3KifIiRkVNwOUJY7VMlrlrFtQRQLv31h7Ujce
NZNaQe+YFnP39XV+TuWGyGYPA+FZcktDPnWc+W5Dujwuv2pqwd6/XduHnFZJ8c/y
iuaqolJJBq/Uiw6J3PbLVl32nDG/4YxW0bVSXXPhSPJaCK29PKEU1A4auOz/xjnB
AwTkac70C7602spvr/FlJy5GhrPk++898tDdd2NXAuod1l0l5Qm9/OTqOD8f8D+h
NFH+n5ddS7Ry4HCflmospuYEDzAS6WPOHnjiPGfVAkI41IWnLKwj6hWR1emgmkto
MklZLPOjfhmQcFjymGHUlIwct+Jwz/Ha2C2IjPYmONQEu3ULjiYj4z/J2vquVRlf
AMX3MJlf3fHRTeHzKQ+57SwFSq6yGWKjJNcuswE5PlVjEMpk3OE1gJNED/hwprDy
jriZ2WnBesfrR5KKy3uZ6AO9J3mL3NL/vY54s/uKRn1phFtDsrsGDJt4qszVVuLl
CK4XJlLo6Gw/ntBrH9ObdZFxhVw9G99tPbRHhaclL10Zg/jKs5yxDz1syDXRjgWg
4DXYiej5Y9LuhoevYS7YSJLfLnR3cfWI+d9Eyo3fMU/Stcxu977R58HHxymbFoEM
9tv1s1phlvg9VbeeJpIZmX0qUOrFdUop20YigCYKA1p+y0sEIOW6l1CAlVaMo5SR
DHYfGp734oIXpvEErchV4GSlPer3qJdqZmgi11MuOAzdIe9ZGAXTiNgV1IaNjmHY
Q5+dc6hTf2Qm7z1RYfhIanwEp5zc8uyZFbcjMZGoE9FdQyvhqdS3kY25wDYQ4fFF
bQQaD///M6LQTYDP2dexiocgnmchYMv946WQF3c89ByMd7o+K1zi/AJXDnv4Wegw
gr3B0s7apD4LIoEVXefW/jLl4XO+FoaVTtjsZTjh68dq+B3K9ePZJySCVGxKSX4t
/AzLj5OJBUUttizImPgTtoKfy7hjtTibqtED7bC27h4BnxUg/roYNr+XKXYDkWv6
xM4oeQJD46kj8xQIlpqnNuKT/SxL8oFiWOEXEDCsaRTQT4If0sYNIOruDbvJIqT4
9CEPja2p9fy8GzzKel9yOIhI6ICNksS7Jy3slMMJUJcG5hkTEoew9yYJ4sKLZ0Ve
kdMeG/2KfmZlznwtIBEhIuTJNBPExmECMwjHDcDhQDid/6zUjOL8HBAx3Pwraxa3
Cj58HHCy49CotjiayRiiA9mEof9MsRwOpFnnHwf4kK894VEQuVoN/sBkUrcDqOg5
H0WP9DdnqhxKhAw9KRsL6V9Ra66sFRCcdtjmQdXaQM+jwkXQoil7VDOFx1fLYd9O
/n8ZtGkpFqz/e1lCDIwYXq+gB9W4OB1+0v0EYKsTbYY8TaVWMgyIKAkQ7xFv8BcO
diomQrIldBJasLfHcvPIoYGzvwK24fKce56bg9bocIYt+xlyqSF044NpKgZGDdXF
Uk5bVbPxSxe1NSBBwjOjXzcyt6DRrwKNDj2LRLOtA5hLpAUGMIEtKeh6IG0TKVZF
xiypuEcnQqAin/nkr9+NFPMWH90E9A+PP75e4gXLhPCj2fiOV8CuRcu2Ryqy1nVY
o4Osz2zGmP5nbEVzf2xppwplw5mz0QubzQK196DKcsNfSfcsZkrwpEfPajKuPZkC
friywiYNXCcrPCM5UygjeTxhFvnSM0sFlJVm/qo3QHtLMBErQDLyvEWz8wj5FwxI
+rXvo0PN5iMajqv5luWJeAkzJIiqD+vSx8epmC2BCvxjYe32Mr3Cvn6VOLBIe96p
pVy2k4g21FUnH9GO/wKsI12l1lRDyesm1ZYIshkFrNTqjeFQ/juLgSIPfvuV4SGc
/l7JDst99Y7dS+UdNEmW3QMgYU0ZLvDL1qqj3J28EcX0wkWwU4KrZQIvZqSBVPLq
Xw5yTSRCmrXCu89lXSytytLihYJXdR4HtTKFzX0gIhEvKWyg7fx6joVrGHI7E5+A
xUD+FwXXGEW7qfqwXbs45SFdlETlbr3UmwHwHgsJW927VIuLPfu/YF/kDfMp6hSL
m40UofIL3DO2QmPw03ADzYRXH5lePlaQ2usXkty3qrookISOdXR6+/Z/gCuYIqaN
HlwK19UN2Y0Jceterc+QA6wLO0C8+f1QMZTmFGEkExmCoLUKUxG+aXxIgpafICUi
SzKIbkZ/TQznCvTg5THJ5kQl3Y8Y/GTZJuTwvHDFvqRxk2zxaV/gaU5ZIz0caQMu
Hdxm3efVH/fcbVc9AkYoxGSyYTXL3OQdQB+aQyezztAq3twSDhGRT/RDTIQNQ/gk
/eSiyn+0pRH1rWPJwQ2LVOGxraymH9UXNj7HTMdmrHD2xynfEjgV5kGJpJSjGixm
j28FeIFaPyuQjxEzuc+JF8nGl6rNDAlOGEvBp97A10/Cu/+Y1aII5C8Xamj07dbS
2bLuo821dfyLcjRRFIbYyn+5OXpe9O1+0zV4ud63QSnfI0wPGEzkmaxSE6aHKKoN
Llg67vub6DlyDGiyxfJEdt+CT0d93pciEThRQCVAcJ8Kb/+o8VhxlllSqEl0XNI9
j+wPsaKVC8HJPnc9O7qMW+wMMLAr0Gts+/9fSxB60a9wvXitQjWjiy+vaCjblzOU
aJlTv/qY7c+Fojv/JPmXNioPBnB5LSNkH3frU2u65uxD3N7+8iBclT4425N/ge/h
yIbT6I5ZzphgDAh58w7+68J2uaqi8C3wJIg0FWKb7s7DgIzj8Mz5XNvcFm230Div
53gMmVLV+rSvb3H6JgRNDoCydLKDf6hhKnDF+Y4qqkQvvC5qWMUtbjPTRWRmZ0JC
hXRU5MbxKHYkeKlTroMZkdcYAKobO2F8IWDTh4Hk7Wk8PdLBkUb5XcM6oaC3XWJY
S4ET2gTxHQ/L3B8pTeLC5t1jfxOyGOGlaCzG/PsbRuYdorpOHrsxz1h3IMgdFluZ
AB0pwZVY1loVSyI+Ui8zoUQ2XBJXHUGhFjLDYa1jSe02EKTBIE7Rms1Hg/1+8kbK
PtFPIzWuCkszs5HmC/rkXzM46I963lwdLHLCYiCrOKX0skzZTsKpcDWYBQjI4DXT
yQMadj4QSFHEilz5H8c6LTgtx0RAb6jMumwNRGKi7SCYTlFemfLUkcalTJtPpvkX
oaObhtnaFN9g7xZkk7ILci16HdePhkhYoUJErCzYOEA9t6J4RUdhmD3FhH6MrE+e
6B2f4J9lnTYwkyCf8z6YIGyqUt87RhWPLRR9a4kQ8tgghvrGIFxp4fXo9mSWvi5v
DRzdx5oLvJTUQzhsgMbE1u6/pMoZAmHlQaD82gYe5gOp2yE2jtHxqSiJP6HHSgzv
Of1ZkZ1zL7jhEcKcQMpaVtOtmeyyiRuzzavZOg7Jlr02Z1wqlWgAn41hiRiX3vFu
cYbWKmPkQ6ZZFjGFPXEgyWgpDtTnVulfa3smUDJyCJmOW8w7B6flOPGj/rl4zaQe
6l5YfRufNa3wl/Z3xRkG9lpNKC16Fjy+Jdd/kmcK2+91gjxkxKEu8rFT3skZ6h+d
SHHEBB9/+lvWT6TZhmnYtSA3exLL2uTqMU1coyrb14sfeauaJTn8aN5Mcg/2UUB7
tfI8A0jwmU7H2bbJRPrTunlR8tMfzrGtsp9uEUdsTQNqLnuV9rpccb+GBwcGPB/d
BR8rYP7IRk+OCbfSNHZatf91lhyFmUYZQdhrPN8/drDq5PrqXBkh19u4NANaLgJr
Wf76WU1L6Exy3OylOCBocu/SxYKAp3FGWDe0vDF1wVupfy5uYV1CUUkWqHQhJHBR
rscUMd8Vg3L4RBpphXWRcrlyY+IL1AVIBS4BGUxinhERNNbfG9QBSsPKeOY/luGo
86Fre+R3jeY4PBlzTIMhnIAcPqygA5p/NQyULglIZccfovv1cpvjlGs0+4D+txLL
MGMQbAYfirVnOjMGNXGED0f+PSA9X+GvOo5dmn5Eb+g65wUJcVnAcP9Dt/fvKWa8
DzctOYsJ5FfimibUGv9KZwpxz7wrNQ2zTaYc632ovuO8T8dp9oY2AMCjqriMI4VC
u9B5NdyE7hYUowu3zqhlFrrqroZBZL9apfzaiS0LYLdVNw4/QtniUhnTYyp8LOK6
5tf7hSjkSJkM/SSy63DYPp0HACGMgTl9yELWRWAboCWfI5nCdTMmIqZSVcGi6Ili
pJhBhQNoYFIcPNd5cgi/o+xdIdyXIneeC+HXuiT+SPqeA/QV4JOSI3+MmGv2Txgs
GR0mm0sGpq6nfedj53Y4gdsB0w20hBW4M1MlqfL7FGQ2vX4Aqx+uThYJUYT1NLBW
jw6Wm+wngJJU1zps1GfNKyya9zphG529EMt/gDpfyn9cJSBD8Udgq/b/8th2Hm2E
UPTZ00y/0FI/hrZO2ol6N9gLdZPB5PRtFhMjZN/lufM6J9kDUN+bszic/4cZ2C0Z
fni6BAYCDLi0sVlDAqmjGiwiAUZjNkMunItrjR73wEWd4V5L4h/2UkGNp0FtRRZp
wTtYcUj+sFLPRSR+XzXGpDYs0aTBOg2RSIs31loOuJBics+iN3Z1LhfBdgcfmwUc
2Q8jAaI+OAtz5VMa2h/RTC3O20PQ6+C8o5KffA9mXhDUIb2e4muNgUv59I7uESiQ
TNEJpToLgB/4MPYpqVspqKrSlBumNKHR6KynFi5cHUK9/BrVFGhrIdP2iqwpomaI
WHjEtlHFX4azRIs9pmh7HH84wWjSs74HGivDt5fZ32TpNWAWtHG/9o7OTQ5cvavG
45XioBVh7KhbcZiKqsX2OR29eGqrYZyoaVCeVWSyetSWWAUzh26J7sozdRwRDuEf
eUZudG9CABWNrbOX+2veK/Z9WIXHg/MFk4Y4DgSjhiDy9YsvZzThl4LOgT1QZGPy
jI67BlLkaWocdl3wjIGi9TIHgOUQ6SW6b3LtcQohv+qMXSBV46nwkqtpOKE0ptdG
8v9rxKsGZBCWQyg5hymC5JZeQKiGHcE0pD/oad5zQwyspI8QwZpiKMkesx9wK2WF
E1jYBj3kC5akxSJCPzhDdJy4yAK9kvgsSXt56IMuMRr+dksbXy2bEDw90lm7hTV9
kxouEPMuV6/9wSOZDPcW+gl1iRrgPt5VOroULz7JKokQEgkNkUWvoRGI5FY53TW6
1LjGp+aaTflPiYQT7DIvt9H8Ccg7T2fo23RwSC4eeUd9iI2F3MSCGHpxxL31Bb3k
B6G4TW9aEh899CXa7kHAyIYA+Bx3FpxCzSpSsi36UJQaDpV1j+yfVsa/0+R2tXHG
/kr9dkD6qsyA+MQ7tpHBtxOTKVRnc+awdDQLza7mvYQwNCuguhft7L7Uka8ISgCt
PTUG45OZkS1hSDdH6A18IOJIt6kC7ewAJA9fUB5SkbAskt7u06cCecfh8oKAjJfF
HZ3Fj0/UrAOClN31qP/vLDmJu5tvd+VNjgypWVhQq+0V67aNObhH+Sk0MoR0fg3K
egQTpQ+FBwcAM+APJH5ICldh1hUIBHgElI/B7lSpUT8mjvKVSspR62qEXppPjI1t
KX0UJHwW8nDNM9Kfp+OecWNL8vkzTCNEuJ00RFdaoFgyIkUOVv6yql8vYdotnfw+
ilu5crGe0YAuUBOXq5dN5qVXXgeRwAdt9gErQyWEjis3ggF7e6vtHh2oAfxCakH7
ayrNqE1XlCM80Nt7JoIJqYOoebqUszFyPQsrhyYyDTIpCKaDvGyxBmhR8E++idv4
7HZ/pDbZo1rIdbj+eRBpeNKXsx2kXYw7Bq3awys+1G93/fcpA4yEuOQWkTuiKT1s
suYwtk47lnEdeBDHL2hzIs11HOeybZwHhPvkvohhVKR/uacFechT2UoAeJY43Pym
IaLteyvXYRyckmpo7EbWiuhjkojY/kJcxNEgeo5wGmKVEPvZHqWE1H/jY0h3Lsig
kMC0xU5t2fgqzfP69+SD1Akh0lWt4OEEU73wKvv1TRcN1FZZdJJ9Fj+hYrFfxDRc
d1P8258CUIO7w5q4uCN6qd++VK0H5Yf0TGOaALHlHMZ56TrMXGg6tXmCLVGQX+j7
82vNpX/XsPtnXMRjELe1QP4vlyQFEVQjYJHOyE4B9q1MZEYsmMdAWSi+ONYVc5lX
ZzJZJG773DTk5n7VvDWFQXxHf2+7+I+08K6UF9XvkLT0kgJMOrPMy+KoUgETau67
f9yqf9S+Ou4t9QRzqoHywawIYEWhlOw8t7kmkaspjlAn6zKsAtZ/W3lb/WzTRq/L
dFIJzLqnJ54WbvuGWFyBF0+WvUsLi/in/0AzlMSSMg6GjSbN3htynyJgN1dvNFbH
Gf0wdw0K6iPHsh2n9tb1BxQXxCiWd0XuEQltAoFxRYzyzRrDSSfVEP33Ht+ff00X
lcK3WfKv5p17PoawzYXTfnvN+5yTyLhS++h/+pUhIreTrym2y0MhZfVW4yrQucV/
tHbyo9gsdmXe6mo5DstjnAXo8PzopOXNOhFHy1zwmaXaMql952WylQ/DbUK7Ngy0
leo/hQotBMTfyBglyJcHOIXQ+VV94LXrhaq3rXclu2NankSq1nB8rSqiYnw+gKlS
wQZFsScikcX0eeg6976Yo9Lp8k3qpECX2Bi+QBHuax8PjuNsUSbNfoiK8FkCIHwF
VVUtG0itjmKA+dJOR2XQbLHd3a5549u53TKj+CBcIFJsP3/D157qLRrVx/abrji3
BKz6pKJRcHiwspTroFqI7Jga79zdoMQAk+CPFCzw9TApyO0RnIjE+eP3WUrewRjm
nHB/rukIuXZ6LPfEtb8NNDsmXT3TXy1qjjQJeQbBbleRSPOGHrHeC3npwzsg/x/s
AUT+4Mj1R2JOB2lmVFnS8grk/ec22wWlVnTk6GpmpjT3ogJFu9XiHwQm+EONmhDa
OloAyOHiOI4TrxIuh0UdIRgPlVIEkjwjTIzp84n0X+2zhlkytBPL9encW+YwWPgs
k2dLxtIquG7bJRb85VD19SwPOROAfVbddg7DsezA3/SPWHR7ggjiPzVO0WAzewUk
59gdJLHuvlY3NsqMFu2YBGU5fmA1BgnEznmX1F+wZNOpItO8OQIyisIN5zy+NzBr
1rjrxSx3xOaln5UPOSz+g7OXMpvIOhLiibxc7Kb4U70lEfrICtORV6RidgGTw5GL
ihoUT9lNd8UDnXM1hl8P2BJdb3ViNUrX0a3uvq6zTvkgmDxxqtJSRnb3E2YfiOgb
6riSjJATrxIAWJy2X/KJHsIdRMOD/vQOjt8QhEKjhmKQazlXGEzbAuySh5JpSSmM
/FhSAUlBt/twY9VKahSLacuTbbaQXB4D8mPY1gp1iDAYpb0bmfwem0ThuEi2trDy
Jz3o1YYsRaaI93tuJvxqyI1tQaSOYFyKKBaiFP2iveT3iVX1kjoGsQbugaVBrFwC
S5ujkF0bf8hYKDF9i9WRo/LhgurOqjHIzto4IwRedqB267kWZZuiDvxiRqHumlSv
Rslzz4fFGWZ8lMCbV/aoh4vcUn3+DG8sWiIFQY2gsbZaPzmwgyKvLG9serbYhKlu
Kt2oRJVp9DSj4B4gTVjaOkTMzTc+hoS1NkFqg6xNjLPTJ96B9lRq6hCTUpDKuUkx
gJs5wQg6DxaZwKcZnj+ji5BZQPlfLr1CaU1F+S1awEgn53PXJZP7LrTImEL5lT1M
CnPfZl5kWJNO3atH0xcHSV2VibP7s3F7PCDS9VimhPNc70EnYQzrsTCe7/qyRtpf
e2VWaZfw0+n7No7IAiU56XWG1zx7PyqFyq3zpJ3v8dtdtD4mv8RjONQ065MMOP8K
ii9RUYy7RaSbr0Dt8/XpJQPwCr9g0RPz7dVns5GfY/8cJ0fLJvymLs1nilXs6AC1
EhRfToQLMGLFH4XBpZk5lWGOImQo05u37Bpz5j6OyJEIDluBIl8sLEV1AQvO8Lsv
qv7zMzJ+bxPb8EMgAmoY3K5U/tHZnSOKCAZoP8+9TERkSOLrclKZZcy6Cnq6vMAF
M8G3MT/C+49/lFa41iCgA/0LtYkgcTpp1DlYjrtrqCI9xFXTArvn2DDlFOUINUbj
LwTafEQ+ATOrL66P6C2CILX1eTcHyfOrG5VEOIn3aAF4rNDC7hvlCjyXd4CtLy7Q
GY0Nu92GlJfe1vsr/z+yIN4h9Aah+RkWA9d5MPBOfMSigfu4YmY1lJFpDbh9XlHN
IF4wD2Um+UJtc1AWVfWpzZU2qraOpNCyi4/NIEe38Ez6IPnpxNfcVf1KxiiyE+AC
kSn6+KO16a2a3b4MZi+x3rYp/UtM5hXhkewPweXSStwmausfknIqKkhfW9bfNS8f
EhjKJs2aw2z4pXMK5b+zQkOdf4Q4FAljlSJ5X7oddlS/VE7vDOZUX2B4FL+MLGtY
4lyHIQK3KcXBsGqF6jzbhHBwaaNl3dy3OuWdC8ukjCpzEGpg1/REtoHKce6TBYVh
98agNW1Ksy6YAB4bexwCgqkNn5hQYZKTIAjCo7paAjTIZKWExSEuVBD+wdVo6d3U
Vs/LkxOs8IwgO19umyBHzg6heFZIVnXPMkJMjPSygIiRnhCa87FWzpdCmIo1kU2l
/voPmM8U2ZIQlbIKFw0Oq6ajE6RruT29cpmPNgNQDKtePWTd9FFH3r0YkNLF4EkU
H/m0YvXkHNmofwRzq8z6nm70Nmp73C/7IFgODucNgYjCO012kRhHlZ8r85hq/Hr7
IbBYJi9KA9H/z3ql760ATXHrjl6IvN0qJtTQcdMnl4PNDifMTD2KMRiHoCYr80H4
BojyGye6jrXIXWdkh8bKfJlvek/nOPh3Fb2qHv4rJ6pbUxFx620Tyz6sTbKeIuyj
h+SJwcyMbyVmerZj7JqyX6FPFGSrWvQOMXJDVs7ywFByv2qzT2qcF64U7+PmKfwr
zrwJBoj1BToQOE04yMWjC9lkFfCGkLS/OBfNjIkJfD0x+XBYN/5mPVQdLMIU7tJ2
cpXc0dzSUcSLTgvpiuUHReaj7e7N+UZAqygnoe6sprKaEYKCJ2WBudet6QKxRHNF
K0boOaxYEjoau7IkKIMdnPN8p7pLNM+WZWNg5WTbW2tjhzonxX9x4hBCc90Tb0Gv
XNpMKPtJ/zvzLo9avwZJsidaQwHL0LnSrBT7m2mJ79J4IrrY2po5ezD9k9tE/C8I
pup1DSKkOaJtagPXF+VePsu/dKKwcR4nuCBfJ4T3smh8DvEC3giJWRO6+vXU1ZvX
W9uF2baRI66wkoz1kMFwLqJiEL2oqoHe8MAFKVmwUHDud5A6GbakwgusOigqXqa2
2nIqSjmL0h8tSbWqFL737X3yEjKHjS2hVjO8I9QVWhHPMBfeGHgHifFCGmRu9V5j
TIJ5iBe3eT7jw7+OP9sjKwlUniUZat6Wd/i4qojP5cKBaocifSU8QbwS6ltASGg9
bm1QpoiHCzQYD8qE/rppXUW176G/6Vnf3FMkppcQv6CBraH2osPPxkK+BV4LkevN
rt4/P6Ih7d5j8Y2/lIOFyTgYOg7y/RGZHvbMeXPpCDN/dd8elGNZNx4WtFlECwgI
rJ168uDYMuATvtKyYlfZEhbZnCKQ1r26QYYB3NnR9POFge+Vno8QM2pTARl0CRmJ
yDYU9dBFhqsSP4iSjzgPx9Z8zuR5XD5r8FfNcVwaGmtxSFwcbIU1uwUJIF9erSJy
rYwr0ffNqnXhEs0BoNjSOWBpDFdGfCwUpYkU20sKjYxteLpLKrlOnhiWAUfTo7mC
PRVwR/pjJ8xUabX+WA7yz/+Exo0ZmEEMDPwryuptKdzSdRVMn2oWPky28AqZ0bON
GWou1NDod6/ubOywAEtMkwF+3k5WiOfHMgB7aP+q0NSJ0EWXhgxVGHtm3J9HaREL
QSYCOfEkin+C6aTCs1XMFLQJj0sMwTjFkb/yDlrdpGbR7FeEj44a9/EmN4QsrirT
ZRSd5EYsLfDet92AvfHhFcrXDArMHMYf8Fosukb0bD827ulgzaoOZGZHF8COsQmi
LIxqAD86ZydHmu17oNiabYVl2EG3IAOtxSNrtNNHvFO+xrPnjoIjXWdVyMEu/Y7K
qXQaD8cPhgcfF73Hg/uj2fMqMp+/FQV6n5gtONAJ+9KL/n3zyALZfDhJ3KEnHD00
ETTfKbPDyK1nMuEbOvBYcY/19irP6CPKR+kP0sMBIVwgRO+a/MD90NmLmkgaBfvv
HUM2luIlTAurFXzXsyFCVEwroXi8W2okw7Hptu5WVMW6L0R7C1vaJDtQ+IPGL54r
DbWpWZhN015dRULZiSNP/HCT8tBLspseVtcO2j+ksoF6gEgWIpGaP2Hr9Ka7DgGq
BcSOaP/0iCK00CRCVUxUwm+cpTuVHhGhmfrPPcIPh4Smzf3+aJ6R2u++pOItfz0U
iQM5IqkjFa2UiLQJVM+QEdkr+7Hs7+SDoh6gotfYDz8mM/wI4HKu1QSow9mC7OaS
Ma2DkviLKDZ83G2A+JlO6AJdXmcHOv4kFsyQhi9AyfeKl2kR63sE55OTb9QRcE+x
cKDeodt1nyflcvgqzlPz+FY07CYP2zJBj3b3x8VpPVG9fM3t7BUjja/eDwkzBGcA
R7BDwh9y9kJpJ2m3fz6xW94awtfm0SWUBhQqZszN8Hq/ZnfoPLWByWJQ6u6nrX6Q
HM426rBQdlLIaQBZ/qR9A0sk1JHzuW1lDAhT4KtB8H4YH3UHIkm9FPGTHdid9mRy
KzqfxLe+pq/AGOmA6ya6oltpi118SPr1O3kzlA2HhudmVblHihDdSlarcRKee6xq
7qYjosStWHvBzDQYvBFVIishsi91QTOaWeXs30emWQn2lGVe3qEpDIF7uZRjsnu/
un2uOgOVzZRVobZ6yCWLJOun7cU49bo5RXDpE/NtBIeMENOUeqmE06KDv3d3Nanf
sJQ3dA9IhlxfdPHWhM5Z8OYm2fVTlCdDAGEFGoTGdHRYaq6IbmLNIHNA+hbwJBD/
pQtIN/FM8nTDs+nFR+s1zN9LCHJsqwrIsPt5yF8ilH7tov2lN3mQL/lcVzyxiEbm
hN4URKJrQrpmJesRvIae/+9Q4HoKbx5Au5R9Ea82e4BZJIm9dAYQyzc0UWVT/a/t
h2ftpmTMszf0tGveNKB/KzggOJXWawe+kT9IS38UAv+Ca+zgftm1AiOpjQu/qXlv
lXuyK8zmHWPKUdVSEKPPTpBlWKvJGTyxSZgtLSWOY9x2T2tIwoTvsAZE1UXOG4cC
uBakm5Wl+1ZqhBFu7HLZn6UP0rb4Yvkry9lJpCEnZzmKM2YK2tIdQrY+RP/lXy4V
PB4iwWBSvoz8xK9jhrCNM9KfyRf4J1SzXicjvtDj8oHikAIdDYO6GjCveAZY+daN
w4HfFx0/T0iNOibTZjqQC+9sy28D1hF0dssaiG1gYik1MrILC6qDdVbPUjqsI8Zn
El3mlGs361rdD0uVJGZaPD3blGDwe41TBNsHW5QohCamZ6kCm54uy1mEISmSayrx
g/gTM6SdgNulh/w80QcDW6FQ20IYtvhVioGcRtduhoQUSzgnI3JUBLVRmZXHOZbX
25EZLSnzYCWjZHIh19oMYWmKNFDUq6a0TAvnUhLMU93tB/Gh6LG7/QWkwBMW+/d7
ND9GexjQ1CPSRy8C49juYDhlFRkdzJam5AQk01+61YLpisWE7ensPLdSf/lwat73
UotqOeg2hjw+40VI/jn03iBmw34FxCiw/1nXKdwc4OA0ThtVCRHg3vlyeuDlkSId
lQ+sE7zLgE+KQDGxvBJYAOagHQzdlf7oM1uREpDMFqBA9RjKyx+Q3o5QKb1TMMrg
pJ28ybysO8Kuwmts76KTMS8AEyDhc9M/uq886KitdmyjhH6NZa0KMM+K9fn+H8Q6
SriKoxVEiy6R8GKbWSRIjnXvDDk+WBZzouLYW2c8RosYYp/s+5ThBaWaZOqdgjnp
Wnhoi6drDGtTVibxhjAqWL6l0Ws/MuFkVGRwm66YwJhePAfj+prqXeuFbbqbnkws
IoUCeLpYgivWoClYYQVwHtITq3zUyLf+hmFBEcZRx9UVIjxT7MqpgMo0Gsgcshq7
QGXwk4YFZUE+31gWhUBBNjXeucwi7OHXzSNlKaXZ1QZNtwHHd1LDdVjWMraIKF4t
8ipa4DUOWlOIaCauc+9SEPHnp574GTdXKT54kXpufHLwcqDLc6Nzr4oseFvHGPpz
tsz7I099IV5Ze10BeJLSESdRComcAn1jKSmBDgvSLLWpO/A/eD7k+zdonGTqo0go
fEEQdIijP+oRtC2hwjqRPJ//imBvyDG0SSepgSin6fbiBBAixpib3mDANHIKw3fm
zSaLp/FXBv35JB/laym+faspF4IBFZUpasUouunON1koJehUqMz2IE2cLfW6GxeT
p3/w6Qn+NReDC6AdbA0rNaBkRAsdpv8xEkkOAt06thqAMaNj/xMY8c+y44eCuvyu
UwPht2P+1cBC5KffZwVPIwsLrhdObYF8b0Iu0qkTblrQFshSTvUfzDKxqSRA9RfE
lFLAgz1UO8IPIQ8i0AFVp0D6EMZkYmp/4sBAh3EzR8QFr0U+ERSp8o/W3hSZ4m/K
lJyZuiVZt7F8PqZDz6nOOvxlCJUZsJ1oJDKPcyeIYpkg4LQhwVLNQwlD0PG0VcUA
u8XNvAvJxqtlxYws+O91DBJ1H4gg+4mcdTzLHiJQw7HO5hJkbFUh4WPJZKBjpQNF
BqEJ57len+Pp+b6YCo3db5JnFfaMuHZGpK9SlssyKrmZROHoyzjeFIwS9iCx8r4q
fBGGtE99M1GPI29Ir/EYMXdhjtljSstJ+wj37rK8hMIjvi6VlPPPwaZ/u2S29+/F
LP+jXMg16ZWycjYpiXZHIK4gRNaBpoc/WjG6oEBcAz6ZOso/YTDxUtSfZgWs0b3m
ASJ2JytnWeWTMBKh9ekWbmXfk5epGwfwH0UtY5Ca2BJAnG40CbTZEhFddZkHSJGU
MGeF4jLMJEZpZ21zfOJl3qVl3BUqiqJkBzJ2bxmXng8vNil/VzndPrgXGVp7ymj2
QEUgMYCp2I0MBYSQ9zaZaRXDKjFM8o4xGdR370EjLj/otC6hKhXLDEFTrf7joTp7
WlYf9J7HrvwERu49t6qROlpkAX6VaLg1ybABbEldrTVgxcwQoMFilJF6oZAaSGSv
ejBGxTRYlCJGcX49W4eAkrNoVonHWVpVa5ovAXDHbPuVUUKuOjPKCLRPKlFO1fQB
VovymfGDsD+Dye/m2y+UcRgGLGrBMhLDTnGSCH4O6Ucs0hdiG2goS9wwDA/uCIFL
HlTuaOQcXaBHTSih7ccl6tZ8Wi4TP+lUCdEWHvvo0HfP1KyvzlIPiMHLDvEt9T7a
MPqldyjtLJSKw0Jz45aB2Ea9F6wYVmAI6OeW/nG/xMtrushDkMr2n93MLZ2ueO6K
lUw2/BC4xCDlya10ST08xqjmEb5/Q49XdtTSkyjDF6LGuxkg8s81OSBM/y/EpGH7
vVGmYz3n1lutT6URoebXMGMu8mmZpJ8R0sZQ8drX4iWEXeDol1h6T+3Dc4iQ79N1
c/KiuLJztTVZjGKlve2D6MsxbaJxWnGPKnlHQUv23rDZbGBOnGaFLjofeqZ3ANBr
TkyremuOvQmZam7VcNXpJDInMnw7gzNCdeHEBcY9jOOD2gsqYPHbA9gKyov3GK3B
56Hb24zWg0fTtG4FQHhZZlKmsZxw8AZ4HZJSIqvwwztoySY4eIYCHQFZCeL04Osk
/WMOvKknvICqorghOEkgWtMLGhe2ojmh6BksNPvTYreZyObfqJbIH+6xSdyjiBvd
k4cn3S3iMVXqvS0csp7HlCXjVdKUmxhzp8x5Jm87DpU0/gJ4nhq5MfxYIhFJhrd1
Dob5Vp0Vj94qKVFjkDDLEHlPxTEzjQOCzfPu26YsZoUQyx5GoRoySqolFzb4gHJ5
RTBc5d8NoLLIPgNGY94MhyDt2+5VHOUMyDV+lWAwfNWCz7tM7baXF2y6A3HK4eYj
tNufbGzgHDxrceysXg7WfmTbKDCVeG3OYWiMxE7Go6QbuiHfvPrSHFMI1ETIbezB
X+R6Vv9WUbovB5LUyQN6FpyLdIwW/GH+PZG2Mi11EhlLZNln8kCAXTktAv2G/anp
vLd8v5tXmu9WdhMITf1y1NXNohq9IL0XDw9swXmD4M7kuegehPAhSwRw/qu0ZI78
XocdMEHHxTPpvmVKeslqOXh0jYQ7D6PRV/7/c2ch+qCcgJ5AADz4N4bfgC94187r
m8T32LzCsb/FexLI83EObwKxeYgBvWPzYPmgFZc1lnjvLRA8/IIROrGGGoINU52t
lv8Pg40mj9aWFEVF/Jk4x5/qbBeE7urERuS2XU7j+6GIdjzEP1mDu4G62tqXyOE9
JTu6MSX+q77q8tt+nP6Cm1S9MPxkMKLsxmJ9dmg9TAI6mGDdWN2OZQDTLyeej7ag
uFgd2RGjHiZ+bpaH1ZVMMm/7n9Ye/tj8fyRxRf6uTITuwSrbojZ2Q/7jWrSMBFd1
XOQqSCkQ6u4ilJRm8VdTcmzUTznJIwCNgG+SX1zC6G+NPbbDJ+3CtKgjOE7unkeX
YmXj3KTww3nX9OF/+pTjhQVGJs2SepTF3igrY1EaU0DrRXHQSHzJO6W+uquKs61c
s5Wej/Y1u09jCdUX/9+a6Qt5vplsr5SW0hwECVqd4GqVGkNqfRa2oCDIEM+sSTh0
VqvaUqX7YXDXW+S0d+76gQhgxxxaflNtuyVt9YJB8n2C0srrAmUFVl7lp3OsyaYI
G4Ly4khpz3CdqBFkE2eKiuzLs4tFs80kttBQ8U+rPW4t7G4+QOHsAO5AmD2GVe+m
dp3s97oRsEnJ2pMWwezvevdiZKmmjPFvz2ihouvnttPyX7b/MAGa01p4UUhBFD3W
1q1tyiTK/vjA/sOO1IJatxDVYRYAnwmxoIpnBpalFRFvjZzi9SeJ4dF8thcKMUAr
eAhu75n1ll9ceoaNMhl+osQ2YWGJ8lGM7BpRcMOAK6DQhKCiRSQ8A9Yn0j3uhz8m
N0ty1BDckSfXtJao3gushc0ki0JQSj/cFP4EmxtFnFJRJyKlHzGNQzImxNprQbOe
rNg2PCH3Lghqb9Qsm/eOKhyETw8lSJU4h9fqSIAQaDMh97fsJqAYYC/SNsXl5FIu
sPBz6s5uDdstS9O8eSoILtsMlVjEx47TVOXVq4wRxn+I/ahY8YKYHqxpAbUW3o9w
X0w1q43IsLaEgK62RRmxs2iv1lrt+kjesfPCWp576QNhwvLrerJleRYnHdzLXaiw
mLRJAdxPhUSBLZSj2jRq47RD5v2rbbmmjS1rSbKhNEzthKaRbyy6LLgrNqoprHbU
V2Z0zkn2GNrKqfTIQC1XaubuNmldqN9HJ57wW9PeJHRjA9FTJAforwP2hbtNjhOw
4EJuDXmuFbTPhMjBYAFI2UAb/chdx/58+PgJlMphuiKvNrOjlnnNVi+dKMgfrkU+
I+fV5VngWwTI9Myc8KWEuyMxnihjhBRf2wxMuhhGLlHq34IpQFsMrMx5Km07v1uA
cHrr4wo2MzLtdCtkmqIpU6WLa/43zAWoWuJLLhU2A8mDhGxjB27YQ/Ach8/YsqvN
GQad+A82H9zUsY86NARxs10bouU7RDk/wAhInv+n8RzjtdcQD4h4mOAwPO8R0+uC
BA+5n+qjyyIOzkjZHXvc5GTmp+1YVVyNSjTZeKXTTjbBiWEBXDOr4tSqvZPZKJXa
isxRRQoJHvH7Hx9ylP5GxcKlGcQ8cIXIWTT946w7d6GbzWVP73FRWuupFmodfAyK
5rKsf6Xl6f30s5zcMmavEIglCeB1lNcS0nw/IJcdfqcHk2ktGxzFfoNSxRB/1wa7
gU7NfWwxZclz8bs0hqHO97zt32YGQVNQEX8c/94LrqNF0acHP1U0OGT2rUvJGgug
r8kwSrjFavo/vEBhSwaXeyfalLgBMWMlapnqowVHjoYWIVsYXW9qUaYsFC/5kFCE
i0kzjNnyh/rC7zjT+qDjEa66QXkTyLzuP6ULRJUcExUsqGNRa7/obMgaIWN6rPYg
Rqa820JKCjWXUHrKnawDyl4wO/5MWcCOyzmce33M97p0iYr04rNS7Yn4vjx9LTMX
7lEzdUrQPxGtVj/x3+0ylxqTBfIxxhFn15HB65ZjwScvj3VuqECPFtPPBcsJEjWO
jrzib0igV8ScozaG+e1YaTFGLm5aJefpkA5CsAaXRGLisk57BfnWFtnC46eUkxFR
hYvC3r0Omax5iI5jg5ZvXirjbddZ/NShi4l4uPzdfhW/Vi+TChLgEryoCBFKIa/M
EtvwYvdGXx/AxRQyzwBvNE3og4nQcBnYlmVx/1JrsjOYnllFApGP/vUMGdb4poFm
jCg2RsBrASC+zgEbDCfgfv4bZuy/6bWmDHvwgcgis8L2Tj5k6u6N23CaWqQHQ6J2
w+CHRjpwuzunPdu/idUBeVpE2bxB8UnrCqpz+kUucULsODmWqUFMnbDF7zEFWQfV
ZPIp349whfldanBn8UzBmSh5Rtao1PgPYiJIS9tomEJeCNxbiNKJbtdXlpwj2MrD
Roi/FItj7gvCznbuPkQzWuTOOcnjO4oz6wsq/EDl/QnbS4mCjbs9tu+NkBEAyyui
U67aFAfgIaXcjhbIfGcYCT2Wfpd7M6CsSybiRnvUgybpvpV5Z8K4Bcif5QTdS44u
FYBz20sJ0ISnKgOca734bZzchXmWBhbrWgznABLYIDOiVnfjKgQPn69Nn4zTqo1t
xzl7pznoKxrLhQBfM0trwNU+knlZqfYt/QyEzsjFyOsTFz18BGPmx13fMXqo8xTY
4W8F7IDLH0fl4ZOeiwj+LKSLwpXTTNBqwDaZB9nuTMz/xj6Nn3w6O3iaqxm3kClo
h2Al06awoKugTJaX6kltfj60pFpx+1Z4azPkpUkL/xLA6IKHncRqOSVMyqtOkf8F
a6v7gi7ISx0nWOVP56yXnI4XMj5HubBvgNuHQtkWx5UxPLNH9TGNmPoQ4fx78wa+
C1KmGPrnzV31P8k+htbumbjetVOi1eFoiPoubKlPKT/h7TFSC51TR3Ykc080Hf2V
ZQukoQcNQRu+xk57B3tXRfItd+AW+erOoGX1PdnZEEF7by8TOS3E7qxs4H+xb8zu
bdf+/ClsTMD0AMa3YD8UPplR9/S+Dy+WW3y1nyTO2HONjecu+yHblko/F75V4pNS
YdIOv/MXcgd7uWNeXlZc7UXGA3Lc14K/pmqzd1UAwfss26M16xrnvWAR/mAK5Tt6
ZEdYMpAKh+7JQNHCnhGpdjyoQv0Ouh8RP/DjFwIboxPgm4JSwCsArUzrqnUwCmRq
HWDp5GCnZ+WFSpyRl4IY2B9wZWyX5Tve5Wi5+sDlHstAOUiTqOW5DThtFbqlsnFN
iKY1g0EflKCtcwmHH6BovlaBPGpGftn0t7X/hZX6Zkg4gnUuG+vE5qrWZemHCAFx
+9HaDPXC0d3S312zi1RRUoKEqZg5NwxcH2NZzpk9yoUPxIx+JaPKaYQLMKEweGKw
n87cT0VGftgd6fBnftBfXkwa7u9e/+ArLhSZJzotydVD8/tucLv0OD9zq9gK2wpJ
IqSOVeJEqQVYvW/5gm0DNl2oRvqKR4ZCOTKazI6DRK0mRft9ln/5bo/yvKON159a
tUzjUlWV6eKN4vNF3tbRyQAZrnYUtW+opoSaO1fcffG2nRie3/0qQ74x96fI014v
hXnQrsMCkJ7/+cr7R54G/kPpDs4RB2MN/iCkNrgDMdwhlFfPaoZZ8g0l9KqEun4C
EGBoBTbRfu/3e4tm86jdBQ68C5eqd+ZlNEStDVIntkiZghKlfZ7vTmJm9RC4ZHEk
DjiDjA0c4bKWAKl/3QB2/ki9BBl5XZE5ImGC116tVxaxDcFRulNZTrnPidLCt4XI
MIu2vsBskklsOFW5W0b3rmvSCsX5H5yxt2xAHbOdyCkxHKe7RSYSUugGKOkVpmPh
I2wj3xcev/RaJUgRzZutB08JjRIu7pjeY+3jR0xi0xT8m1/blZmm2BytfNrMs2+N
Y2M42v7b6ecfZHM4LNJR7H/Dwvq+AMnHYZN1uNc76SVSIrf74yrdqFZLSTuOOdmG
5NYrWSnGUyQTLzTxTuyY9JcVsqr0CH2+upiIxkWzWraZRDteMYJM11CI3PC6eIL/
/xs6ud7e59ncHayhPuBGd3o31317xvp9CjWhTXvsPr5CdD6cFeqJgi/IsvVVjy6P
XIV9NTOCn50hGcpkrVAgca9ZLJWB2ZR83q33/X8UVo4vY+wONVl0zcSyQVwtompZ
nKEbaxv5SvuyyjI1j4vex6Knle+5936DkVZPpvrKA+h3gjUUxzkhUL0zFzULAyWX
/rYHKCiST4cGGFnicV3PP1IQhK8rry6Q6RYGuIYcVhHjJwQ89av5SNillpf2rjDe
NRXbyD3FlcWCovrr0fupUqK3YzfmghKGJpoNPQJEKcWTdABD9LSLdgMVSdUOgAjY
vnPm8u/Y3q+NuZtMi9tMVdtXLT5MDZBxy+ep9QiStMTdLO9Xt/ecdnQpFY5/hYuh
DpP0TxBjoo5h5zJBjPGFoDFU8oDi8nBmpz9TwmDwrFiO3U5VFFLV469XXRRsFhii
1cnQ7BljovEzLHXd74XZ58p9EY86cfxo1L05IpyKWaw0827bQ/r9NpnjVjg6BvLc
Kd4GIrwQbnsAMEe7SEfBJjVIleAmbmGekbjzeaNKdu86DkQApTWiVPc1P5Ub3b3A
gY0d7LMsX0WjnDo+Vcm3XMuQ4rtmxTaEabMBQb3XO5cF5aZEtHPjN0g70YLhE48w
i3MNlZzoqRAmike1Q2u7AiU/yAxTXsUUFWI2bB1OkV2+EVvDDzpfIqAqfRyos2x3
L2YhFb+cWwI3wOR92Zimt23nNky4yLoBckLhb9xKJ0/gqV0KoAT3aaezoPbyi3Hm
u000Kw71WneUQ3nnFpA7s3iXeKc4GdFBj6RLMpHwPX4beM7WIKh7EL2gjg4cAQo4
LXIbYAUPF/Fx1sVHcWbITeWjGWIEbH2g9kGN6N+7ziKHF6pLLu540jMl7IYuQ/WJ
MzV3Utco4RFlFG7zjKDlpGE24GTDnKzF3WGe0iDOAwwYtQLmQh1BQX0RL66yugBT
XSzUjCGm71eaHP35/PwRBZBKXGOkK6k/I1CXs10XbBBYEWcsKICA4CoXpF58Qvix
4Z73GH+Yy/ZO4JSR5yrHGhuBZAzHWTfUdHLQ3dXOTqw2sTuO2EILhyHaLRMv0xLZ
F0syG6piGqvD5iVsBqrc8TjvSBMw2JmCJR7vBwBktiMpcZlW5ayLITATQrNIc8pv
r7/Ij56U6/ghJoRA5ubufXh35lMst9YN00Fuo60YWs48/yN1pLPnjMOXrURSOaLk
N0kfJyiYLLgdLfmyl1GQVrMdymLbUe7T31xMkeEX2DV/IQcN1FQXJDFEsp103/FS
mn6U2MvEQ9tcOOC5UHJA5oSNSXoceSGy4vlabK6OxhtkmaWt6qrRjKQW3VInFtOB
0/QBHxh6fSuT7GtD8eXrU46e3MXR55p2GiIMVj387dq+Uy+FzdGOpdD2wOX/YM5G
Hop+VCHtCs5PuXm8fZLf0Ex4Hc5Y0IkDVZFe1xxXi01dsKIXm0qXPZW4CfRhxKIW
24OoT+PAV+xn8f8LdlFHYSn7PnuMB7HXy6PnwGUCZkrZR+YQIMbHG3xLJlyajgKg
smu0hAtuMT5T8snHkYqOXenh2POXPT1XSzHkFNqtD/yZYIDNiPIVJz0lkEHTfgjB
x2S4fvqMTaW536rLOguvd+Iw65Sw72vwo1oeRjg1k/lzwwb2gYrxXhQeg+rk3Htn
IK0/SCH2EN2d96efdIOmcJAMR99NjmMupxvW+vr55NsjKg8ndsaMX/KSSr3Z0Qca
8M4z1SgDtx68b+Sjktv6ZXwPXMea5L+H0iuxjocVFBxp9f7XEgWCgRm/upgl6GH6
0oNYqTLIoIV2rohHeyv6vO5ib91ioZgeXsNynfDIc2+jYwHQBekRxauk4iIyA/9r
IgaHUH7IRc73kxZS01rLmZfIrQylGC0fNeH1VCH0myGejvd8ttPCptl9SjiEii8U
U/A+vhZgybNmAzYuAmXGL9ssgrD7lY3ROXYOrm/fcjkl3wbhzYeQO/t3GIoA4Xfr
SWapoqqMIQMz/Ti9JeP6VNFNbHWpBEirB7qHU+Gkviqw52jDaa1/Gd7RcSVUSnSv
TweL/jACpR27qonEWWFZfrHh0G59fER0MshvUqJi5M4SOS/x6Gahchk2V2as7yeN
Eclbj0RfzkB7Kd9D0Fe498A3HQm+n3VZ5OZvx172NZvUbftWAjD5lLOr88gftsUj
F7PSGADOmmIr5Y/CWav0PlGi5MxDKCO6UBR4DO9odm/llFayLfUx2k4DhmGGXz9l
OosjNF2U/JyzLaOIK2Km5GT4PCrbKxKmFK8SkYaLLh1LF9D1ZSWgdNRTJZL2pzRo
qOzMLu/7G6OuyoFHva9KH66w835haOIRylgPrVLaR8WwgTwcwL48E3Vefig63AvZ
aPiTmJr+VPeDoswGXKE6dAgok0eE3BWudP6HvGKpUfKNsY94U6q0yeR8lWL3g0ly
OgqQRPVxwahvQcap3Iif73i38A0Ett1izvQNg9GeoQXdC9wMeBCJEIG1NfUTS4mo
Z8XxXTeklQc6VqLll+GJ8c1fFmfOVRkFvcgB3dulWm6eK31W7h8wkfBIzS2BOUnM
wq+gFmCcuU8yHwLGMsh3YIKpoNdmRcDP7gecZ3tP1Jz4zdl0Hx7Uy0Cfd4UUxqP3
qP+mQVSZGZ4OLO1EQ4pLjrAI0kDP0go34YFbsUuz9OXGpXQ7r+6jldMU6+X/Lc+R
58hdtRGNd51dsGSCKWa1i6rW7b+Txub8PcJlpDkCxoxQMgYsLGyp+plQjgMWYZpJ
qF1pala9pSUzvVLZjzfKTO1xWxIm1NmAx7rnsrVHg2PCc3c2Vq9BQMKWRBG7DTc7
xT1cTJWUm3gBI6Mf5gn/ZJ3P3j/30lvF8Zvyw37FSTwGQJFzQZCGE6Z8zNc4yBxZ
Ze9InClUhy4Wf4cM/lKtIW70IpIrLW7Tapqsh5p6YG8zaBDgIPSz5g4TT+4y+1pf
yrl/GJO0pi7EeIfQP6lGYC7QPuK49WhXv8sUHbmLeYbND5UIfgqxNmg6jUUyg2io
BOqFUP2udNzw0HnTHYOPMiixEjxcL98dr6x612LrXwbXJ72k3sryIt0dkovVRbb1
toPrSqs0P6O5/eZUIJTaG8w3l+zY4Qw7jEIrbYEnXi8jvHk0OwUG3UwamgucO+bj
W/eRs9gNsfDWQbSoagCptHnu5KRw+exyExOLmi6cFE0YB0iOzLp06xsi7PTZPe8w
GpXvN4S6hbAY3awXvam6voa/UmRzH1XyMF8Izb8O4gQjToam/2M+rmcbIU2ofkWA
rUt8zD+UdcSr5llyy3GZYnDqRHw6KxVkuXDTqQP8jg/4PBIOTX8nHwb2uj7P3zeV
6QVKygKu5ZvQjRv0eByMsKOQmMzswRMB16kIR0VBSJLvLMC+g8NWzUBfQ5carysD
YgWI5ONNlDKUHsXR5yd/9bOwnXMXnc12xBKhLxkAJqZ9me5BKDWmKrYmQHyg3kxT
AJgIjnXSvCs7Tv5FeeAc9DwmZZXDKlSGzZ1RDV3HGbS5ETXIcTfB1pM+jS7Sh62V
FU+/pTBjDcKqtTHvwjLtx5LheQNOuGfxOiz6iKv4xZyXb7p/K/PZa+NNNHdTP4x9
JSCypjcY2nFaTytqJ5uV7895pobOLmGsHEvJlB9xgVtfd9/nRLuSt3W+2swKjzKt
O6QWCsdCLBVCBeS/3h0k1obWAjySmbKZV3PMmrCuT2eEy/oo48MXxNHadAyhtZzU
O9RB1L5wNObcRHUaC21s0KT/6AlanmnZnDW14H0sK5ChbC/2X4CGdxjr8UIJGBhY
Jir9Wpwqo3+EEdWgyj0moD7TosBFKjnu4TE63b4LJQ8TfuRsvXlULO6fjXWR2mxS
lXz9Ya4/3CDb4YQ6hd5SbqhK8qI/UIaT0GVeRLymiZNJgeOLwP5Ce7tlrxnqVAVm
yZPw7TrwSSdwxHMVUUtXkP1KnxqJuukj/IbYg0PhO0aYK+hKWORoIlRKYG36Woge
/SDZNjVarnl+ZQM3ZyvJ7TMiOnGLxBzr0TeScVSywyLd7hR2LCFkEYOWf+m1gYJA
w3tdOpq/JVTvzVCQHrMj2t3E3JU6GBUWQCeKzuVrk0iwHgkGfGGXqywm5YAVQlAv
qUhVAIAEW0iIo2zs92queU4Hapci470ZqSMoatIn0rjZsUchHEqUBoYPOajgHNcr
Fa1ArYur1KhCpm7jlYcwPdyA+H8P8MmuJKtKhVL9MQfnsUf8Mif/sicQNu+R4CoY
npNQ3Jlw8VWtVLcELg3Nos/+t9+s1NKrZh9zZAlDGCgYV+8FV1D+4L+xfajP/Hdh
S+5zeUWRPJ+W+3uUkuesjUrIt7/9glrUpyXMCZMLxMBYtQc7+hPi1JVk4u0N7nOv
vYaiCoWtWpZJR/Hjvzv4pcumSTH0dDhAlg7OvoX5zvbCah5DK1+ltcwgxV+EjajN
5oN1WWg5GLmVEhAkbNlpUj0fNLFTaOV8L1t7cdEH1iVmIE/vGIFYd1UT1Gq1im7P
vM03ertc/gxX/vL1dT0kV0FpcKu+kGJwezIKLgja8A2Ey82N260K9hxuDdQVJLfe
tO9zwJtTmwxKHDLgN3tEekprL8/VFqvX23GWSDnErP6lpBrMbSDph5coSbcuEaRt
RKi8/c2UguOdERCG6FtxdSPy0IOpMVYtBkcV/td3H1ThWte2x0+q90MyD8qvym8a
dr3DDU7TPCxWnbJrjnPLHsI2YrAZYbb8WJqU5iIjxkq/6PMJkfyffBjlPf0ROdHF
mOokFFB3OtHgyRNWL5EY6rUADurQjz/ELOtwbyUE78MLF5i/WWuPOU2DwqSqWExA
FeouZMJW4P8MYpLr8iAxcW54EGdMYbF1vEona4wsyQa09ODkog1VVMkUlPrt0a4/
pnnUHafAES6/BV+c2F0p4EegitB0SNeLNmsVCNpAm9ucdFtL+zq/M6K/xpnq3xsL
YkLEjY3c4RfJpoO/5RtyjxLSev+pC7u0USRZ0eFxaCq1TBOp38YNhP6fscYaKVd5
uuXwO6/JG3Hn7Dx9ObaOmfEIBfCuPQ0V3mzuimEC1qLhxicZMBtIFqg7cKSsOdiL
K2qkz+S2YEePEMYo2KSkGbfJwDc2nGG5ryxflrArsHC+gHlEnpZs+qb1NCDen1tk
5ESZPqELhIQpLnFUffs6PEweA4iZusPp+6LsM/UqVSqa0EWM7iam8jiiHYLWP62I
kbQT/0Vbk5cNdC6yOOhXwFUhn5tDOGi11cW2hlL14VV64lP0CzmQ6vG+3FZ++p6l
uF7DNxTE6nAXdVdNxaDFHb6h2b14dV9S9TaVPotckhdJnkHYPB+In/hEdd9Fp+5G
BL9caH2nH3sIKyilve+TvRwEg/zJCFX00tMOMNpmED0SpkGjB83gsQHNdoHilrez
Zj+vLjF9B/meQ/DTnB3QXB8d4L1btGukAHqb6XTMjwQFxoSz4m79ZvPdEdBo8AU4
E4r1jqboICgBbgNgpylpDyg4XOzdHHlx4Bft/JTp9t09ZPNXMX46oMdM2XedgyUV
yszTwvMSzMMuw8gV+jzQQsYWdiKyhMiOsNdaQNIlEHGjnTJP4pj1A/+1aMRekT+/
ZqNooDphPwQTV0nwyFXJbnHD6zXGcWfoOiAf/6uyAM5XHemVxF2IPd/YlGKrDAEL
XTXpTNTDArj7Wd347ScBjC+JxpqcKpOAZGDVWeE2Te0xkuYbOmaWX9ulRPSuPAxd
VfS4alGZfl5LqMW/yqLTNUYChsvS5f6toGbs2RZun0OeoIDQfqiwp1U7avqpBzGz
TUmr7qT3vzMmHZaU6TFOMnP4vyOV47Msx8E1zzciOgAW9rzA3JVpGyXzqZbYOkCL
jsjm01EaQJEy9gJ6YnCUEEoIFqH4NYivyOhbXFqQHGq8fmb7y7FVdVcVuPWyCSN0
Kv7hDB1W0o1gpcUFayuy2fm7aJzsGWfyuvYnvEAEo9K4V0E56uQegCzONgWljuvg
lDWresrkhBZVWwXPx3eVosrwz/6Zsefay5GTaJAlGHtS6yj+QoKsLcuWfkTEmtg6
nW0vqdl/ze7A+ESy0UBY3vnRnDmVZQJB/eG+5JRB/fzcUmePhayAj05nRZ6+PLAR
tHLXisBEnzEo3bDNHsKP5HsI8opu/nO82sDgKOV0lUcCC7SIJW5nvQvwRLlqBIC+
8EBTXZWappB7OKHLXex4Px7VX9scx0agVMkRopY5a8cHaQNzoBQrkdYsUZEdbtPp
GbTtoJsZVcb2ZaHbWBNtpCdgsQ0y+S0cDd9WzrEtb5Vc4/tHaA+Tizu5EN0aQPC/
D+eBTSggDJujgwluBNgI2e3FXt3lkAM2Os/jHEJLZ+bvlSrTF450OIE0Oxit+lc/
4xnvnQt0ooQIE2/u06loaiPxz5oeoK9faFSrhuWFekpFZKc0o02ycQwIpytZ/TmL
JvZaqtrvYDAmsRimGhK1tM3NwKcE/ileMxhoBXcV0AakFTts+QB5t5sbrreb80+N
O0MRaPsGc69RNAlVQ9yUj+mdmPhcTgxQyOi03zcfzc8HoDpD5m6+BoiUyItLe3nA
uQ5q1+UZrckSX7Jqsy1jjXjGaCACuFORgYYwbruahCLyTRgjVZ6Lr8tNnu+dicYA
h0BkAiYEMMUWancGYR06nPugfuCBv8g/P10aBZKx5z6/HqEVfprcCb3IBGJ59Q0g
9qpmjHB2YDwXevBty0hq2RMNNA9hHWJds9tfiJopP/kbhvGWTLm0zA5US0KoQW0P
aEGuRebjJ4Kb0j7fEUOseuE9SHjqqeVTRMwJabscV5yn4YY67fhM0Q+yxIMmEiv+
aXvJhxLiDDUnW3+4GQZdf4lO6625FEX1GtDkJ4FYiIWuL5BlbaS0ZZKzE+25r6Va
+knX3kBI5b7sE2vYXboRoF72JThjfpoZaF61CsTTH+lrTwXTRPEPgjbAhaAVjYw6
4wEctHE6TbQ2f+WroWXgy5NeVOSCS30Qhk0ePQBAWXvVi8rSqhgh4pJw2+rpSzP0
2Mos3jkz/bZ0k+OxYsjC+xkf6iW1M3vdZ2A50+xF7uoi8WtoOukiJzy/hsbm1Ehz
a8CFx0w9anh2LGQNDplN473U29inxLbuUZ14EGyx0zg9PNc9hEWUrWwJdiEMPhPp
RELhQ/5Svs/rR+7cgCCOV4jbcrmM5z0Sxr/UqKIeoRzNkeRQKTukcx9U/nC1Qps0
fCEiBpoNnepdqtyRyqDwsqb6KecCdwmpAF79/qN+WrfFxvqn/xiPuPfBRMOpq/4u
syVxkCOsEHbxyxe/lLZXImj17JPfpBi04hlpPSJrg8zzUt3q7DrAySulcGTYPPuG
WtlkDvG3HSDKyawdJVoboAgyLHfFESNZRL3K54Q+j3FYwLjzubf4vcOFkvs3xaGv
NSLVPugDpt0PERCpZWZjf3wVKdDtfPMhP9LAiY26VmDMc0+h2x+FMTVd5ggpXBgK
q69m6bOFX1uXbdGkRJIq5ZI/rU/eqnklNlhhUpf19wnQmVutQ08S4ZYXgITVLFoK
yLC6fSbocYUrSWpW+B+4D+q7n23o9swsU9JvP8jsXRQXuZx19q5VRSHxQ1b9PopM
AIUsycZgvTfyJ2KTo+CBdNTEO0iak7mgmk5RmrvuDJsyApOEVKoVswzKpcnxvJzD
1m4rA1wcDxfOqMYYl2uyYejE/ffFoM69ZNynpY9SmabeF5ABpP1zYgtLSccoqIgR
3QiqjalGc5z8SGYeSebnfBZG8RYyCjDzMIx2w50BPvRocs3S80fYUnSTgp4PaqQO
NpCYZbmcfR/HAfXNBn8akCyflSY/Egry6JxZmKmP8AE/YlCr+/EItG67R6G+cQoR
ZUJqLsxhN6LYX/uCtQWivtbdEjzHYcZnRtjXM1pkR+cEZEUVeUdxx+oTui9c9+G3
xxFmak+YNBzQbDGXnpkp4W4sVir15OQ5Zt6XjunvFa6ArPBujRF92HqBLddai1M9
zJDv4X90bzLc9wkwXJFmueIqGIjXwtvXhsvNGmUVWvVS5iYQuLvDHVjyscGFJZwX
WzkBcZMRSGQqh3ytrO7mgT1cLuEmJ4xn7DDUTZykvKoqjdj/dmrhXcEc5MLhVL5B
u6hHVg8kbM2KWRqBDL903T6QgYzKsDl/SJWAEOOowOyd/+aHAPoCcupmLZK9NGDi
Xc9NXE16ogoqVnT438yCL0gTWkUf6/ERQ1qXODsbjODKoaic1pNugCGowbXIZ3f4
QHoI+zikuqABaaXv4s6vWfmDbGTecMPiX0IOhrhY2IrhTLIl5Xhc3qHEz7gWC2d0
SysIxyaIi+OswHPzVPfH0iiPDYNR6fSgLDFmEDGKpwhbfmGGq0XT3lOIfLj8NoRF
F+reHBGUSwDYI9ZssBDJH8FO85QX48jzzgubPuuAfoX20EH4cmluXcn/k8Ts2YyX
j7qKCOw6p+1TGQFN2KM+6zM01JthiFNVmiQWzua80VVu6TPuDpUSV6eAV85PVGm0
MJ/fK5blYQ7CyusqDUYDL4mHnDjssGdcEu9m8f/SIYa3QWnuoEeyJffAQ/Ymf+Z7
MWJczSRwimR7nJXwn8a43nHrT5ysg72ptvVPxx7ulE++wAhcj+xgdey+HB+DZ2P4
IEBoQrAomh1OTHWRwb2cH4KqR34gFopSdnP9vI8CnRVqjUCnhkXZePCSRwKPhI+h
PLtZUrYrWOlYUH1I+9mCDVFHNpbx8NnZ5/U+lo/IfYWRm2PPkCk2D7zDA4NQOPsX
Fx3EvZED3J+Vllphm3wBBKymgd6xQJlnDqArlABrW/nsPaMx0P3EaG+xOmy8tltv
0+lHGEKOd8eJTpolt0Kd2w2HVTKZJ7DTMhoXh7QHBucvfG9js3162rgnnWyhDpmM
K0TgqY9tn3FdV4dgFEV58/nN4BIOfIxSIDUVVrI3FWYW2t7zk0LFL9FyEcG3i4v7
v9fg0lgxtsxf8ZP5tXX2iULTLupuwbOCyg6k7zi4vedtfCn8D8h0+lxMTsgL5uz5
iucFD2tmlnUK8Wh2kypcGMc8H4jAixUW7Cx6I2/+xyog28hFwFDt97ID+Enec8Cb
L8/ngnQ861/f7w2/36x/2Rj8f3ZHDF6c5jCamEGtN5qmYCY3wt3/Ff9omZCIUZJP
0W9WngZzav1IVVEZbKx0vtaoPkhJ6lfBPLC7eBEDcrGyMKip3/ZQTZRsODWux6a2
yrakxpTBPQTnyD7IxSFm0vrq2TATEUTy+goI85JxH+MJGjPq/awZyHf7wOw8H59F
omzxzDWLNDad06jERDlI/dNBIeXq4KrRjl+79oWtMh292+/CFst37NWYEzAdy2Sk
9FQBjNyAAvyWtcYeI0zSiLbWK2x/6tGH8daZTKv7H53M6826ba6B6XnSm+ECnQOp
Em51mn973hCQdKDIVL7ySlWInhQSs/NMGnlZtnfoT/p45cE/716V+p3gZ3jaZM+m
htqWwyLghOULYIRHtoqTCvvd6cm3TX7g8GAu0wM04sAYkTohTXu0DCNsTQxiGyot
vA/u7zgvZDjS/+zDBZ+DGF0RhCZqSFpQ0/RD+8dajhFawaeXUVY6oh2eUufP011X
zTiaUOp4e5I6D63jboesZzEy9SlrhVNe3sEqeZrI7U6F9GGcPZJogkcMvsoh6+AC
g0OxvzTjK41eiM1yf2d28rpj63Z5GzyV27QE8iU1FkVl0UjxVCg5q7v5Z6xCLY2h
6thrjFGHKQEVkhTEPxTp7dhDmpI4XMvD6p1db8apYsc7BkMIhemulqjah2GdorzT
DuHPNkvDY+UQmIWyH6EXN8Wq4/CMxFOr4fhqP9jK9bfDjlyWe+XMgkzj0S3evpFy
gU0I/LXAxIUWSyr4Hbm+HaEsH1Pu5I0OaLvSrXDPNBNNWQwxvHQgegthCANnBtYz
lxcfxwzdHTZVtiplzP92WgkF+2nW40GUzaP5BqKKQNaWrMhhd2SdxizNp5wR3gO2
uB7FvQBq1kXiPbIiSLPwiSorL1iPjq7/5EYMOTfqM4t1697L28Oo65kf5kuvap/h
m86MhPDA4rBROVwvmWsqU5fAljj8WbzbN3UIAIvE4VQC85xLIwvCIdtvPx6iPKy4
5VZGbNuAvEpxLcrbKubXRbbCFvg7Fo3BsnLyHYKvBe4u57m8HN3/qo4VTNzCy0pF
BANCNpF2pwcfsM14kZJe4n5gWyV9p2tHZyyDeDGmF6iPxSGuIe8jXeX9qU2o59Dv
9oeij7z3l3ww36usAkkZsAdTCFAGiNcpLzVB0Wcf9Ef9qpNxxubScoOMDxKeM9BW
BelqLARxgY1xRDDGT4/PPxDmNyV2x0OFMnMqAD9hR4mfU6y6UYC5VP6/RiJHS4xF
kB6WfOz7V6ocrqbQdvZDeM3qRZQIVl2D6HABAtK+guikB893vxdnreFm7bOWKcy/
QTfvGR1zOfkvwt+z9adKhVAj5rPNRUrTmz1H5/8hyV1ncteNSq5TaOxRn10BEpV7
jBMezeXLvegChXrpmbbqllL4vN+JX/R8XhLW/LlQ1BOh3/Sx7CDwgqgQlAtrDGMh
7R+O+ZtHuzkSs29UeXrV0pEWW9pU/f5xb0iDVFwXv+F5p2lTMHfpvoV0oX8OV4gB
wIThTjnp+8CCcr90gnbTnDgDhoUNOsaH/YZliLhDtYpPMOQH6oskBwQNon+aV4Wn
CNcRihjqwedxB+0I/PXLeNuqIwIMXHeaneGfxllREosPAmnhqftaiHtsmZ9UBcaW
QCm3XHpSocARf7Sj+izNA8jXW1gIw5T89meTR6Xr5jl/0aA8ALWsbhfbmz3d+Kj4
hz+8fcbP9FdZ3XXgcC/8oQqJiVP2wvVPYOeZuYTtNZK+B8ggqR9RCgc3YfL0uWcT
kyhtKO13jy0xlIKla5m1U7aEsBy+XPfZbJYGA49Z/q3Kc6npGNhugDTtG/sRKWiN
wzZb1Gq0+2Hal0qpLeKdyUJoetuFubeSByubfREQWg42tlKiIvbBGhHEGi53wzCi
P9wKeBCFeIGH8mLg1zeADdCJHghRydLhPmvlnQ0lSwOjSBUkbSFpPUvKamYZQ3CN
YwPqKP6kcCz9Al70bJJNHobGc+wr4YPCAlsF8f2v1DYQDAQwAycI5JTibp4HmxG1
TYtIEf8YyyXbF4pVB+658F1/Daq24Yxu99rqLF9WbUCfVCNNPDiZCAVBZIb6MIXB
iFuf0UkrN0S4xcolZ9Yuj6kgjtY4pKJeZNewmw/EMT12mrNDFIkzj0dHfAxCv10M
3bdkLl4ChDdJkpOqxq2SNidxIY1O22qmU6q1F5FHfbXxh7MhVfskte3EIsCGbuDB
ujqdozx8A0D9QHa+M0bx+fOidduhFDw8k+6GeLF51DYMO9Umior1FbxCrTv1NUhW
OJCSy94RjSGVsFOyInF+NCr0yDcXkTmZq1amQKHEp0xjFVxI4Tb8vk1hQorB+Wlt
sjKxb4a/RFM55LuwPS3szf+cBgaFbQYaBdsjMqdjmY/IwL1ULv3Iryt9Jt590iFe
q1D+PP/C0cPW63ToCQDTI3IRTNzIYAbaQCOW/f1KmpIAagFgN6lehczY7qQ/7Ij9
BTnQDCYPTcgw5DK6CDvpOPsi7Rltco1E10Fw4cQcvzfpJd+IShYlIzIFKW87CgZc
N1jiKS3X8AWOBb3w7t0UT+9DJRYo8BrQR/b8w8IYrlm7uYsw+jn2HBNxF4XTCTIU
h+p7XfSOzyHbLa9A03f2IssD20bvA5cwWvl0Q8cvHokChwS+EGsO7XFddTYeOI8p
RItCYSxWRLOYTrIBzEhRUzCC1DAGRDqWIgc6C+jYvEYO2ZYdQ9GKoPCL2JhDWVSd
+KE43v1g4yyZ0dFMh6XeAgyoEYBDtxHH4zhE4LD6rBV0S9ffGHQsDkhSi5ej9KdC
5fR9J8/qmhvr4KOyGEgyz2KOyVYz5o/9AgnBOhI3Bxphin1sp1R9J8FQ5sO7Ia3W
qIUfbAFPZy85w8iIYTbNGM0o3mNtKxnXKclkj42h6cYd0unDJvEvM2dy8lP1nKAc
YY0pZt5HQZJae3r07TQSiZocRsnZtobDCBAoSzSa2U8tgmiltf1L60SHusGmSYxu
cc9ErEIwra3ZGgFwQH/nNiNdB1Gec3qwd/G33K4JTrxntEd7Er4As79HsP/Zfh9+
KSzga4rRx60osCyywe0TQLkV1B36oCzGRXz57WxshKfsYq53oTvNbBlOhwMoH+gB
OB/sgWSVFmyo1j5OcYVugqFON5EzfcuzH0rRjRnq3v/8eLk8y8X29L6Mlwd5i/LE
0daXk3KavRyhNrl+AfZkfQLyMX50hZ0JzzMlVktX2VVXiMK1x6TCkVSnDcbS3QDr
/HX4fK1lcBfFYAwYR4UDauX8FROLJI/xw+RQMt/I2ZcHJKxKatVOLKVi1BkZc9lF
X1vCanX+1iq0mafwdBvbPng3LIgE9sFwOslPkcbMjutnF1Jysy4gbteysNdOarEv
sWMRTudDpskWDdPJhOAhIUVlZlCYAtg0+r/xKNBG9NneGSctcGdmX2iTZ48wsOjs
ZO+2WIxKh08Zxxjk1voIQCHgyYLrpCX2yNcI6wG81MS2robMCnbjBNfbLlVxipK4
MojobceTomgy2RctCJSn2+nzlGa9LRd1c6UR7ohO0O+SCwASL3Ugduq9XOCmA3ML
vlksZvqa1k6VvXfyzSeMeH19wIL2mKX1Grz/wIv122m2eYpB6hF/xnzr82N4XqWa
y2qE1dcyywW3wRRHbVxh2ZTUFdzPbcZsyZqF0/2Ap7fzWrUGH6IdJ9skGqMinOqU
ExngDfDioIHt4pzNGBoC4QjKnZSrs07txciypAhksDDjqNpZT391vSD9Y2eN3EQR
OaTgbsx/80GjrzW0PYusxzu6zDCr5XGP0WmPONmBoefFtM3zvYywDytMSRPxLmLo
Gr2YMUq7rLLS3+Oj97713HuS3jO7PucFLxZW+vIj40eBO1BGz8wiWHJexMIor3qn
0qKi7dnzCCgCQVrW73CsfA9zRNo6cRdWXZkQLdmsVStH76eQnAaHhlouReGui4k9
c6DMcxPnTV0zA3543OaCw70Ehh9X1xRuy13VmT79W2vIld9Jvm11WeTqmSEemydz
yc/S4m478NQUOcCSVgH4Jon9bqVBonvQ/bZ2outiwMqfEG2JVqp8y72cGfzApoOB
LAnWBG1JyNmMlPP0gYsBNWYmMwBoHNPgJFEyDXeCJU4R/6clG3dtjlIV/mIfJqaU
ytusYtlUgP2nS1svWuligjCX+hf14RclsSPGAjIOzKt5iKBlwbBgiDalzObXwolA
ie28ye8aURZfHrgH/aytBW8lja9AqkEJZiRvW91O/MolAoasv3zwjPAOu7GSXyCw
hy0mICDu92iAaztivmF95bhKhL+ln0+jVor/zxLT1CHxtCdGoVr5R0G+/IQXvQjz
7HXZOSFk5zpeCqI/qpkrIEY/RrCrWyNhrxamWTjx76tuT5X2whxJIeSC0Won/BX7
ChRy6F+tHjuoRJoQFzvzIOsG5rTHgb0IpiB3HgWKqyENgYGk7Yrzml2Q9MQubFhq
rv8nOrBPBINzcvLm3Q+LAdaYOot0fiZnjlsAVdzmLujxZzXmE0a40RsCh3Aydh+b
ASrR8nohJi8HaALi0zJqtjhUHbSaKK49QKfDie429KMD/dArMhLPKBJgnEk0LXCd
EZt7g1589Bok+Sie6bb0aG9yKkw3eBUpFF5us4aO8YPZ0fqi5Ym2g/VQpomOP6zx
D5F0eL048bolY7DEOt5X5cMyHkw4KtxJBHvzJiko7p3q7I+9s/ngezJwMyaot5Gp
55C4HQmRHp5kBg+817KQFpoqkjG42oagYR3DG1ZQZB/E4kkUjnNgxNZxQv3I2lNX
UaCzwipRoAs7IsUfH2orXL/XABfL/F/86TtquIw3/GuzAx1Wy/SEIP1CkD+m6VLZ
g3uoMvkWKf4lIABRHVDw3PEOiVxghDQqeUmElq1ZwTRjMfI77cZ6BiOtT14v5K9H
ZfhrGUPuNrRX5K16u6/3LRl4WEVSdi7vDzQ2/Wpf4/TFxix+Tg4G5Nkc0IK6669G
Edu3vin1VMJj8099g+ucmuLYuZ1S8TgH7VtdpjyKdB0rNBynXCTFLm4HaZH6TEA8
RO0r6oikyBS+eA6whnFoTwOxkczwhCAukTeNiXHbFr0L0/tEi+z+Df16s7PNcMVM
a+3HNPap/Fn4Cm+fbr02W+7G1WtzytjX1VaEuTBxKRBXAe0389D/GavVv3pWnE0z
74ObQEF82WRMvmAjnfjERnkFEoNei1H97jC+YNBS59p35iMXN2YT52cfTDK8Z5Qr
fkCSDpCQOPSqCCj6aBNgbTjW7t2cE66Uycpb4WF9YuETjSziKeFndBlxV/1p1MuB
akfayBrDuzxazsgYHnZUZYedxcW2IujCRf6DHFE7Tm1w4jm6iUrpikxAHK9rZM3n
BLtoYgFm0SeQI85UIqXIZG/JdtsDtho3icEB5i3+Q64P4q0BzY1ee8z/aDKNy5Dr
Nr8w7hzGpDBs6V9WjTYwWOVlr+AdigDJvVKgPpqrYhSeKo3sYc0xWvFs8GXdmMXW
hONY7Loha1IR05LxDi+ue+FqVlKyCuYSD1raaCmdSlPu7/tdcyixrelCF0Xjrm9S
TXX5JaUDAABoKx6btubW7LvyrassyOARgYl3sHaDMWPI0/2JM2qPzYEL4DxTwR+D
ncPJwQQQsngJ83zJKMwJUYFFPcUhaooUTm4WTxxfIu8gQy15HVED95FeppkhyQNl
m9O705x1tOArvH4PEu/XDwNGxUe8YKkLCb7wlPqI9JCiuER16PJGsEevRlWOKt1l
VyI26upAhbCLPHDNXfwEt0Y8cYJ/13ofZC7AMAqqWHYJNcwuZYHLNStbvshJNNDG
kCA58w3w6vziYUCq7FrX8hHTJ/CVKc7tSDCo8N8Nat6ZAdvuhnj4BvLVWKSX89/S
FnTIiptEz5vKzAO9dX+WEio9ieQFmljzs0gbB+vwwCyPy+op9CppHJ250IDU1B8X
Ojn/lG1bEasks99Sald4ENRb5MtZRJ+YA/rNFvwqVs4T25SOIOJOp2AXLcegiByY
ZxAe40lgKixYxP9ouQ1NAEk2V3wm+UESvliHcWhWMIvAoOfK7x8l63e8vNE/uC4o
WeLatkb3uuqzEGCBRUOzYfWWMLUigfb3Ir29FjD54tw925uUi8KFLl8c9yz+S78/
VxouaCGpLXRe6ESjlfTGj1bi8oP/KgQzNSWm3DvPhn6k8qxSE4z7B+uFaTL2De/v
AVsKPNDJN+rHW19WuWCFWDU6FTxz/idBOjcUawW8FbLdTMTvGUZnDrkWRCcOncEt
qNGQBi4OWPb4S9L5UiE8O4SIfZXzPoA6+qyKkQimK1GqOMMgtTL51LC2sjDzpXI8
7d2U1KCIvwsvsrYSFZMLit/olGYhVJecnq6nqBxPda52EO6mKSodISMjwD1a60Ms
dIM/RJogtfy6BZ+IM4AT5Q+kMDRiEOfN5lqkIXDX+eGIC2tT64hJJJGOcgWHFZM+
jhyP4BlIRsUQDYQ1WOFyfTVkn6AThfWwEXYHyHaqHYyaVROIo4GpxA6g/lWWtgBT
pirAnnyuvOVidruCJzYwH6/kjtw051F+MZBOUAtRnI4QLU+TjJHTAEt0UZoZteNb
38ZG/SsJm+AF+Y6ZcHlewZOH5ZlrGwXzhVrYTBY68wxnHLyo+cjKmV7M7k7oT+OX
PlRqDbeZKkAAStcAb4t936glhs+mZbL7uNTJw1QOtmO1V8ktp1O6paHVeXScgK2s
K5V5UsreUynk5x3n6U533wie5+8KJYDUKq3LVWRll/wuKUscCV8yWtpJpdD6akHA
KVpSRzKyY7oqCHXyK5hiK7NUFI43WO8rRqbijRYJYwwyJbG8rJK0f7tp/aFIdue3
xwYSUJ1d/k6fNAcVr2PYU3fOl4SbLllYwGdbRHInQVEZ1VhzhAV9JbrjivvFqIoQ
q3apSYdhmrswOl6OpzB9mXsTlp6cw0lydxiJor9NAfcENRXsVxQV1JaMDFva2d1R
PVqSz06fY9VOqqCtaMwkHBF7V11tXjEfQNv8HRgRJF+MV9YGPfTuI8wwSqw+KHom
P5a2dfdf0kcGK3qZBUWnAK9ELYDdaeScl5gG0I0nhZeF2Y/VIlx2u5TzlTdLO2gB
TsxHhyubJy8oYpKqaz9or/CYG/z0S4iRIpjwMzLZV2v5GkpHthxr1X1cIDYyVSey
emiuwhW8f8Elhe0A/RTuhbMHSvjtK8P8w9s+AUMQxGaH+K6ks4EVnLx/e4wWT/hL
djG6Rvadl1zgBiaS6NnWlhsFBysdAaXFpAZ1Y6vXV3bb+dyPxI7PY3eBz7MEwkW0
TWVMhuW1krKyxxwFKSYWC/ZGNpFrMkPOXTJWznU6xHpyv5SgpAFg8GcTVb/r1Xg1
fRrXn7YnmYlNInB43DjH046yl0ckD8vyNWfSbcshBuqsBlJq0dsQE+tRZ7MwNT2Z
PyMiGOdDKyn9R/CLpXys+hPI4WTq71a2U/bAK2rduZzWVi6X/of1ROcop8OwBc7v
AUBOsXYCjeL9zYzwQ4tluL5kcIvXX5A1R8dSzWxR1ZFERkUMTH+u4+mQ5k2auT+4
HZGY+f1d/zd/4eUztfU1zy1Uj5D3feot4E/hWo/heEp1IHgn1ZjO8MAiS1puvdZ1
urPE6ZDHvdhCJZFTzYQplaUdhCBLtoIAV1Lbdm+tnNMtuiFC3XJgYvrKGCNtTB2A
bZm1GqFgadKcqqJDI/Qpe3A++ERyeI41eLEvRVWpW2Gsh+srh/sIBCXzwKQ7Vwdd
Eb21nWb0P+rcDM1tIheObnTeBa+9kP1AlpDz67gxSoUT/2t0+H79qeNC564zftr7
CjkWMeci7xPcAKN4olxIxH8sPSFLFGTfWc3ds3E5bci7cZm5wqrjlWQSHst2t0eH
MWh/LYta6q5Mu5q+YsxfEGkAFxSJhaBAruRh3uddKc1OOd6JqKbzpWRISU1r7CCl
/ymdGmSVQua6KpziRKS2psB1tQXILJmN4s8J9581UqaU+Qpvo2jDbfK61YehXLkS
ApaGbFdpzx+tqSgJJaXBk7h1C62xf5pzfhvh2MjXPII/AGuKBi5KMp60WSI5Kdx5
35vny6T9B2cb+xQ0hd8WTp/6DJkuuAYDplu90QuBOmZJi9bF36yTpBW02Q7KZez+
bauI9sBOj8DtpNTttty3rAfrBA5QKpgKosFD9OOYWbCb9zMpaS0UC40AvlDZBwwL
Z1gyNmyUhsAwWh1YRDILCBy3Zc6JYLWDr2lHFUhL3D/jNWX4kRqVamZiMiXZyYzk
+nvnKsvGotjPs73fXz19ytIb1vidamSs90BO9HJf+N19XmUR2jwxCl/SH0X84UOY
R6BQsx6TKNVe/Up/tq22unOydI3EMi8lrJP8sG/W7kgje25fJbh6hiVIet/NB+Bl
1u7FB0ypW6v8tOExHAudgFUGJLgv2lA+8rwBl9pNyfP4BoXTKnMPoPvo/Y4Z1eiR
XHA6WXSaNp9dHvVeNgjfG220vGkBEQ4kR3y0St/rPmDEP+zqznqT+K19MDEWPBZf
psuJHHpvTa/fjgWWBwZ7mHtvo7ivunUv9aY4quLraFvVOv8CgBYWBWtUYQCiqx9b
sOTWfKDpli0WGmxO1CttWUyvYaqzrKJ4szdfcMrdAn08DC6fFBp/oA8ocX5ykMHV
gCtmJ365GmMErJvoyYbjTFF5WhFyXMngBRTZhbzrzkhQOf+i2aQ6Ft3cXL+9QaFt
y7QBI4aXPgO0F0cFB+MFVGIQ8hY0CbVMnNt/qpvWvrW5+ayGrSYNkFPZlu/pSmY2
UujNb1KZAcQsl0aSWBNwRYupJeAj1Wzv6lX/iFH48oqSGzH5QQ08ZA3ZlmO4zJ/t
gsRzt7sQRdAD3YAatq888BAEF9ymplNwQsbBKgjGMcrTSdgDFhteZvNbHAKs9Ifg
P0rA6TalEph28wpGHZVCjHDjt+FGoYd8oEa1n0s7UkTHHqiallVebHxRJfU2No4N
ycvGmrvsYdBFhd1HB3v5XjpB0stttmpYtRFn0PkJS7TGteTbivklb7xW8H2QUDHm
qDYN7sr74eqH+evBIeaEeMBHTDyxDRoirQ4oXGVec+yP5E9PHVOU8/aaB9qtHi1R
0D/cV0RsCULNq6h+53VQkpFZg6eggOPqOlW4VLGdBvf7W/JuuqQsVcV86KPg6DGN
EwHCJPnqKR2bFPMRNFAPZrOo5Vw3aajrn+/qnqNHYOEws0h3e42mVb3sH0E07oes
fqz22dyKKAuClnJVnUjde+yAVTRBzDlkn5B/IkbkyV7lWc1NbHr1FqS6WVt15g5o
oMzkdBUuzUzvyAPUwAZ3EmDcVbu5cQMcAKa43tXi/Gn98w/TV1MNmD35HRB5GKcM
nTsdwacHDC4Cke5WL5eQyPxY0IYIT3zyVA1CQt+FOMdhGFFck3bQVBC7MQ9Y333p
9zEEpIvL5PNbiF5ZzWYSPewUV3AsUjZv/IlBo+yNbdPJjJyL0zOKd+QWuwIKHfNd
hdKDmTHeg3jAiXI17apq5wa8gvC76NkXRoDlQaFqCgfQnNnoEydCQH03xIEjVlCQ
Me1P4ry7WeMs7JiiOYDg5n18nXKbC+2upAdhycAKI+shfZ2wTpqvx3UAnFxGyBEm
oBhqeZn1+AmlqObCvf7QdVTdpApEHsmmAG0aBr0x3/GREK+PpJgRNtc38GP9DQV4
gwxBM956SIEHZzs8ws9X1F3YcoMMg68ErD2Lu4UKcG/Qiq1GvUEWYlfHBWMDVWSC
JE8oiJTD9tylVJGUDuI3RjqCmESEskzCX6t01w4ei47mnuKvxmOHvhaaNX4nAv/F
sJoSlKE4Qqltk4Kco78pcTql8l2V8Zo29YldTZ6poy0zFLvZcJTU5hUhRFynLNgZ
r9U1DRpz6sT8iwjV3Y4OHkc8k3KGeKAA//VUSAyRWAnYmrSWsJuZE09h1TLX1ETj
iyJlxdjEYPgJpoivtfNU4eSTBYji2slsBx+62USZ4bBqQ6GhBKW3MGyM6z+UxbB6
+ZelLUy5Wd2DjB5Ub3oM9x3fTu39f1vCzlt6jgZhFRAVq07pxZcm4re/Yfx6QYFU
2OfPa5cqvB6QFuv22yJ4luQUxOxO5PSguGG+XwPBlE5Q4cZZI6ORVyx/pO+2PbqX
EeFjpdHLyE3Os0kfVtZlK13lAhBfFZuMiMeVK4GaT/GFt5frDc8kz0+J6sVAi9n4
LzK7suCVni49h0BhyQPOyxPl++WMKzeuOZ2LdhzMgaw/jfSla7MIFQ6enRb28ObH
+ubu7GrBfrJNzcgshdwAf1tnoklPpScjzOBlDIbMZBzNqCJOchTiq8p6VV9GekWB
lZHSmiRIwCN88BV2yqh0F9eKpCKhjLzG69IXi15osS24gCPJjmTbGuUnR9xW+FaX
tJGYIhn5Nqqqh35pLDHXOynOeg6n9ydRkADKC8AYh5PZSJyGzknjvN6vTarrtRli
SrzdytBthVS+Z4Pgfqkg0U6vk1WvCzl+xxXnhq9SZPa4/tzGmyh3c/Qnit2pjUI5
xtQl8LkKQleeWi17ZB9oV9vazipBNJzAYFFamB/1smgyy4oGK7O6i5kW4g6pX+RH
OrBRIOqnBU4FqtQf0q8RxUq4Dt0Fdp19UuH3LOgvqE5PV7m3aPSckSMAIGNKAt8d
h8MVYjlQ1Y6sdTeus9i7DlFy0XuFYQ08+XI5dDjrOf4ZtEV89lIkm+/B7Ntio4JQ
uNL3F7MYhm8qcV3H0NNEYNsGUlh4sXDR+aT0sb16XeVbJI70F5EzUPQ20aeY9Lle
WOhj17gPR5cW5byIRw4hKOX5lzhZetS0CMoe1TY4XZOkMQODAkWy/rIlMG/EpN7y
FRg0lmPVixgfTU99zqqaJiFtZNLw6y0MjSHKkpXpQ2cHyClGWZ2STiU9ZqxXL1DC
gAr0VCmoTNAiHdXPkFkjYDXghD8HUofnQTGn0dCzWCgt3essQu66RUnHZsyaOx8r
zhK8du8mnYPyzWX1Gk8i5x7wOf1l7/nQWlo4NndsEpNMtRAIrnjwkfHKgT/Ac9wc
CY3ooVpWOXqcN5fNy4t74Nce88+ZKtz6Exl8piwg8wYK8svwSWYMmIIrFIw+yO68
S2JOU9Yf8Dz5VLt3hh5+VjAaM5ner6gHMDivPzxWhfEBlwWSZmrwSd1sSZ2usdg4
A49F6uZxInHLGFF+kryjOrUDLOHR6mMGFuYv0/bmTe2G23O15VHyDWn2DK6enlnc
OTpdSrokUqI6bgr+l0eYnKxNbCxZ6IlAb3dIDTlVoAxrDmCqOvvPIcTU4RIkdLx4
8L1jzAxv/8syhmB/WRNH5GmKd8YlEuCxD8l8zB/B9KyGHj+X4JLoh4Wr+BJUksTL
txVX4m2KsJykz8UBkpIktMUImfJ/O6DO8SysbSRigo2dbQtEX9qWocM+U6vNNn6+
mS9HfVCqJugCFFcrtFnu5Z/1uN4Cz+5lhdXna4FVOFv5xPU6jPb7yBnN77+54vNR
IIh5OsYj6rLM2qTWtTCX9TairjoscSSD+PadTZ3GfZ+G27I76T4FGNzcsjX+euDn
hPLPJpvgfq9uLWc5AT8gakPTJGl74jNwODfs1IqCT6zBgvewg+JFqq0We1HD5EES
BKdghvfz+h8ch5rikVG0aOQkchESjTcMq80G7NEDHNDsim4ulkFgfq0fJxOuDCr+
yFTDsyCYhjTVRE385vU/pATnrY5XzWKeqj94GN5XQurUlGzZqGXFIywHly3bkCIo
IaHsfuhwOvXY9yfNH22lfraPDHR4SohbrL606qUjLPTrv1fqaiUc6sKJi76Yrh9d
D3NbkIs1972xSPQQ7XHlz0F3QsisO97a+WOeeuuYxgyzVK5ecBoyZ3sOzzUKUrcp
FjrrY7HT8BfHm7WMmnNbwLgI9yVXzogemtdnrFJkA1grwIKmqGAXbKFw2ef82fJH
XADQ+6chJtTIP3Rxj/3zFZZx0GiUgX4zUEA1DS0oHWFG8JJH7+eRozAyEcJnaqiY
qUmzqnTYt4sFnNNq5EflnRfbOO1qrJkCXmoS6XS7t92tV9WjVZfl2dVcdgzvAIKl
b9q5WLoag8/Rg14ckBn6RT0iBESNYgyywg3YBZNgvV5pJmX0lvhIMp91R8vT6U/H
EbMBM25U0p+sTzWX/QMRggWUKGLwK/xKuVIjUkyOyk4pYNJnxkJPpsNww6QvJV4n
PwT2WLllxfYs3ibOTYXIURtDWjN/6iWOtUujqPyIRmj8Ev8sBpdbuIL9crxbYjcl
7ocy/kFQ0/vQ+QzLPnv9ry/XLgZ56HrhPVudFLvg2tRsTz4YdkxruZ5tLYU9wg89
zvL4hrrRxK/o9p5MH9pc7vtPlg4MaOOr+H/qmF7Bz9n1jmlynlk9Dq66LEtFpIgL
hjhAJHT+F5c9Wj00Q27/JuGPnDXcPeUP8KCCpoLEebB2aoYxyEyy7ZHXms6A/NLK
JAh/VjAo4/5L2rf7DSVqlxt5RprlULbXT9PNHKywLT8bv8q37K+f7CXNk3qYusoz
9sL8/al4bWqzN910w8nM9gUtwIh2NmRGLVutMfWUdNUEi/VeENSWBq38b1KH0Gt4
ZdtKd7n4lruzKahnahkEB1XqxtQyrAGBMsmTcmZBVN9UQFKX0M0Kr3LbqisDRTWr
DtCXXmaYbVB7ZqmQUc4RYwJVBO4s4saGMILe3rN7Oqfi2WhxnR9zWGsR1d4EYUtf
9QLVEuM+K8nII+qJRp89H8dzjaFzBmY7ckoZuSv2ksicMBPfvbO0zB4L4+uBKlb4
4+YhUfTCfg1KM+1dlJmoqPjQPsaRX53cZG5V2CT0l9vljMAQMbY4HWE3A928XlQn
UooIqD7bFok8dMBUYzkgSPQQ4awbjz1JcagpPfkyo9tlrEGw8ZNPhGIC7ZBKQMVY
4xc2+K9E9Fq9lXUZz0TrwsC4RpihutoJO11v03sqJxn410KYFq5iEMLTfB9bTOy8
Vmzn+W/iSymNHq3djZtI7ef8+w7wllbjGMdAkVa7Iu19iQJFrXR78i7D9g1oqO2t
48i0A34G8+NgmbPRAobZ7/RcuedfdfOoX3mDIMD8Dix1lKGb7gxiGEXJz3eqj0Dp
slR8JDgNGTyrv+jRzfFHfMPHYl27h48fdNX6+erqv1ciK6tQDME//ee+wlNN6BAD
DzIsa6BldjfnNbVLxNwcH2ZTVHF8TANeE6i0FAs5Kves0PPHwtsXEYVjigHB1s3n
UBJk3HyBWoNt8h29RD3gcrxSsNnQJBMRFwXCGpyEd7GYdeDXNnr4HPuQDv7K2ipZ
z7YzzRaovzKG8oNXXsX6QYpfnaaea7bFwA9850fPKGSN6oERnYstuzbtgpPzK4/0
jKybT2jrDeTDsfWeNwRwQkFTSU2VNLw3D38uM66lglO4WIV3GpJobMoGxXEd8fWi
eN5Lv0ltwyJOhCLNB2wFEcURk/YnzTpF3dQmJvDrplzpVwn3/+whYZ428DwUN+vB
bFXIaWNyc+5/ist7u95jpw9t1hTQnvRmE690HFxd2QLxuQNrEawKbUWdpVpxEQ2a
R7RfNchoE8dtKEFgIqVY6VkCkEes6cKjkNg2aYh/g/wvshs34ggK+ZZCaKuQUOJE
RyuySMW9IMKW0CP1cxKE1FsM9bLON3LxqVY30YOXEFSn2rycTR3BKrzxwrVQ5vZ6
0Qwr6hlxBYpyfH5JNFssyovVlB4QQGb0oeBtH9oK+AYaRmkAxG+e6GYeJyl1XDaB
rjy2x9tiL9urhZhoUSRqB8SALjaUbd/UawnJ9i5tnaMhELVTtDSL/ogJYB3iFFg7
T9yaWFsylg0aKSe6UsOEnzzKmZcjfzKLsXh3gDNJhTsF1Ped4AFHc49qRSB2f9Ro
XotCRVc1YDsUp9KhmbcC6N4j3Pr5RL91nwgx3pJehWgdwnSdFnyQG+rP7cXJ1lyK
yYD7BiA/LQJyf+eaa5GjVONuMJ0V8G6voxUMExCcSesx2VJu6MXtOxmr5gIYbpfw
HY6qNQC+DJ6Kp9sN2CxxE7NrjD6Iif/0DEWoOnVT5BG4sFav/UEO/4/r95cqjdKu
nd0lE2Q08bWxYVeiatmjhn+2Ts/8w+NVQ1/izTfXfgwhyZmvpBZbQSCdWz1wtf7+
8uzKbArA+Wfry9c6vW51zSicASedwnz1tJT6f2fmUbv38I2POLxClpGVTxTsTSEd
K4L6GX6nnUQdD+62h9+U0GZH8v3CGwmk9kzQL89ESMVpLqb/nYiGEKlj0rK7syYA
bioxdlzHt4cKZdOMpk5bgMNbtYzu0KdJ9NW36b3pbtjc31rvY1VNik0BSivhdYWR
HJC0PzQYpDJLvH7QHwOfhS1q+AjazQQa2Ik7oMQZssjogmRQAKA5mXMbZxKF3dBU
h3T8HkrveEMKPu+/zoBWM4gub0veb8mF8E1JiBVzd9klC7+0th8hlWZos0o4thzM
j4sN1tu7uzdvIEDYY3hGtoiIWG2h3v7RI/UO9Re3rW0zbMHMGy/vsEkC5xlf7UbP
CT4X2IcYNousQU+IYS2+w1s8ojlyezQionwOFyKgv++dp3V/Z8pJsmW2jonSh8hd
f8ZkkWWjrzJG3jv0Y1TSZVoFWdGAVggG44kc2tI65JPuWEcKHyXJZyptjbPG0qty
DQjTs9pPJDQzq6h+OqEVA8KmQsQLBhIT4DKlfrDeb86XOXzrRuWfN3kkz04IBWQ2
Non6J+weZjQRKBOSYv9iCERDHBagmLU5VbAL/SFOsOs1wcozyIC2MLdJr3Q47hUY
awSij9OzdJHTS9zpcZRAAMzEYOoeIxviYbU5XR82S7CIePrFkrS9EDQQzKYovDDr
HmcGf9OUtxgzTkwix9VrllVPw4p3ULfIxzvyagXSRNOblgxb9duiHzoFFvZaKtlX
RP7+D9Bw2GzI3PWdNSpCVIIoBCjK3nAI21qssc+36LzCktMKjuIClGMCYRIN+/KV
WSgmGXJE8ehPi892RfqRfOjIiBRwIrnmkqy4QgIvLX5hozp4H9mzVr/UeIWZScU0
InMsIvm5ANZ1ijoNaS7OLsziV6RXLWSfmvbRmD/KhwycBYT4qGchkxJkH/Kn2s3G
/b39lvfg0AEcRzwjy7IsLYztHoZsKVz/xYbqKmGgcgouFlN6WD9SDFb065ab59jp
IHCHkscyAeVn5lg98lIYGZ5MD/xL1YTAkARJyCe/3o7fA4ts6QIT0D8rh4Z5XayS
cLTPFJtypqBA33OmRceBDvq4I5EtSWjjSrlG9vp3dqZwWiyPPiUolMwdmkuhEuDi
bSjywwY6jLTasMtySm1dGoWj/pLrgjPL6TRMq1xqqwcF8GLHnMXCe0AOJwmr89xm
1d6MNBbM9l3CpZy4ojwhDhxk7sbyAphs92SG2V6H0xWNSFykbh0YYa7pc2UhM/Mw
+eOIRkg5p1ogY+mVWaqikrsLBsaYM4u5Nj+OBMkR3WbFSKqWT7yHj3WvWFCnDwY8
ggHQu6yBGn09V29NaY4FEuA3OoJ1tQZFFkGXB3bqFqwqMmTIw6xTUo54h5biaXOR
uY8EaxEYBA6Pp35Ac/3S0alsnioI8/1gMoHjw542DM2tcTHsGirPFXkJBqTesF5x
P2me4Ps76uSmXsaAiPQ9KWZsT0/t+Iwx2ZNoIB4FFjQpXQdpBSDnnLRHCljAbvVM
EDuhiCjjDhIOol3/Qu/6SZH1SCtxF9f4GkhgN+AXVIi+Mj3EDkbQo5fsaPaBpxRF
8kbZGQMvsBJ0sstYanXBMqU5lG8EF8yBl1eI9ONb0esrTSzpw4TXgAXz/Hhk7GHE
Rnx7CHBmz8MNEEdIl8g9eNkcnjSrAuvlZNVk3H1aDUracI+Yw6duj6CPwtB2CSdI
EInfjHjGqO8DocLq4hSpFOhYthT1FqeE9GOdBoBcoYlRg27nvZTuXL3cN82LY1Dg
Sa2vaHWUau1dIiliTuouED/ks+F4altZKrhLu/erIGTYwETQDxwrVJSgVjHySY6G
cV0WukWW+HIe6PrHfGewcT1SHGCj/hpxX2JmHFdRU49O71HnhTmFKuxCfI4Xfi0R
GrcsFyvp669Kn4+2gIPR/5Dmi2H4oMwFErv+pgCprCSUeH/a57CFCpyzfK9/eMpt
XXn5SC4qTDcG39TV5SiDD2gq9hKKA8RSaa0TCIxnAk5D0B9RUfOakNj1owTf5gVD
/PRzBVtjnBmDV3htvV6bjfLCJfIyXeMknQRq0OjOPS+3a//bcCyOjSE+kE7MBHdo
KEAhvLQLO5b40BI+HE9AEaljJ/yTcWdyASnMccnaeTpjHAJaBrmYbWMaSW19xIvw
sxGkBslwkRTjut4IP5VnXuJRvMlumERAP/UatvuvLUqk15ufXmGTRI6Z/KLuCUYE
+c9qRGoMEWfgR4gbuqMcPzdwDEX1AMQeMgFgy5iNChH3eCc/T3qFuI38Ltz3lSv3
5POSt+iaICDxbEkbFvZHfqMvBevWzNBOvAWjdSiRzLazxHb90Zo4zbsKk+7fYv7Q
V2FG4VO4lHtUi9ASRJfBDZJCssPENn9UKdzgRmZLqsrqVfQEzaFoRbulcIT2TOvv
iUX42C1ATDdpFELErpHCMj49th9sBlo4EuDTBXaVdVdVNdG4GZzoRoxfhegi8xIX
ojvtABs4LOL0axwutiWFCi3YUc9NeAaJSeznJpLI2nEMvRNYeNraX4qXks1+dqwp
l491uRNL1kCf0hTDavbRjoMavkuNSlNICN79gG+VaDjUU7WEZh+OPv+wdqPuwe/2
lRMvqVqaGgF+OVF66ra8SatCFmzVapHh7qfTvitTtdGdmMTZf7Rim10DOiEscyPg
Cy6tnK6BDTAmkSkysJUt91n56YFmT/piyxMUocmHKEdOlSdy0qDsnIqdIgisUSHq
PWFQL9/WycOMY/0z3XdRiWtKMIFWDQyoZsN1qy7q0GN0UsZYGYY/6PQnoQOvFdtT
EwzqtPZcnMyH/do7/zasuPtFPxgKl1oN1LcjRAgXeU2v1Se0pkeuGprmeSXxCfJW
51NXsblPk/Ju5LSvtK3zTI93RX/tXL/6zbp5++IIdV4pKntO7nhD49EpZTrITlsi
VWCjMRO2kWTJVmy6SYCJleizdzV3eQdLgxx1wDce5y0kIbOztVxwn19IEITrnPxS
E6wDqGFFTVxI3bY7Qs1qRCsW8DVpKe78GrOgWhOTQ68zNQQKjxPZvpZEUDFDZfXW
HL8SXVvuCAbE1r+7IgWZZsR9WCM6p6IT+STVDQUlP1tmXdSdk/MkFVkxghWH6WcU
V6kS4xqaiCIAky14N+/y8zcV/o+jRGO9i5od/nYD6Z/mjGXjGJ/p2YPEta4IH7Hy
QHqjqs+/pqMH/JS0ZR7EgVRGAKNF55BClpc7VbXIOyeBRbnzu6lcpVNfU0DE9dfg
GoQq4zZnW+MP8SyHEUcq3V5/rF77yOKTXqb2CqPkMVpGbVRpfb3xsMzzP4AkbHD8
S3LqL7NZxjNFUptoDYxvyQ9PXieXujZ1zwmN69/YXi66rirVVJrmbPVlHQp8wHuy
pI6JphYFYA9eRdwPm6MLT3VfJ4PuudSeJI9SN9sY/xipqW5X4UQX02TgtA9VYFyg
MkRWMjVEZ6voWzYtj762nrMs+ufVYlSxj8egE0P696ZhQKVB+USWoGq3IArN2KRl
sbKA1ltuu5WLFL9GfJWfUrR2EAmoe181klLxnSemsPlaMeke5/l69XD6N67dwG5+
pADIZzY/RaS9PwnouzjUDXvrPfr3FJgZK3a2wvMBoP60IU/AQ/upqG+J+dkpitDS
oS1UHYkTLtnG7LYFMRB/L/L4fyxnKCSWk/OzIz2LyCfmDOcao7nd/RADvy7VHoeL
60rA53mlmkdge4v6r22LrZAfzdn4oW+iEgUoL5S2Dh5WsbwkcjPOrabqAOoiea1G
bIYRJAU8BJS/5IXj61GAyaJDttnd+JRZb12F4vzrHAlv9LfvHDaj9yjyztw7tL+L
Oa2587o1IfEFxWLUw0u7R1AkQvShVycNNsm1c/zmUP8rV/lxj5Rl4Dk8trMccI9Z
Xg+vkG6kHIqxwFH5u95C4LOVw53CcWGIy+O+wG5BylEJ0XdPs70mcLCpozyD2smQ
cggaQ2t7lvpuicsvpJrcK2nuZHo6yTw5S/G3I9oQ2joC9P3jC+gc44BKa59xyqA+
huDni6ELdeg0D+TV2DxIgeFAeA2iqGKvdaw0wYSPQNmvcf5eDlsI8wcSZC/iQ2X4
oPMcqQJ6XvW70dWV5fbEies2Acyyw836vheTQ1da/LectM/hIq/ai6W4MgnbXtq1
LLXayBQ2IhIB7NgB1RqRXHsWHslb6Zqw5P1Z9PDYrXmQufgtw/TuP+d+u1M9SIzA
MJsEOelO2BpR2GuxyMjnFQuVDHFUEVkUzKH42gprPPXCPBjs2BsvBA2fvxBLmnnt
Czr1DpStaT7WTbiXMw3fq7A3qiQ/p6pDHgaLiBP3h4JMC5COBmhGufwFbDB9f1DC
JR/+atwZW/8cdwtGL1zJTxjaAq5iwjzBQztjYOI3BxG7iiB/SlJQAIoQhtKROSu1
8/3qplKG3jGpxzzOM3nDYATitDSpyr2+kwUeKrj/37ER2ACCw1FOsFU6m4P60Zc0
TTJD1NudclKRYTnh2nKVyUjABA2uQEAoskqq8N9w401gne2kRaqSu7hAXhb7vs3a
MxW6kaZdWZEErADzgPuv/kzPm9PKoHJin0CSj/5VvSCCFgAWvi5kZJys0wRHxbZe
7V5vrR9ZcJ1tilYMUwMTAjDRyxMQnIIddXl3S/9xMK9+UFDj3oaMX/hqA2krTj8k
Mcc6bpsK7LhJ/lvafLEpAmCLmg8GaU8Z4Z8W25siAbDBXlGoG7tlMV3YEl6kF12t
QXCTx/CDDpFrWsP/MuDTOJhw81gPNMOfYzqnVuccvwscVbeBLRvPyHZn9Lm+IU2J
YrsxL+V47i8w6pCXouG4NS6X0Sa37MCAyY/A9KcPMfMgfBd2x+1cwGCvCl1jz7G2
eyQZW3fvgsUy+BYYH+KGJqmwyc4GrPY8kQ/FXKHDJhJodxJLCN3uDhjjlziOCGFT
a2IzaTU4V2OIhhedtCJUNqfl22EI0HWTTusjpGMisf2iZRsyHeaFi/yKBBfe/SwY
aL1vcfKrtJAo7jIZeH17GwWJ5O7cYrG6nQKJ32ZtrI7PLkKzF4pDNi+Ze+TCJZkT
CfH5J0KDHXHJ/iCkkDmrQcP8U/G/OusvaN5Wm4Vc/gbDjnY498CScZh2nuXHrDGY
+aFJHotGZNNHQaTBtcJkbPkd0SmW8SKT+I+v6xBFlEfxeQ1JFiQzAK3i5ajN2sP2
AJhxPR4o1FUkKCDX+71AVhobySoXq/1L8yt5hPdF7t4qUsIkKtZrx0yUBlxEa4BH
zrmRN6ylMddDnfq5kKsEk91p8pe4JPEAsxctICEEoT5b6QZw/mIgKPO0lRoixUXz
NWBxbzLDmJZM+LT/tUG8fLFbLaATwyrethC1bk6N9AQhQO9VSNT3WOf+ghCgH2MI
HfOoU2+hpqEkfiHYSJBR0eLKsuw1MWG8Sj5WiYhJdewTymCy0jVqDGFPXKvLwUNR
tDtg2dNjzqG1QTxS8DMjJDTBL5AQnR4EVcRWfDeqI81P/IjkVEjBOZlC1JQF1E0I
swEPsrN/mMgmwQkEKxa3+nxTrpInuBrQs9XNgy/6OuITB/uMeQS506WWlZIQTVzU
pWEOSPziKVzVqeRivwEmqV6svNwYlDJIRU95wTrSwqHcRPIzf0iWyQg6h2phR+ZM
kpaxnSkG9uAgrJw4DtnqajZcJEoEVy4rjDxpENBSfpiM63mtdzum6NcDNm6Kv+km
GjkvWz+CJca7UtVKxhWR2ZITXEHPXY06ssH8APDdpa1gZ8WFGfvLjkcns1wFJToE
R7OWOvzSVapzjpB6yjxBP3gK16e+VmYoz9/AtMWK2ZB2ncZa3J0dhMzqliNEpQAk
Nn7HzPDc4D2cp/ihL1PfRTlUWAu1u6P+YxVPaB+H6VqGjnX3ttbCVfLaFocdVhoK
yRsAZlqBDVEG4yPESt6zfm+EZdR/oEOgmi3Jv4r/pPu1XJQtHZdNMQri+yRxu2a5
IkrjtI/vaAjllm1y82sO/HT4cesh83wMdc6kzTTQadLqfWhVNuSx6nFF+QwBUynt
Lerb7pDGxQN8+FYvxKVqdNeE7nmJ9ofB6ZohULrm9HHhJ12B8zjz6nvecphm4shg
lQ/Uw0csWruQCRUjApgufsZMNcUpCy8louGf9qXj89dlpBGuGZb9XXgyF0lb8fgX
EjWzGAyH0ydz2QexPsQXGFWrrazVZNfNtTzl4VBVXyZ/v+T8GGgxnRK1N1Vxn4Cn
uGdjd9VzXF9kidx50rWf/5V5z8UoXhvfaM9YHTz4GpeFmUbb44B0JG7CjdsbkqUR
LaFHNffalMXNKXiCD6dISe9oElpOX4yBNnc1mPL1d/DQgdJOOJyfdQNtcLnEIfQX
IN9RB6yiMpvZuJ6ead8AgYZjRMM80TAxQ/2U1YyVfTzPRIZbpR+wlYavOUcK2kZO
mNGo5LWrKcejCteyJqab4QaM9Q+uOwkGZb+u0YMJlAConD91OVINL7i6s5g3r7V4
8QLqe6d08E1od94wpd+39zCiEYSgf9VfwotjrCUvgpjA1h3gPxkMklclkh/ww6O/
8t5WHAGX9wknPvEpJ5I8u35/tJ9VNdoge+xrsV7wYzNMzyET37GhZZmZlxuHaflH
QimmKAdmmr2rh4t8AdxGnz6Kq40mgFTCgoiLiqNG0p0dPfmOd6hgrYCE1Bks+das
VtBzplryw4bRteO9qCxN2XYX0l5snmF1oLQEGXJObBcdAncJfM5QQSs/EVYHES8C
MytjtnRErf5nPqGIQI+wzib7SbzIqqtAQBHhIukcqlFvO3Ppoz3bjZFClRLJ9Lx3
PA39g+FaHYwpNJuaPBxiSzUumGFZ6KaRf0+zbXJmC1tK2vrhuz/4E6HFFlkTT7Lp
hD5aFcWlWOj1jUvIKAdeTTNZfWe+Ca3y8Un9sWtjnrydNpSCIrmhH2Zs4/RSs8/O
aHgol9yldLpnId3R6xLiRmsM71Gk3SNyDrVLsBTmCXjWYilOAGEh2IZZpgToAarY
/Z2DFrU6WKKvz/i8Jy/dd0gdPP9PG+hXymsgMAR3nSETUo5n+m8VmGogpx+32kQk
XR21rjvJdSDXyWsbTNOiTHExX+9f6du1wklyVTOlSMBms/DxEemdBKFgqv2X9kIs
XdSDqbbJQQtd2lfLOq5oOGCHnIbkHIdeFmcvyKhSpBFvXWR7lpMDMd2/4kRKWzC/
KKPF52iK+Xh8ggoeyrfEs9QMAy+wJGUD+oS0t8xdXGgIwge9XcgXuc2/9hpxHvrH
/clggXkhXVIF64bGYbvj27yge2Ry/I19qSrt8efRKpv3PikwmDmOJbpd6mf9xvFd
xJafxLPPJDYuNOO1FYAGyxf/7wNk/WvRppyb+GkuCNCvDEw5NVLBwQvpxj4M8y1H
QGITUrovi03EuESs3LXLvCEnJpw6s4th1C6zV/N7INRFWbnfDCJ8xnViHI9yKrPV
SNxYbaz1CFKwVdZ4bLLz1fWv0wwoy/hfR+HFhnaMg+FsdOVF815R6DxieT4P7LVD
FKvEv4P7bX6o/tJUp0fmtMCpI1r2iIa/364o0qr1ZPZtBEVyaGEm3fsPlKAmYB/Q
Tt98Ceg0XVmj9G7YK4659jf21g9ko98TvZP7spXZV1F6l41ifQoERh0a1cD64pRm
a03EYipn7PsiSoNGbetOn7Q8ZrcudDtTHEDA1I6thIxvtWIonFPfOxWEVHcj8CGH
H8w0521J1Qx/BQsvDt9nwnBo2W5EH5j6UVST9XGSfin46RacV/q1/AFrgncOCPl9
RO1J7w1OtgxNSbYywj3hnJkqU5PVJlqk/UMybeySe6f853anS5DIwwWKKr/0dkhV
7KghKv4YiXkE2F4u8WnFTzH0AYBy3a8KGffeJc9499L/RpRzn5rm3Rs11hOYMscZ
ExHG1RJStAC8QiB87Zs+FAQS0exyGAHPSP8itNpD68tw30JK5Uy3tj2g6K+e3Bak
tcWvYTHzGW9KG6xRKnFj2SBm571mGo3kG1G3leKKsmtxBHG8f8QliRilADJUgwfj
KdNkiLRQV4lzqbSrF6i/Pzk9MfE1mNE8AEM5WckzGQX+YSiXIxACpEwEZxdT3Ji5
j9RlG0rvOytdAShRuWcepI/UWWeGRUk9knRZzNz5UyE01tZMLsvhVxQcoal9rNZR
rAhe9PsN+rm+yvv2cXZUGfK+cm9rLYdFaTx83Yyb6kSivH77H64edutmtga9e+Sn
oPMwNcLBklEW2QAyEenaaEeS1j4b3S3uzjXyTVICSnxVW2q8npI1UnuD3v/BX8DQ
SChiGI36JLOnnlPK0uJwAvmKNL1mabsnyO4HaY4JH3NfInXDeMWh9K6VGcubs/W6
lb8vhOXQXpf8prnpqKCrDIdkr+OgqW1WWgKpIkl4Q1RWlHQjwT6lnhMM6hAiLbbL
hTtJEJtHvcF+gBS8fGy3FXeBIdWXeEToROpzJz0ed6c+dBm1ReFA0RS4TmCDKvDh
hg8JD92ycC7ZqPNXYc2bZRyqlgr8cn+cyTHv4hsWuloP0BXWS3mSOhpB+/UZBgA5
Nx9fNj6t7hSZxT/wa3pz8oB+lyHF0q70a90hx6bs0zk9cVvlWW4P7oPRXn1lRTnJ
XfXnp/6HZPwk7OeKUOXun8ZlKXGVDWHtg0DnZ5c4SEt1Udi42yRxhxT4UUKykAes
4hIlubSMKSmtXjsKHpGenJaTQtJ3/ug/HJovkEyAkjiK7P+JPuE0NOuR9M/XnB4E
pyqiZoK5XDQUZTd1CVNkvFoVQHQmQ1OGRB90uZACufcdJR3oZMTnL1OZChKs7VFd
GuYou1aozBbNV+euZyE+RvYzBsSU5Jknbf1BAcTU+Jl8inD91QpHa0TCnO3LcYB/
coeada9DQgNHVOkR7b/IOe9Dh33Z0jcV1C6D4LUqM5VFRGO8zNKS15gT06wyctNM
MWnfXcCMArBwxmUMrRGwLo5Gc/Fbc3mEEnyNJxqN8TOVnXAMSCfjBbhyzl99RgIa
MorH/Ys7u8SfxeEIgUvUoxkbLAWr90O5h7pjYQTTg8vq7orGL6lH6IYxh7WhZbeN
Y3pBan/BmpaPAXiNx0lnqyOJL3+6IATPcWa3SwWc0YQR/Pq6GXj4G6QejnHhulSY
S/pTVlfgym8Id4zfHgFhZE2dR6WSnBw6wL3qF5wIItOSY9CzJln2Qv+bSwC2218z
jmbUj6DllDkvS1u1YQIlgNHW9MtAbI5oGBGoQMtUEkFSdxH1XOCCOrAMZvqq49JE
lq2v4ebup2Qf4uYBVE2qBBUthMdwIlZPd1d55eaB+Qx7xBKjitG7ICNivjGBJ14R
k6XsSzb3vEFls4l/iB6U8Z6914sW0/9LMN+TA3H0lY5w2YbP75Jq/NCyjFrpM0kL
UPJFXOR1X0RV0FDqim6F71ll3131QOwZ1tV7EbfyUksO+0SN6KUe9KmoDGFDXgdm
luZoXoDABi9xxyY0Yt2GpMz1r4Pn3/VNQfpnpHNOxvk9rlWb+SGZGEtT+/Xu9oSP
cfs9iO+RSUDPtD6I8s4h4Lo9lhsMo1wshHVE0eP5B3Lnkzp/+5biD3ANel68WdFf
GXvNegFTlnfbSB+fHOwfEzr1QQGd7H4ZDaQczsD8SYIq0ixfYLEvU+eOHN6AdNNp
W7irsY6544s5A14JOE7UCEpZtYN2YONfWsfDSGkhxp1IsrUCD4TmT1tVVubIRf4d
B2lbAogprDMS5imlOCFaGqGR/SxqrughzQob+gGP9/QguoUto6zNLW2HRsHLLBGW
bL8r12JZ5/1jV28EEYh3/tzbFR426GW3oUjWwi6hDSK7QP1g0crqp4zAhcjL6z3U
l/gMiEKyk7hHevXSyCREdnssJntfej7Brkovb32ndU/5OPwGzneT6sphF0PG4rCe
zzPJlJvweVhz5wF8GqONu0Yw58HfGwAC1G/knZ5TizT/JeqqqULpyiPW+uOZrqCE
FHw3tVjJ2KN3XBUd2LhsLVwLM9SRV8WSsd1FTMhxGiNvD+FNOj3Mso7+dGBH5nzi
NwSh0TrI97S1tFnApSoBOyhT3+e32AXAMY+Fap3W9MEj5pq0zNepZKcAZuzi3fYX
QMShY597WdrtiBG2kmk7MEFdz92v7uX2z7H1W7ST7NxefqzudrxNFFDwCyig7tKN
xQuDYXZF/UjOuD2pc8uvuFEXJgH0/86PwXCLi8Odeuy34x2zhAnvTc7MNvVOX1dT
dM+tgNbeSmukzVySVZgqMdLHtirFk0DCWak9z1iI5K60S0tma/5xOOvpL9SILVbp
Adp8m92bsIB8MQ+soaTK8XtgZvvZn40XsEeVdNyI6RRZFmnlamApkoRX7FWfAnqS
D8IqcbQM5ieLN/FqmWYP5vL1mKKIogGlMArYvrOMjv3Z6E21Hr1/sQPzr0i7aX48
p/qiIUS+f9aypPjOHPI9evGXcNc4MEcndNoxPrsDK0MzCAnmnoEsdi2juPPjpEB7
AVQUKIlowuEk1kLN+LOhyWT8LnqpPI9Ft86BXCCSj+F2iyps725JlrBrF8VkH4Wz
Tcbof1JihyHO6J2zKKBcwgVIvek+kCD1TKFrRHSiLjMMCENkzvyKsyFJY3RMl2IF
8HSPx8DzrWJy7bV9wG9iWeR7Kk7ERfAuaVZrWv76cpw4kY2SRW1oclkwprDWVOwq
v3yNkWV3qo8k5SYvB4utWxSaypgk9RJA/4/Nl9MnmDrkyHrCQoOwuQoetpfUW5wz
zWtGORaVMtTIGom++41vw+xuSKepaL40bPBxh5DH53+CkwXwe2SWWBco/iroPIdn
SKpwb0jQZsFbtHHFzZ6re4bXZYVvBgvZpQGaL72NWXVWJNZpxvlfVkuc5u+STdtn
vDZqxUmKKUkVr9ZYrv8r0CYHD2Qovncct51xz9Np4/j0WKnpMQ2StrRy3ywQKzcG
nMI9lTeb7ozX5UQlkaLJRwnpMtqjzRTXPJzd0ADyKONc/Q5NS2MPYOmx8NF7gvcN
FUFtykwttV7Xh1N71n0FztcySv5PQmsS2EG2ClWrWZZswS2bEp78pV87QGcro1A5
rPRIRClQ5f2qzBRfDaeH14UcUMIO8Tl/IBobseH1csEll3DnT9TJX2seujjyXvYa
cq6Ab0xk2SzSqmVrMpe+8qVRGZnjSyVfC/dhx9HVJR1TYwN5n06ERtpbafpGjPgt
ERY37EKhoeKenB6Kz366hLe9wlmV0zgCrJyezCBbLmlHBj4Jte4DHfqzDQSoRYTD
s7vrFVY4l7AAT8oKc12ko75B8+x3Jc7jkmyIb7IvbWemO/4HJ9Bz0xIqYzEDoTIw
Vn5EnjSr2IFQTImaFOQrB3wVXGLhuHAbjQB4Nec0cc9H6WMqv0enguh2BwOFe2mX
z2V1QJ/CZxpgMtHvL1E7lh35FeZZzklv8ln5aaBpLQsHeJtUfAMCMQffavUEP+dt
RT6fpV1g4hL5GYgeNVU6kyLSwOn2VgAZxG0uhXjp6EZHS2vUE9sF5SWEIkLF/L9J
ayU2HKMfClQHfmC20cxt7pCrqU8SMVEMJnRaDZJr3GprxfQKE2tPW6K8XoA+Oelj
+P15IuNPHEYnJm9YQyTNtFK67HYnIlFgzj7YpMIlmJsHfeN2p7KKxAsjsPKjjl17
bLbMHmqW5lLK9QzkcmVET2mJzCVi2Uo3DINFAkM4PqwCEodv6ClA/u0fKAvWA/Cp
EuQJslrMH7e/snY9ggNwg0fisZaHhrbKgGWh75sRJ62utwDUjoh8lIdjWYQMxKwV
flf2185jkDq8aUC0R0ct0oXHPtDvnq/wW475/Rzmhn/0OC6gI/WVETh0AM9BKtNl
sFyvQXPJn/5xetxNS7o1I0QynnWdzqWL7Se2u2vWttVPR7Aes/vAUKTP2jEJYaG9
dAnl/3zkszbzWQVBG4FX3tCe8/Vr6L42LwutSRZyzlQ8T/B3jXqhdxwAqO74s5/S
AorXLm0Frzdy4PPY0B/89xC8Vl9O+RrLTfjYgGKndC2HwOxkGllUYVm53RvLWFpu
T94xdz8LugzUIZjFQn0pp2p5SRzcybjXz46kap6CrPFs3pOgVxZRkwpFoU3Rh51e
wV981b9Nyj4PeiLRzOL1gBsi6vMwly8SsQ0oDSZWSSS9XJie5s/5V57/BfCtRcMa
nlFvdr/nMiAXCxXJG+pzJ7p9QSYGl/Sdpb7RrzDgvuy6cuRVr5fy6oYuBd+XYM/e
LeJ1X/hoQLLggU5Stek1IB2z3X2EGVD5ur3SQ/W+xmrB/MSlUlpYiqtJMJIgptMK
Ds5XCTBOLphqYUaAehkePUUgxil+1XpQ5Et5022ZITBSIYh2P8iVjGWpv13ISrSw
cwr3822TTw/MymEcs40uFAO7vZw8xAsENsPPZ/DRJJ3ggbthCFA/Fq0XYZm7fSQN
BGys4gryOYz92UuIdYKG8hB6ao/Ff/PA9zoed361da9uFZpj1RrT0eFrmnWFQAwx
GTGfFoDVfz1RL09thcqg86plw+3yznwbMHwQ+uLQLUcJipE91/5BTU18GOaqTiQT
jWbKS4dApUQW64eHLjYs4J5/UyNWmlpGs25Py6JhR1+MW4R8S3GnaE9O8h1ceTED
QYcFJ0Zb/tcu4tYSIOik8nFiQF/CLVcDxcv8drilAyTpm49QViAVCK4+l7U41Bng
gti6G1CFlrpxI90YASFxk1hLPbepF70qxLPd3Ww1tTNr4+fsCWhxzbtLl0e7bAQY
bYlUad+dPwO83bWd7NUbk/j2+6OV7Rw1Z+Fr0Cu9g1wiLvV6RYbc7rRpaz3+b8/V
SriylmRnIZZCR4zeWiFPPakFY8noR20ipQiG6s7nJFBdWILQOWTXEjhTzwC9ll3R
OYbbZTl4llyIwjj/Xz6pfVvIlrnCD7UVcAfOlFwHPZNTPMBSIMgVt9QuscpS1jy4
TUR94439d5pTZ5DQbvcUKMOyi4fE5DQSM+5f0sTAq05hzedS1Cy5tFVRP3yVFd+D
Gm2N5d/o2rpKgbuhZKTHlxGlUTQzMHwjScf6SxaLuqMr+DSDOsTxLTzlA/XSnQ+m
BLesQ3JORf5gBkF//C+x5LAu14ws4We2eUV5KpG1epwcO8i+rwqN3PZOS3Wejq1g
UYeJ+U44GksgS6FUPJPk4vhMuWCmZy/QwqqpIjDpYSlmOXiakQZAhZRLUseUXaiF
b6vpL1FgENxH+QeL751PjjGXhtchP5swqibgkMz61aywTv/EQQCefmWZ1HBkl7o4
UPHmDpwhvuyObacH+owf4takVkjJ+IblhWTX0HBs2bYWGOEY5AdLLc8WmAJdn9Zg
uDumQcSHSzaeo3rQNCqT6Zdx9tt8KRb6mbpbh3g/sEJyP+qTgqkyGGEVfIHLGu7j
dvKCtI50nJJXSHmX41c13+wSSV38tgojvhUWq6O4rBtwenD0bSUD8u+jti4zV7tx
pvdb0oXUSF2ZUo07hFy7L9hXjquKMiWbk3SuumjvUI6akyP3jCTfIoUgKu1S6S+C
f+2MRsBb3iiBgWkq6yFvLc4r43sSLELIFoZEgK3vWpmTXBRJ8jvNZN0F3WRlsbSH
1TOO6j7KZFyG4WTL55+kF6RBazg2QANTS4IxmB5rya9V9MlTpdSxTQ8j9woST2LB
CoYaz533zEBFAb3BcIuZAqgVnscUfIJjy+ONLbijq98sf/zDppsjtTszu6yFwf38
HiCb7p3MjopzcMSauYqYK8k4ReLHE3Ah8ZHzd8vz2AOhXa1HxItKXpmvPj0iAexc
X3bW97cqNmRbhWwSURfrFWCgpMqEhrj65MYns7qTPTYbkZcUDHYF5fUsDIodcu/Z
W8KwlvAMZWNxcoxQZKZ5W3M77bWI3fIgAMmuW4id+i7zGErUM8+nurU5a3kDXOdN
Dc9fxR5bdRjBYY+CPxkuqXx9kN8hCAWowhrGEpsNSBh58pbJMU9pNFLXe5K2YqtO
qPghaN0T7bkXvIgAG1DLiOT1z1r0jMlMf1U0D8pkLukql3m1WjW7z65/p5DFJSuS
Vto3G/1FnzgbMUDpyb5Nw32gfOGxrBaXZ0VY70FXUNF1VbvZzfKX/749WAxRWHQ7
S/HAlXRw1U/r42wYk3DDMKOK79kpHPVGVSyhqdt8BCSVpyyHphcSjWTeCXc8SBi3
0gXp744krrih6/q3k6yCrBN+sZh4sed9MgUBt5KLLkQ2pFD8q8Xv8Lr4HJbzAcHu
sn/5F5sUUBr7keO1Aecd+30PQ4ILCeD10MVmWhB6IXuyuZqhGFEtT6iy1UIEoOqZ
EF64+02CuzCizirdM2/ep6zn8X0EUc9cma74sfDzzZMOoR8jVc9h1uxRYGpcZSur
+aqN29jpL4tHaOqzolt+Y1rMWsQL6lO/UglaOCuMA9MdC+4ZlkwBWfvLZwJCXFhu
dYBJEOw730rt0o0S8BZCEO3cx7dmFQRk8MnjsabQ9t0oEo4XgrlXOvy/i25REgHE
OThMivXaNJoA5iFK91UhiUkwyw9g7x1TWgZ8GPetkxdXGFl//D6VEAyyV2m9F+aL
SloQS9g/Sn0QQ72zZhi/nIN4GIJVC6uQLmZn/T87aewPZqYcbPsmp4zk6V2wl1J1
nvAy/fuIS0pUUttPf71ldVJpbg0U6Z6Xy9fPQ/ABz5ZnA5bt2Zu4lUuETCZtf/+F
jgPOKcdlYqaAL0cpl5wqAzU/2rGBMxxxrnCg3QLHpAJvAynn3Y07x8JgupmznT6o
gWhft9YLcyYnrbZrDGhTZJlbkIWy4oiAESBIXl3/p21Dzt2DZOIojk86B8p8h6AY
GQEX1QTcx2Gu/nP3HZBuxKH67USledyzCPSLLQtwkQs1OCCRw2/vP4sO2ZetUbZF
RSxh2j8CcodsLCHeikAMkQWZDwS/iei0q8jy+d2g2oU7g5ty1+5372Z5R+IoHaAl
5Cfr7L9wUayWqt/KoOXuMpD/YEKclAjJcfKrngGGJxRIk/+G1gRj6e8Q4TnwAq1Z
W75n8E88lqAx20/kuVgCTsP7hs9z5/0PfnG7WRQfe7mhrcVch3SPqcPpZ61WBU8D
BDip+JhUyUAj1hIyLL0dL79SgcPFEZzAERVprlAqn420yAtAL121nb2N+xdAMhG8
bbGT6tYwMrmEA6HR0K3295z4PsvVJEcz0YRxjIxdsdAZSIiugr37QfJtH8VmsNAX
JQFbpxU5hbV1wxkUWD9/bwtJS3B97849P5K8OCz56pezPjhCO9rSKAW/mWUBGvj9
XdLE55Pr1rz1h8+kI/DBA4NHMkpDM6DvKl+vpshIEALyVdQMnORUg359yyI8PDS9
o0Qj/mjaPJx8sPBB1nYzBPBPnJQffdaKoVpEnqHryxRKlPxxIJe1TvuGymGbPJvn
62CUt9FxQYQmDQoso/wvK77Gf+ZRvNLOOv9bNyduo8RGAqhEAOnegakdk4uyDcvz
ymZNPoYQ7W1hRjSPNiebmJlsgpbeR1Yz72WViXkY9Zicyv78fG3r20SSXqTFnBSr
Ir6gggjxPeRcIgDdz9jgIHRPXkjNBlR9tL9cDx1mWhVfxASlKA1fD8tT+o4zeu1g
dsGGg2Ppn30EYQh6/Ig0xlZLlv/q8I8bjLMmjI42+Cm5IR/+2mFmoRkaBhSiLm4c
BUCmWSwJN0zUYqv+h7spTy/nHx5nNXjnsP37C5rzNfCUZ4UopFgl8+iXspIN/4J5
R1QbSGudOWSfLATOJkbgTZgKgKtuDho/HVYQpmTemDsZKwx8SIgn8OdP6yh5T2F+
aeG2rhGxj4mAnlAqR+CstnqIc9zyEMijzwiM93b5dRJ8Z5MfA7D3rWzncbk0fvxh
lDhlCPmGJFQXO+TYC7FMt7BA1+lxyA9pOZ/tiGK0nnt8HpasF++BMmplWA4amIMD
EnfqlRQL7MuxK3Vc4PAeYSMJBQ5+gMccWt8xV1zgvI7wHaLtFWSbUWN56ZuXNGv8
IUtpe52KFgkRADL7gPJrV1A6+A5s4obLOPXJpEs5burLMfGhEGSmlTaaRcOH2bue
K35IAs97wwl/+tDQXkwHOh0IyO03Q0lb/kd0ATWMX9KmtVgNAPijFHDfhEMFCZfp
NWzqyvwZLAAKblC0DhssCJZ1TAhjFDLj+FqseH9c1UQl3wKUMr9eHIyuDJA1rrEX
JHz673v4irMwo2igHkEUb/fzlyTIELqoRsWpBf0AN18B0mOWNUGrOoLFYUaQQ+QZ
DanGbIlYwzUEoV/7oLlqVzNh1HIf46bAJB7dVgULTEp6ua679nohGUpkkY174xp4
MjDUdB0kCXA63beYLKWCauuNb9rqvqY/QLrQgYh3Z/cf3AMx+OYW96gTm2T2K7fA
VnzYG+uDZb8v0BmM8wAggxr8e4X8u8Y+TQ5i+zZ//uGsCsTnYoc7dqhNxdq1ZDki
8rWx56efhA5ib5SLXcA4tQQ2jeAqI8CW9N6bMI80smS7v1v1G6ffjeLlF0gF5SDn
vfMvEvKtBFjrZs3bAntyDzwFjQpvFzoGzKu2H/miDJOlxHploEcVSDEpH7bsxQwI
W2V13wqBVIEqgPesE0ojS+UzmIkehNxB73XczkOuzOGUTpeJQQNwUuFD8iNa4YLp
uXFFQuApkSleEcgcb6DNYoqKQFbyFOfA59w2vPgntTAtWeu1O+RpU2Mawdpo+6ew
Elo54UbgaISBrCcv9yPMiShxRdulLFKr+YKMrxQBKjHKp/VjbGLHHav7fzDBnjd1
k7RhiI38jwpR6duILVxhE8UTZ+IwF0KIvoSbthFt2Gr4YLeVW3C7OSoTged3oW85
kxH1LUa+weqfBQYPOIdutT/Y+kmrYILRkj/+p0POgeoZiEYr7mofzwacNWPURMio
9RW9bK9Ni2f6Z3NaqvNeaJyrFin8hZzl3NrlTQM4g+YlOqgb4/j7wwIOHI4GnvxD
pETxkdO1tQYmiRQGFQgCxngBfOm1I8jlp4chkKtVSe4FtF55guTSp5pMULw9JtW6
exmC0TfXnLX8xrvTJ3IUOkL7RyqI2yAPu/L36WMxEueRnQQFfeV0u/lgqxrRmvoo
TNhaZI9pH/iLH6rsPQDUV/GMNvQarYc3qM9aHwBbsQfMYXfzCCC/SvxQJMGxxYeF
LuL84F5XOEQPWk8mWVwKvgQG9e1U1IAGi5jXqIPQCpMteyuj93UYrFHGFey0JUc4
bPyyE0+kyANhZ9vewpTv2U5+UKWC37MU5M1x8a6j79BngcQfEhGb+nuyqPPpZOU6
ULHbiorggtBvDoxfFxk6x+9/FHqqbyR9g06ph/z2awYuMYCHs4ndyNw7YPofoNC4
WxZevolnkv6zPhZKWQi0fWyN6xcNUyfJsctZtcONBRzg26XppARf8kgtVpdrGNSj
zgL6ek/HNiv4/2puCX6zWdO81oY2TeyyjVnzzplAnPgRmmB29ln4l1vKrnDrml4F
ipeEelt3lEx8qy6cMnt+wfwJIM7xLjTkerK0Yqhv9bRS+osMFZparKYzFG9qCzWu
APX+GMDQyCScdQuptVF3M2cdbR49kDzXz2g0CJS08igaOgkBb+39Z8SsKTBTlT4S
2sTBZRKIysedTioVeDT2y1r4k40YQBWnv8RkXasM6+tLvh78vmbcXrfBB+BjAhFD
nDR6cy6467PE5+0NGu8+DWJzBI7YzgMKANexPH5KTZGe8noKcgVeCPWnD+OHTBSk
K1IDZkqtOb21DxNJBmEy7iKiktBez5MAr8rAggzJYP33QccsIhtNWm83CYQOqDwv
2rAdQrs6IwA+OGDye79f1EyNqDpC6rt+D6qGSQ29i9sNu7Sp62MRVDRkJaEeb7/S
GhcIgxr0+YsAQaPjIasulCUurM/VSCflMt17ATJtFjZp2gDyBug0V8ZAzz36f4cN
WcIwRR5BkLby3LFubGEmeAOl45JIyLgl0Bgtpx+fHg3tso3RkBpPexlMc1FRM9EK
CJ/QLxCc4qtMwQgJ3wBZdKZFneB2+4poY/GnJC0jhwoH2BNKfe9MjGbsGOL2Cohb
ceFyRGk1yJamlE5AwsGyTMpxhrgQRVip3Wsm98rUipMOO8Qtf16RKIPCtZBEZGNw
xRi5y6paFDz1BZp+Dcm8cRQ/0YcTXgyfcvm+iKLs8a0KHEw8Y7pKsii0FYrNlJ4T
KVECzhfvHZP9PzOET8DyrZGHM8EFzFCrTtgsrUXC0Y4SzDippXuthihD3n/qgZGF
dF1Nh7K0/CRDOtJiaqJGikbNbPFStuJADFCYA38QrhRCeec12+lkPd/1PRVh6h+A
vHhPjdhHIMjt3qCCxjIzByO5DRdWBCC6/ffnfdCd9wlTuuT52QCuby2OpuW3+VBJ
bHI5pftKrZAkDz1qh5O2AkZewoQU5WM1KfOt737dKcB/W76iHwKG534pLzvcFin7
t/rBzHONl4qOio8gDiwrp7Zu6oEFc7OBWlGHJJkAL2te5Cm+euYdM+q8lucIZ3Vt
bv66ek3c+JT5ZV+UrVfl8bCucj4TJl0TydQTT0g4huAoXjG52puxtnQkg/9s8kuA
sY286dRGHmoeyLZTP8ipCPnjC5ro/kVQZ8ExefPCAaSkEJxT8lskV/IdrSz+z1Np
m7LsUJ367ElDrXCm3ctSGUzx3a9Uk6wbu+syxQEvs1K23vIkEAG5Bi/uU46RLxKd
55UwOBC3PhqjTbJs4jT6agRQJfWhLAPc2vWxxcyR8ZmTE6+m0mh559J2/CrtA3MU
pPxDRwC4mREE0AH55hmCR6CBN2tC95tGpx2tOrnE0Io2L2On1Fo7UJcqJVX5+J+9
Bv/zgiFr8aJxUcCgdNIWvMOpxpJ82sjIm9EjaMTxYPeZz5mw9TVVjoV6OrUu8nqE
eGpEeR6Sg+5Hq4szQjJvy86a5RvLOlSoaP68UmjktmDYGbdOa8g6unVJ3aDY6KMQ
pUkkYWRumFoeMD5JtGMsdMtZckd0QekAxdFLeD2dz0A7pOZnBEr82UGQqtySZHQq
sAkgAU4cerJCXu/K6Ne/REWwGd2yl2tb9/x0+uwmWW/NyMXHu8KqdQc0lEQuqo+O
FUXwmAJxhCXFnAMkJwqElJhTyv7Z1t7fYsy97Io61AFjh831RIGQ9QjmsVQ14EkI
hLzNB+h5yf6mNH76FWHKtoltK3MDJ6pMmNWJiw56liv/TOFKHHa6MvwprbuK1GAR
jFE9qHQ8F/tZldOzcA/QDb4+GHPNeyryIpSkcLdewUB+CT+Ph3BcUPolxnd4BqCf
CmqGS1y7cBOgRifkO3VQy0xec/Q4ER8RnXtAlxA5klrRdzoe4PWJUNo4z27eA9qb
xgIxxdjXQqOdVe7urFFJKGuArHwElPxP10t3QZVKQiQ1QI4Zm1KxtZHsc9EQV6xu
r7UdQ87q7EXwLgB1ifHvhanwOR6peiVGbSj9IEBXzQYWjHVeixe1fEFtlSWOnLAf
NjyZkabVUFQL38Q4GkQ+yaNX2hp8VNEIAoKBYOh3UKLmo/rSzrFUyZjSkXqPF/4L
3fzvpK3l5MC+keXADhPWDeOkXAYdkJcooE2J4ydGeKoLfKXgRQbaZPo+wJtNzQ6H
bNlcuGWQyztHI42hNkgfR2xoDN5yQEuSGUtzMlIaci23ern0w0BtFTnpzlZQ+Y6U
u/bg3Y205ClWOj+mL3RV8V33Wx7Q4JJmKHmUA6mibfQnR/0Sj45Kh7mZubIe3dt0
J+bDG37DSeHvtNreeR9dxNvUi3Inz0JGxBGPKOV7lVkg5hMD06TwKxsSvUBNQrhf
kXRIWOXL81AlosVvFaQ4xDvB2jKVYVaIXREL0+bLz/uVESHz6pGaeV3JuzQPsT3w
o8H1qtB5neBMIvTCKZe5XYa8l6qGq9IdKr3jVo4hPrIIXVArBFpB3d0uvgYooxqq
w2RXA+gwKDhGU6BktFEoIlqA3Vrpq3AcUY4M2sKV+RZNj4GhgHqtXWlGdbVIlXWV
O78eDfr3/HNmyr5m2jcA9eC0y3BzpI6ICXgVkXraPD/S3afqOjNggmo2XB05ZyFv
upO2/RwmIWDARiGdr7vV6E7Q3EerHt7P3Q0PLOeFtcdeciMCU5UQtXtnaKekofXK
S1SqiF/wzh6ZZo5ZEDottz/8M1P9EIkKsALAAWLj51Fr9E+HusViUvVxPgPAL4HF
L+wJyi8TNcjupC7NAGJi+yTXeWO6wlF6cfnfq44Iz5/9SzDWN3fZ/9x9U6xz7FEZ
MyMzoNqScyRsTtK6K6x/ZrumX6upqcPHpUkOYoiGc5t3Rn5bG/UtPDs0D5uuxmVI
NSQwQ6hoIBW8rTDj85bdTJP72+AoiFn66mTT9K3xO0Vf3PDITet4t1372jD7Xq9q
lgEtglHcH+KrVZFRskHig1lvIqvz1Mu2zwqDAxuARYSFu5/IuVJauBsHaWZ38Up8
/buDIwVqBSvsCSY447LY98dGalviWloLq+wt1sszfvD0omxHxBsaIw6JmiMJVnuq
qMLtordeJmG9IYsbAJz8aYhlFpd6DUOLzcufcUCNwxp8e5NowwSZ7ROdhvh2oiNP
AagnaCpnnGbGw2bqfTKHkgqCtoTSQgtnq+kSGiNIEGgPCDkwQcYQ1ZkN/wj0yTS+
VAKyQYxIgZrTo8U/Ymu5Bz5+u98mYx+ElotyJnCtul823WEuJjd23gZiNNMSpS1j
0n+iogmlB46DT/7cNKS8k/kCUzylHFD2RVXx37qj4WaxICclNtUhtUDaFOQFzp+G
01XrL6nTU6WQheeRZT02c8RUHCHRHz7woc3HhCkWPFyncVsa7Ulj5FdS+euyQYT4
kjxuQF1ooN/HWqwoAf5u5Da1QfJJR6A3dYSaKriiczsGdOPlGmg05P166hEHFwVL
FcmbUC6CM+E333Ue+NVZ+G8IY+h3jDkJQ/77LH5G7eiMV5i/9WUl5fqSwOL2TBSq
olxJ6gNR7/vlzGTjTW7awUCQXXUnHVDz6h7r0EFXo0tNO75El4rlh9J/vLwLbT5w
s+bweh/r36rIXx1vVeO+oQsJTyD4bnSTErUN1p0BJ8M1di1/ucyDooZxFE57ftjZ
2PDaUtZ8FYA0ZYlPWYu89oWhn2uI30iVBKLZ7zhf9UxLA2rHF6BdQitpKTz7X+Dc
fy18EcGNIV6Urtd5EhbZ9IjdcUI2Yb0JzclYbg2In/71HyN+f8VCjM9hfyAYpQiV
1nU6rqH8GP716v/1ZifvURjATiJsV6i3ePHA/h2qm0t6ClaPr/TQITZGzP7zZPFP
ahqihyVIEU2gnRECWaXnR0neoH1Au9uysJKBKl1SH8ocMwIJ/MQNzhA6qbuBJyZO
sZv72JZCff4SoGvidu7zvF1+yhXccIdxNZfItzH09bfhvldWXSrI8StVUPh/BeIy
YsfPgkAq/Jw5PRCveea2rX+mQaMFrWDXf5bunS6Plhwym6vsal/SByb6RHf4Xl/P
ZelScyo2djIiNHGlVzeFpkwJ5yyaJbILC3I/gVx0dwIQErHNIWOOrfC6mdc48DJt
T1W7ZM3RmMvx1yBplD7AVD/yLZhAEjzm6P7Cm4pR5QJspS6xTrcLHu2g7gQROitq
iXavP2CwrjLt+VfZ7RCTE0DifYFoge9FhF6bEboUZNcD8FV4yGbffw29nn2wzZRu
mZPDjpiEUka+60zk916jjW5FQAj8Out2D/52ZjIQ4OjTr2OSLlzjm78+/w0NmT4y
q09WFKiOabuOL8pwtXXF6jtuNjKyLZNm3y73dLGS0MeLA8E/7K56GSNEihD24pcm
D4LE59i7V0oPrVH7aUdo1N75lrT6TDtb6nlAmQm+u57hixOjeLS/q5YPxydig/V6
xNXC4F1p7i+QCU9lWr7SUv/RjXJEwMaydA6ogT5Rb5bkMfUPmwCK6SeHdKkLgp1H
U8oY3z5K+0RMAnQYopqbAh/1CRnvajNKcHj6pES9AKo/qv5suxNx4otmmctrYoZl
YHxUT6lqV1WuiaaS/rc0CvFKRL1FJLPDJwODYJGsxyd9OMIkWFgy3lj39X4q3uv/
PCxUAjHhom4zPQxo1t5Ni7ON1HFayBLcXEcAmee3gPSTUR3t8loxDu8CvPxLDI/W
X2diQeLPWEKikucuOtRFSsCG8QoWbwkGdrs6SRQ5ha0QsyLer/Dz8X7sV/MnJXNP
OxDdC9oh1S3zs7IsFmgy0nZBKATg2I/NMt/uPrsagdhLewglSSPauMFrT6225+Gs
b6TMJyj8kKzT3Ory7WdyYJpIpPfdApBGH2o0IErMWDlEpA3ZvpJQP4onmbbf1lOv
YwTuWaFpd4DLfP8NDYtRLoXSWQj+OADB+xF9ZeubJh9LYjCpIZ/hrLMNqj1omYPy
J6jHQV7jFMZWwROc/x18uWvAKfbYe1whVwgfv7HPIxaML5d/GaYaJ2plxzyhaMVS
vg+a2lg+eWBHaTabxlUxP5C7eATkov3rhfu333K4GPDcimy6CM+/4Fcm7iiuKf31
JH9uf+sf1qkTPT7iY/tFGqKhJtWi0ZtmBszllQEYeJHdEKTFrsUYzSQMUhjA5Bub
qg8D9JnRoZRAA3ZCYCt1VaMX7bJWmNgGWAMbGAw5p2o00RJP/ko9dgeQ+gGDclMc
KFGLdsK7499qRJHpXOD6JkX5zmAXuAwSe5ih8CKyHeroBJFhrVtSq2siT5WGCsdc
yZHxaRQDqyQAXsY1Yk9CJ1PSWZtWnsgzW7O8b69u1P4R73rDnOIhTijO9Bq/wlE+
1CWIbn1W5khKDEETqUuIwBuAZ5FSz2HYfR/9kSV8LpqwYcjF1PuUHa4tiBF0j0Ea
wE1CexBYtlODKNf1Q2zlDZG973AWMSUjJccAd0SXAgsfuY/g8BsSDP9JqRKTfenW
IeNpVbkgbSOzXxw0bHKiEmq4SYWzrP8U/GCXc3NEzUq3qxjVMRIT95THNyGCHFyC
oDs2dAtLFcIWhnk5bB1iGbrgludj+GxbY9wf686V8kWaD0yeOdlaZhYcFtQJpDYg
HIKSpL6qaVZdYjGeg37gHjafv3h1KlfF1mUfyUUM/vfzsIFzSuotL/3ivbMwJIRr
ozv1tzE5gHWoIGLbvXWJ9j+2yWSnNFENYG/OrtE7Py7vThQHaFQTMb3t+JSAWQ6G
hXjSMcnQpzfIRKkyxly8KV1j9/GGBbnvWIALHLHxlpiM7wnnfKXOPwI2GVaddtn/
pmEmI5muHRmG7lqoalXK32vwnwKfN4bqSjFsngwcn3+g1/copnagjiZn/jkaieJ6
h5xfIq4M0Ul0sB2c+uT+nQwJgLOjzjvfbGKKx/4MbiNqhLTIUSa3RgG4EtoTZckq
C5ttWKb4kfRh6h4pIMwI+eAphcLh+pyBXjFdtHwmCuhFmVMic2vOd90oV+CFJvAY
0O9pGPI55lkj99T+kk1Pa/TAR6LhbjvpWDbR5d0hFAe9tEUDPRueJrC+0SXkII6y
rjarcCjzZJybkKuyRZW66xaNECrNfka+VocOj847gRi+Z2suWH8eO1gcytvmrl3Z
qQdJyNlrGGrVyqsCEm2XVTlP2EjjLI0ukIcGv7cSKLSx0Wq7YpAKKqx64He3uYoh
btDFQ5qZlWfoQ9MMTZ4Yl+UCG/gz2q2IwNqXuOQ5thvAFtFMdMIPDmTJEtOisD47
r2jRAZbAszArs7AYYhAmuYXGIe8lAKVyWOWi/HPDmU/+jANyoaFQ/q0Y5HO7ph7S
+k5dKTLOX0hWNwJ+TnVN3cuH0q6SzMu5iy8qTweFGhVF57Smxoin5hBtHU7hLjr3
OmuuaTtMY7j46P+9dRgLk4Rd7tpYV1CMLp9k59Dy7VdZqlVBPMteqRymHrfBceE6
29F+3EsZpnHMXDrfKoSV+EolQtTxL3bsjk26EjsCb6Vnk4+egVmP6vLuQsnryGXu
1FHICYe84Rnk+1NNW0DmKYpzQNfOyGsGLIZc0eqJIaT5Y24MoT+tp/aTGDDdgeYS
4HMri/2buJou6/ytTRSmcWs5OX6cikuYns2WxgQPBZ8umiYv6qQHMZSf7d2c9oqU
tlN09DRH78Z+6RaJWiOyTEMK/D4/hV4GaRDvJXaWz/4Bgcpe8kDFsMUjwcaNg8ju
mQ63R5GsS7aeJA23/R12vW9Qt1HYiKxcDFHB3YEt8T/41NGd1glTB1Ri6gd3P9lM
tNtr/MAeSrWWLszjmDcLaeg5c43WxWCaveZiZoN6iGU9Ej2oU+5gMfcb4SMzhWrI
7j909x+Odb+lNdBQg/FfEkI6Ssjb93Tq0fWdpeGCy0gsqrK6H8N/UoeuU+qbNHCu
q8B+isOz6dJ05rY8f+PUOcBq+TjHG+hfKtLIZXMbihBGIkddaEcgHKz+ZXwjOy+k
legqRu4h1MBMU5XeF3GZfyP2/YDN1tiBUik4v2FuV1an0LC7rml43A5t4oS8fuSr
ffh0zUp3MviwJPpHmpZoBU8xT/Bc80/gZbL1y83WWZizz7Ev4RSlEoHYBMVsDqkW
oiA0OayL7H4NrCAg9IAZcc/0zEtO17YrDTYKIscsQfi4qoCEDBWzCUTqLl1ZWQBb
1CNRw+rWo7kaxVwJajICYDK7y162P7WU7e1cLeCMrgSHCoBFGjwIuXwdhLxL1Uxa
OuloA4J3IpBOvjRfikhjwPx1HEtifH4bHSFAUH/4HXgxUz0FSdZhMaciTigyVkJP
mqgaRCDaMf9bq1kk7IXYJ3RgEpPy4FbJxvoEF8zY0ZPDpv5aW6Ls4nFfh91K10NB
FIg244owPc6A7F+2JY8SZiws9abrMyhgjTuVk9tRs18QbMlicD1MtaMtBIsebQyU
ic1bCd3BtEtTWwASCeOjimjuGR1H+TAcUIFab35M7YqPTPw9nSxPse77W8c4CPvA
wddh6ThGtXtblh5z1P/kSVLVQJaetiEC0dvAXUa49SNhsPv/E2KmFgtisoLzepJy
QN+XttGbZcsv5MNG5uG5i7ZSbyZx53fxJH+EFQrmte8O+hvpxRfoypp0MUYE57gQ
hUQN2aYSPK7yBr5Id3U5hhEAlYI0B48sW2WCJT1XuzHuzL767VF3G9/3Yx33xNGN
R9/MkK1Gxh5uZrtvFyG49VA4ehfbiQjX2zEEjnaV2ctNyL/Or1aDovgD5P3aMwah
vPvugENM92fEynHZTi159cpJ56PYXDl9TGNwkCjK+IYKfCzjiMXliRP3pD+0eCam
rk0R/f6d3nkZ9hWA57hhQAJW3xcn6KmAbJ7ON13ydQd3tTl6omjiN60r5kEC+LJu
rJBDfEkgphgEM/AeZkMaHtVrvWnNndm6N4jcT5v1UvoKBqly39UdliNE6AgEP2rK
I0Mk1NSJTaE4glPzWIKb3+4C5n7GA/LC6+wC6PjKA4uNfd1+qVzCIu2JBYVGDqeu
FwrUMFCizp8XBe8Qe1gJG7nxtzuhaTYUojnvbVY2yQf40a8qj4+UIBoSnreaSGe7
JkBP909n74Ulha6kDTeuuSuf/w/YjnR5pNtX8aKgJT7hNqnTlffKL4ufvzhZ/oHu
pwIEh7FU+DxowZ8OwqMuRSv68kE9OmDiqkmCBfDaeeY1bzgLCF54nLO9USNu/12i
9mar3EemqaBH9W0P74MHMLfaIE9fM1o6HEo7Wv1/LpsuHt4RIC/XNmP/u0K4NU8C
Rcvt4RFJgB5ygS42TxnNXsdjH6Lmfni/o9uBgZhvlw1JVxYzvct2YAh2FyLZ8wBJ
6XZtzDWqKMXLFGqmi4MUZk68Gr6vSOv3N7u6cS74UO2PU5bjEQdxbupqArADS/6Y
kz/lvgI5nXrU1L97c+CUkfJZMm4wF8y/wykMX2R0h1XFt5VZOjbgnJPWwcOBftkH
HFmPg93uwxLYxuP47NCqEvfzE1cDovs/GdoKYzy6i7H3seWnc3e7ySbGhhnrnGvO
rMp3omiCNsVS22p7FkzGmZH6RHKt7+UOQniz7/ThxlOdWxZJlYY5oCaGd7jfGDKF
3jUDNjI24kJPQHCbFt/oIkIJRkcweISrV06iDNGQifZyxWxE4HidyG7GeWEafXq+
3507Y9CY4T8lz4ByPMxsXpyNlRk1c0IPEz48IH3eB6pgQz+gRhiFETdZoawGryuI
4zkKuT1bimoP/LQkQTNcCRN+iUPpWBvBeh7v4O2pwxbCJBstVMmUUmaiLaLQjKWH
sN+9sGphAPneYrR+gycvd75qBYIpkDIoZ7MTGuaItSZ3Ae6iq/3WrBAUXEdMjaQ9
3HDo81oh3IkdUs3o6vF5d3yVOElaycA1eBu4Yfh3ozrflpDb5Cq5mUFYAqnzf4gu
AM/a8Gc4FUIZTdEt0qgvo6keDA1UmmTYGs2F6SOX6IJzxjQkjjWh0ufG/kk7fBiD
Wmu+pFcons4zX8UU/3mPMiT8amp3v6AssQ+zVEDNo4Psujh7D4McQIMYzBR+B3iz
pYH0awJEKlqR1jThBBC8hhDGLFFvM8NHIM1Khdg53h9JVFx25+7Ds3DwO2UL/uMJ
7Nfd1/HSzWfzX/MtZz7+Hqgt1sYlKBpx+9sYKRzb/S61/+yDMKUZNjqMlc8W92eG
6JL212rLHVhS4ds80dziSdH6J+YaPsutIkKqQguCATPW+R/6g6pnmfOT/ZnZoGwM
aNM/9yUbT5DEaieunZq9+nT3DcF7PMnXmP9dcus4HTCMjxpE9LzLM8Wxw6tz3Zhj
4wNG7eZ7Qw8DoGcbRjJiLBYmpmwfEBAazDToSONGsOo/XAVUbnCtqqMvsN6Nt1a8
zKo8SQIfLoaIVePrQmkXcUcWnPH0rw5aaB8G1Rrr+Bcc9lrM5/QZhZj+6Dwxt/os
LZL+0/5/bwq+Q6MRW5EQ5Ho5M7bsNX81cPAGeWUPz0MfwnACPVTv25M0C2i+G+/G
ggzSDvM8NRfRpADtKuAaydGpeX7BP0z8b2PdxIhfHNcTyEmmW8b3PkUrqMYZ314R
so6n2BFVTw5tuLua+kxSNou0is+X61TFhkYE5c/Iir0WUFiJUeQf9FUkTZ4v8enu
D31BunEma0gUMue/Ezd1fOvNOYfXeALDW0q87QLTv7AxlKpj+r+p4kpZuHwP3Q1V
6h0i4OGgFR79K3TSv8407qGb3joUCA/OuDj2Y0sGTDxntjByGNQmydvEYMU39NV0
dfu8YD3mb0f8mWxK/E4vDoSAzHYufawHgnKS89m8C3YA5YWxRXn3PqMfHC/GptPV
ztGhFy91t0MzFDFp+Y/ICmmczbYpPzdBm9XWyxXNDta13juq926rJu1gNCXMcjvA
aUs2vVbMTAia3vvamZ0URw5LzUdHwWevkPNhX+bECLsH65A4RVCMCowRt1vP9yNS
uO4QOHxcmebF++RM63jIjYxGZbrN22uhm5ffY7ConXU2R3bmSuSu1pmXffCUQTxA
tdfl3OCaYpuQxfDUy6C0s8eG70GyiIiZ3mfOyxSn3BT9BCFObBrcPGnX6wXG+Prp
kcqOy9dLere7KNpLAqYKLmN7pDjw6B5l1lxbJsSrBO6BbVTINBVHdwUkZpmNjCCm
XvbF2kjrwd88qe+VxDM5VE/cRIuCPqJkekhc4Ld7h46oMUnAdfoTKOkUH/WHbIYD
uSatFbK0d2YMkmbeU54jwpckp7jtIJdemSZFA2ezQCdbAjfhzC6y1tE1Qf2bfBel
TgD6b7yvCLP6mTmk1YEv9w0V8g7caDvmThHEMmT4Sa7tUVhCPsZaiR7iaJ2bjle0
e0XrnRZ1HIge9qiyuBMSEXUVK9CKHDFHfMSErB4csLuxoRZRZoqMOx0hpjkhIWIx
z/kEndqxxcfTLSitJQLMj9jv/uO3A5NiDbjdHlA5r5E/nAsmKho7iPVtD3HL/Y2f
2jdtPcFx36CmxtRN6ejXOsev6FMb9m7zmkfyXs1++Z1XkP1BSnalV1S8NIl/lLb1
XRpQa+oaZThUrbaUaAcZXxTGg9PFn/6ceB+4SXx6EMxbYwduwcE0ZNRiVTIdHmFy
Y4wjKQXo8zJf9h14E9afbXjznKvQ4sY7lr62S9FTUIm2L/sjQ4lqPi/lj12LiQpR
mA7c2MCOXMbDcKha2z2GdPqA/Y7ZqyJisQ5/4XdEJ2LMFQShKdbYYkg65y93jCYX
eWObtkvm8k20XD26GxnQdV1o9keN2OJp33n0vzUjphjw4t1O+I32Tqs1Rjp6ZSaY
vO/+ROH0VnMMCLEsvZGcH1UuHei2so0NEQmTVbPI80NNnmYIyjkOmT+/E8Vol+Az
r//Z7i/CRn1NkGkmBLUaDR/gv6r+zxGJjHYYdZ7qdTgihwKxragNxHy1GkeaB3s/
ayH2Vk/E8ax+jFP9v6WMUWiZFHrVLEvy5xoMtlSSesRpAlh0QmwCNzlgkdOxXvoB
We0jvdB6vqVHVZGuHRswcU+htD7hsUEnfJIx7iUzPKGVSzTY6zoV2P77Vzp/zD+4
7ZqGdYWkfyJFJSio0peZ178e/KWmNwODvhEUIoTiQS82Ml7wKIpLwB/8RkhT4eO6
jirt0cP4ZBmCpMaCWirHjR2I0SvA4BVmxTzjTOu6P/fgzM03qLIhJQb/G7y6PdPp
U30Ow+FcEHwdMq88QQPp22Ix3dgFMzDNTHVeHU53qqofKTB7EZiHhkHc4dZd1VFp
W6mfBLegZEFBdDfvFa60Sg9y5a5OpcXOC+3kgC/J2P5dzTKJ/vtPoTq0h56mL5n1
rjH4ywRGtTkPgP4zZztZlHBYYAprFE26LLHKf1utko7n6UT0ymv4/+wWwWbjiVZP
4mj/7E3YvF1rq6LAOFteN5u27YbcMga2mugokXqnqXcklr0o2Fye2x4+W/iUy4MI
iFd929/06PtGOssX0/MQbX8nqvQV+S1LUmJLKwKzJjLZHkNPdYdn6jG6fcwKXzfQ
32zPr/m2N0EeOeB5UueC/hRTWDjW1v5TQeay4ZtXASWCRyYfG5w5zH9QV7vHirNe
z/4YF0dQbKYYc78cibiWJzfsiCJs4czV272Kqyji3Qnj6Q8u9nfZ4lyZK7K6QH/s
MG+9RgSTf2hZJGFex+zZb1Zqe3ckzorM6lce8bTDB5kMbVHP16xYLsgWUjOBM2Iv
GcgpOrjkE7R2OrhaKQmBb+YfY+54u5nOard17KKJuVcs/7wiCioAj7zCydMgdmw0
ihQU1Q+kqdtZJEqqX9ENPA1qk6m1rpxT5BAlkUgIbUCVGLvK/CVoq66SSb07/lvo
/uOF5T1HhKzHJ7cSwWc9g445vN/thqUnnFZwAIU1wILezOcWW11TLyb2lsQflqj+
RWCe9CEJ5KETD6QJyY1aIEKMUylXQ6yq3R/CRVL+YG1JkdUK6NqjEDMwSxFvN67y
WHiqh9iT7PwJA4kDYPbjq3yNi5QLLdMK6tXVmMYShGthAnBEuhou7410ykE+IJ2q
cCt2CduVXVtb8y17OQ9LEJBtR0eStAhiZYBrUR4OJRA4Zl2O+7qfW8yKeSWkcCfH
FtBaeeer3WFkfOw28mHzK7bGnXZ+jUoUGkONjWBY/znJ8ZkhHt4EP0H7i/hFgL4B
sqdw3hUvzOd0WeHlXXOOwGYE8a9e9sJLDVPWKjGq+mUCXrj1UvcZrBREYC5xaruV
fuFTXXxXMlv61ne64jr7YLdp996coeUeq/6YwKrTi9029CsQPkgSQWh/C55IeKoH
HZtrsGgrJVSEH0sE08kV93Qwa8FUsAG1KUK01ERfkMIy+ggPkm4gkLj94hUBBFAJ
c3CtO5UWti1T91WXbZzwmAV6ebjeSWXJu+OunndGtXrj1xK0Wr8fmx6MCXD8U2Ok
8kA1NliWzUooqNc59RvsRy7Sg6s6aTg4yhXFEOYI3dsYqfsB8D1tvGZ3dRAiMRMh
dnCCGIgSn84XP+UurZSv61Hepm6O5zxqc9UBPDcLcZVuw8q8JdvAgYWpZnZQxrSH
l9VifZsggHdbHE0YGs9CkEDF1141gy7JtKRaa4j4h7jM8uLl5o4QeDiDEd3Yucct
lypaOyZ+DEk3UYVrHZW/6Jjo8q0Jfu/y1BVkheKiP2Rz0jnE2YsTHCRKkuyW/w9s
cJwbd1DUfYCK2QVHrRZkY+PsRZP1OT0dzTrXNlos8mwuoGg5S1r/VX3+OySdK8RU
/wum695O1AYNbkew671eC9j5qeUjId7W/GhJOhOjd9jHeeWRl4dDPZ8hQLalRLOh
iAhyJflCTOswmhNWAuloe9lSHNsvzriAC2ggFpjugtOmdkjZu/jeXNTdUG1+m7sR
rBM+aRAGUAw3wL4TQs2D1h4EaIqYobYRnUS8VZMXHRsP2R6gzKOMvslLBgAWPPwM
zCHsc/nbV8fv89q8YkZMdQrKRI3wum9rhcRQk6Zgat0Kw8JscLSbC47+zSze/lu6
NVouGbOF+O5LY8AQSfqMVCAOFGmBIuuCcEb9wOfg8LyjS/GmhI4EivXGpuv9yxsk
2/n6zUq5oowIsz5FfNG23NazPbQKKQwKwxKOwWBHZb1qFoGUhda+tEVK5D0eAuPF
htaO35aYNWVNzZsl6ngmZseWL/OB1LjG252LQyuy/Yjy3UBVdgt0ky78D6/VenUP
ThkMa+n+QTJA2dUkqzObLGJwtqJKt8XDqJOs5bIwvFveiOei2Op61wm6b7E7oD4o
DaKGVKrnwahIdzmNhmkr4v1PtxXAQOvyO7kiqzoInju/VacCOgkN6VkOdzY45J+o
NLqLYmz22NYbvji9Dq9HVMtebtWA0+jdn3ve7hLEGozBkkTteii5cnvxsGd44WzE
rc4RSU7zsZxjmBtGSLF/+urrJr6UMKmbf13qqVktIS/KYteE6JauViXLawhAjJaS
dOVN/TRXe80Ppfxef72m9efcVyOL9qoQNrGPbw7sZx6lPsYZ9Ut2GmA2S06aCEMv
GiyzplJtgg1r/a/4LsxyzSE6gGVXJ24eMtUl2wRFj7qQhZX0Y/urYDQBiVRK/l3c
4a5lXERXZsrljXvAKu7e8EDXpPORL9UQmL1JwBUN2u3FKdiIP/yAuDuSfb19kc5o
sVpo4DkNySQpZAkkzJ+IsKegB+tEubPNOZMYuhB4zGWxWngESC5J26e8EKbdsI95
rp5lfsZKcRS5s9ZNw2aQMlGxqudZ93P9IRTaj7JxIX9bmDp0WPGjM0filvb+hvI3
HALGtvWJlq89W1pDwNomo804CH5Tkpkow0+cWvqttM5x8TdI6HXXgBRF510O2w5i
EdEkZn0sEOiJErc9Bj5HjRygYPrp0DdyjdECaP+gBsKdBt6jvB/IH/pt8ETyQYb7
hX456RNiCztn5E8iu4TIdKPbgQGqWrnTjc0IGgpvSBhVHymqz33wUrLKNPWqpqjz
JuodqCVRLSJWwwntr69QohaTTe0pE7YcqaaKpjWHKDgIjd43R8e2bITh4rr+Pu8z
FwCEyNKLk+jUfPM6XdUKjfjEZYyEPA+hvfPtmWdUIW+Y+31jC+L1TVxg9oEmzui5
9wr71j6UpPkMOCO0WwAr34cixgu71WGbwPT2M8lXAo4doBgjpM1xr8B5Z7TYP+Pu
x8m0jhK8q/11z556DSBIUMWJB7YMyv/uNF4CQL/PfwoNkPo/4uATtpwWmk3QfMfF
nYgVgBFjmO4bHg0TbODatjpF8oeoJvuog57iilBEYXHsom0SRMh56nCPJ+XPcNyM
4GngNX6W3Pa+dlB5T/UwyYqT32frzqLG+ndlfMJvfjPnDTC6NPi5FGq/ZBUVyo0L
S7o/YV6KeWEo/2aTlnpG0XIZ6mL9siYcDqoZxPHL9nIRhAq2BsqoqWQbNQAw2z00
9528kp1LiM6uPtA8u/SKcuz8Y9hnA8bxpzWnVeeI4qYuzns0Di+/QnTRmogMXtDn
iA1oGfUSx5+XJzogZfp9ziZnSJ4puJI+K0gOKjSsVEajkQ/dPHNYob2yhgAgKU/I
bVEDOW9/hmzeZ3oVlSHuQCuAIU+JgKgouBdKZpEtuGS89l18QcYGM3kKLzfub4CJ
BNx1x1So5djJoEeyo2zKbWG2ZMjRDzP0eJ/rY0W9e+Nuhoqz0FeZzMb9QGEK1R9K
Czpc0C4kOkqZA1HpP3RUXttmIfI2BkxpDrJaWVTmTq8S2BjWEqgRaJxZW4oVek9j
LwbJuPVNH530fb6jLpdU8VcccvxxhxUGpLAN+XlxH85Pan39Q9Jr2QbYTZMI4jpG
7qAutIdnF0uCeYHYel4cvvy1/lYDpHgOiVDMwdoz/ZJIqWB9f2+mlQyDBk2xvj8J
1Nj0glpsP3A2H7P5p8Zc0A/N014oF4cQZ4B3XaKuaYCZjQIoSb4ICKUndJ4pCAlh
wqfjyvPlPgD9VG2yNnmMJnKTn2ILr/xZjmSqRHvsTeh0U8iSrqZDD5dgY6aLkwik
t/YDwjrXtIiksU/EXIvWAzqfFplTT7wPSUJKJFTH6JTEdP3rXE//DF5wyUGP4qH4
l2koK6bDat4rZk/RDvG+OfvjZQIDMa59ndhuA4r1k59l7DsBvG1xSbrlZflkNX8A
IDqJtAoAeXuWCMRT+fpvXveiieh/iHiVVo7loP7g47Fo6CVyLHT2Ga/oiC0Nbmkg
kVLEWeMHUQHAb6wc/XmopAZNq1gUZ0FfhYQfGIIFIQ7NDuoE6V7ctvSHcKNIGwOR
Xy7Zr8RroiHaXJ3FDI5/kSBR37JpKaEpu5WfC84KdjceoBQvGlCzrjZhuCNJo5BL
rL7RBHQ8BjkJr9+K4/IF3tqtIwvvTl5mo9jRjdzNMX7oHKhZ/S116zMgcSlLs6L0
Eg0eZWSh6oeIikwmY/c8QQmYzpgkUFIGFOdoQg/AQd1xOS84UR29Vl11gO3SDYmL
ZhSc2/wMU6nqj6DKuPVeuUXj1/7GQFSaC80Iki+rVlYWI3NojNlVJzL3Ie80/RPW
y3TC4ICW9/8iqrjixb7PHq39GNGC3NCwl8y6Xvm5EZ2Da1ftNkADqSlCGxCsPILF
/0ij2mP9I1uMkYt6jJ4urVaeDQgr0J+UKdICLYWorLctzW90jcj+yq/7m/sw/PUd
xU8kJN9UqiLd/3XB8iwXX04sT/YsFx6XQHLL05XqE186rYn9CL23TPNxqPiYpDPh
MfxsUs8GD6PxhIDNGC0MU2geeIFQXXS5Ia3z97cDqoQGKL17uhXaQp6bfLzDph4Y
vUYrusQI2wK5Cjn38wKK+HpBlXQlWmzJhMz7xQG+rrK4fmdctEtuHthTc0MCL54c
WgytaddfNjpUT9aYR/2BlNBb9LeH6pQJ6bmY1wG8kzZE48Rfer64QyQ2jv435xYI
D2HjXZtjMhpZqmlb9vCAia4sgYI9q11k/rJNy6Dvsd5FcH0Wr5/EOwgV9SvJQtKs
LvBa1LteLjbkl4uSeRvhGYKCy9B8fTA7PkD0F9okbIaMXsL+nOC91srnXv+73NNK
r6CwHST3GnvDS2oukC8Tc9NjzilYXbTFkcugrgPYV6iVc+hI6aw2rWGUnEtADpmD
orPakBNt2z8sDiMkaYdUKxCaCQ5INykZ/i5CUQvRNYH6o0/gUNBll6fr7Y/DzCoO
2VSht0i1aJUtZy3S/fm8beYOARgoC+h6B7JMZCzOmPgDAssc+hUQIlLarlZKMlgl
jo5a0hS96man9no9XjSOpdSrM2fkwlJk6cKHkzkJXzgnkYzXw7C3y55PvwX0tJMg
6X4ke2JiuVTOjfVHXNwPkklyiVrX9MfTrGJ2bv0zflyVo+d8Y7BqxZQ97JnK36aF
VKRX9vZKu2s8uIFVze7UbWgIh5ecBzhkCY8fVPwCZ8ZpIV7raeSQEL1sWUzbaIOo
Jl/VM5bXAH4Qf0ra8rMymRzFIfQW0cWEp23ovKZt1F4ig5EpZy87LUi2elzi6Qyx
jUduJycD+zH9EVOP3X79cZLgSggYnqiEtcSRQmZQU/91CgJsKkGjzWMvwfM9JA2w
q0XtJ+1Vp6C9xne7LE4SaN5MnQ4409h2BP5rtMwfZ3CZakygC6qgFbausgJA3pAM
FZNFbeVdkrC0ec1OEtdjG4rtAuOgRTmGQHiI0PCxd7KU8xsUGOEbDq8btdk+sn2O
WLnDORIgKL2foyblvrlRnlMZUgmPfs4WfWVdbfilO+NHCSDHf7NxoXa37zFuAhUT
QbfeeEMiPjwU6Wfs8BgHaWCZ6qctenPPSg/H9AMPhvl9zjpaHqGo5YUl0+uBQcsD
XNxURrvk+QFiRyKvyQRsnEWZ3CnnAdc8A1TeL7VfBtzVJ/g/NxRaP58DenFsGZkH
S6b5ORAP7A/OG989UT19yNtF9TVpmHwQOJqm/O1y7I7nIiEL4nV3dBmGEfncT0kg
k7zUmGnRfsCNphcvNBJPuyp35uQAa9dmMO19BJatEawxFD3z1VeV5SEOd9owIgPB
4Dz9XIDY04taKIBgBVmQjCoMDgK5PWJWs8gm+1LzwSz8YZml6UKIq0Ccye3VlaiN
CnLVL6Igvx8QBT9iiR4ijc1UJYJRgcbKIa6MzRUo1AgB+JpSqonjQyJfa9GYKwmG
FyHLy08mVP3uR8P1dfvI7IblD9/QZ3yX9CLP8hdG6jxFWt6XeFop3o+bdy0BcMBd
ghNmw6o9neh+cAAwhACRyrLZrvzzADDauL5qDk4HG5yryLFjyjKH6KyI52x3Lrv7
5A6bAwBAjAbL3bt6jorzBbs3iQT3ha2v/XpkGL54GMJwGzFuZlLgvtfOFxT5MsVL
RlzoaQKkdlRrcDuKQpwnd4oRgN2VKvhpSdjDD+7CgjtI50jNvJbxQshjVkLoo4Vj
rybdYuMwddJRLzLRXy1q4xhcNP0uLGGq07PHovOhxvXhRHC2OIv55g6HSy670qty
/YvoaHhqCI8tkdHH0jUz8dWfwZ1JvyqmLKl76dzKK43FlBNIKE3BUmIhkXKQpQTH
u7QRphGhmoTfNF6FsYKTzLuB53jffQFMARwUNW6Ijfcl80I+2yMy9NsrHLCYTY6K
RzDqo3FhkLeTF3xUAtk7PRw9fo+FSU/aONDEYYnsblg6M9c+4JzvJtTKph2Hi1lp
lDQiG4zy8RxkNqKtT53NDm9XW5bmGusD4YyMVLeC82MSv8YhttrmCmrY2f7bZdiq
eHx7UkvEFOh7K6zzRcAINwQqKEURclhmUX2SN7Vp8sIXQRHOaCjEiP65Tg9Q88mS
/kUKc/cvIFeAkoOllh9FDj6bOiLpNzCSEEIOuh85GxoW6X3xCgzBoWgr5mmnPkmB
KSzHSlxQql68YdtHt7dHwOpd2K7Ac8u2VbPBUxlNf98nX/sXRJjPsSDyHunqf2gP
KSm/qCNvQ4HdT8YWL9SK2C+6L7rkE7B7MvfKLIZAmrVxbzroOHh0Eep8Pz4Fy0pn
sktHo9tAh7CFt+kkJ0rui/JW9KnTsJdONVypKv5E/w8j1cnO3BWYxqoiIPfKk5Q8
PA5omrUg/uUYw5ae14tKjKNuiXkTdEcMQ4k+DSl+WjKp7dGlxdWjAiPO+RXufoWp
QHvrmTyEywu2eA7q6ILY8YYAC4+oU5FHZkKb1TE22WQWlezvXi2QUOE6GUKCQp3k
6fTahPJuJ1zIuBqBqZ/eREDuG3H1GdwQkF5OlHz51UC1XOfP3SjybB1R0Tyhb3yi
blrDZAFp8QybTM/eATL8I3WkGN3BYe2g2lT2NoYj+RwxsPFZWGPaCOgsCyZXkZ/J
xjxZVK2Q19K13lw4nqIo4X4+AmD/61k238SP8dw5N1CT9YwgKQuxeDH1+H/USuol
Puwk3V50kHgm1dYCSIq8SitQdySkubQ/k1be9x3BOM10mI3WfK3FuXWB3gI9tE/z
bGc4sDiziC2XzEr/7PgChZJuXKHX+BLq0BLm3Ei+mf0I3Grilfe2Kg1N2ZK45JVF
mVjGBdT3dhE/Q2tvCjC+O7J1N8ZWeC5Dg/UbPlAMsw7BgpZQfBr+eVfivAE81b2V
ME2va6GIo+RS6mJngYWppZewUb4AqkNBhVnLOPj/yJFraPbo+DTJm4PmzRRiuPNp
PZ13w/Wncu0Pn8QUTTJzpsT8cJQ9poTAovouIMtIBmTfSUx5Fzd8QvE8h1YTpIWz
gSAfS1qOk8y6dNaVVluyPmO1jvE4QftD+Tb3un2MNNu/CJzXRYANfRNi9ugjtqn+
rhoJ6twBWtRXFSerGtNlOSR0exy28hSrqlv0nsw1YJtvLYgYPIE7dOSE3+AFrLS1
BZWaJBWZPHVoYWtFdAuUxsVvPMjJY8jqxOuEf7/kPkMLxjwrjtBMx8xxHs8fMXCx
Rpoheuc1/yNSqalUslhImbonElyU2wmBohCX7/4AwVIGXi1hqQ1pCjElwSk3HWyl
jhiAZWM0zW/aO4v+SSVvbK9xAQc+HUfk8hHc3BGd6xJWG4T7hJKPjmJ1r8WX6Ioc
bhi6eFmwciGCpWIAZY4ofOLsIxChKFCZcQnog78QgrIcV3sx+PwKE+25yshgWzko
fwBNLF/IDBeMn22Wqq5LKJ7tB2LiOkyjzXZOSUcoT0pR9R7Jrj7Lgn0Ury7gB0d2
f0SEhITVo3FQ4BX89zNiiipDez9QvN8bFRj91Do1b8kt5y0ndFYPsVkyS3lXlKhG
ABlj1Ug2wjz5e2n4nRB0kxjfdAS0aNFpLzuNJV98RA3SMOWC2qwbIOq42tFHKKC7
EjQrq9QPL5uDOiC6LcsFynRxC2O3GGnOMBDu9am7R6XlIQ7Ji+5trCfNTzAsibXQ
FU0JsjOi0c5hxYd6VCioaSg+vuWhfAAB7zsv0TA6f1mzp3yoADVnzr+Pda7mtmu6
II50rdEDfJ5e54rcqf55UBT2omim3CYuJx2+YuxN4HMqS/YTCJPxFxVwVETtqRGJ
1irN9+25sjIp+D6uuWVYI/ly1Bj5RsYobhyUok9pYi/My02RcbnAKTzR3PGNHjLI
JqDg+5qPzSEEj9HJT5wJJiIa/nvms8g3qSE/c8Q5ilhfQ5fiiK/5e8e3+VCvSA9C
gvyCRXloo+NkpvmLSzWlRjPHtg4sKm5SVTzWsopt39b54SdTLDP5T2V6ah8GeiGY
s24K6+80RCE76Xy0L7f9zqv9E1DKl7N3xfa373+QEW0FAUo/B73fw6456JAo2zw/
KaTWvJHdiLyrPjpwjNMBZc2+IckYpt8yQqi0Cw5ygftZhEyFqP3lKlv1IP8CJKFQ
jQJDPINMrYK91gKwiAqBxo77JWqpT+FTX0EWILs2pNvSWpwrfjFa1HyuDtjTq0+7
uigA8MIu+sAtj/lG0bSZvBhPneop24SfAQAjFjPlMDU/A0cF/yiZDJtaD0ifFL//
lL1wDy+CuomA41dt4bFOohmb1RAWWTR7x4Xa4I6bUKKveUuu5deUxrQfPWhYZpw9
7wk0KeDgxYIkJb6/IjNMy0owyFuWDREuqEt6gmd7ba9SEaLwdAanU54OdAI8DHlu
ELRakyI2C/v1hT5GajP7VHouTR/lqVAVI9JEqFoU4CWfnI/iM/1hPDkYi1szoarO
V1Z+qXElbB8gN0nqIQQpLwWxysdD7TUdbIThAEYsHhdXKgnLyZ11MCCJpI1yii4O
oVjikKbGJBQGZ1vUqquMKqpYikEStncuBM7cZED34ak7w0WMQvDk2hIfPDxCpDT0
6xdWwJXPXBJ2efA5UnRfhtRCmfx/Zljr1UZL+1/VJfzZxoqCp/E3KvTSU46CsRgD
iz8n9aTJS9JCmM2ITvUXTz7bqFggth2OpJIpFKFyjEUsOuYIJVt+2wgyGppukRkf
CG9/Wr4GJA/K5GVqq0upQUMj0Gr7cPP6kr9/7nqlsPz4nbkiApTjQBJGa5jQODfO
JV/HC6EhK0cL/4sU/vy4F640R7I3N6doyNiMC1P6+WCYVRMm/BXj8nJteyiX2cyd
5R1ylsBTKPfc8naDENyO8jRDWj2Jk5/hABSygwgOGdp3ybbdq68wkk0rSlhj3oPZ
dhCnqyFz84/jKR9nki3Kn+5ZjPopiMr0FjTgFSYnkt/xJMUdYHa3Hmle7VSTBZ3X
d1KWObQ+6ioHhr+nlWbesqybnVK0YrfEV1KdmFplNtNVwXymMsRWGVHYwHBqapTp
pep9ZG5dR0nSmfWSTrbgKyHcjr6bGEzi7/4mEYVWQONOXizox8RU8RuOitvj7BXw
WGGe+Mlh0nb6k8sj3VwLhl5GNgEP9iMQN9u/eydBA1e0cLxYabpyfMSODzQ/W7LP
u3moK/5muGeOm1JuxhIROPIDwiC/SGCicLMhzm6ZxJDYY9Kr/bXsTH8EspWP3B9G
PqSX1QtVOTTRgYy/d6SR24cpbXV4FEmJHHioLUUGgELv0caUi/fSIepPtFPG/zFR
58/5gCFS2kN5+jJqCGlVbarKvEbRVSyHRcjX/EVgGtNX3orPnkmrVhX1bqasJJEE
w7/xcN+mhB53vJhg+7pQiLwb/rx2U3LM1tT7e8pIQuzl27SNvvUfJSnND3s1G7hI
XnelInAqnDp6KLRnERmLBQoJ9eHTmDWZhek9PVYP7aU9Hvriy0TK/21BMikiBH0t
KjUDCLEPl+Nllu6L3FUdJs93RzAgjbYpVS1g4ULbI8o7nbaIM7TSHvduzAdSni+o
L4eMIHYR4UX/u6g2ltWsRta+JPhQTYOL6luAH65sXojtp1fJMe3acfI+i2676FNh
Om2+eDSF+mcBPxK0gRbogz+3Oau8vQupPz5wcM4ABE1RQ79mGm/HseoOOhVpydw2
rDQBza/qkWu3Doa+iRAXWazl92x2g1/KD4tpNzywOI9CG5WSME0ee++Wu1kc78Px
Y6nbvt6czsB2qehSQjnK5ehgJv3s3OlHRtc4Bo0ElzjuKkE+mNOqFUPHFQymnp6h
OnVLVe8MAPSX/WmvU/Hz6RJfoTdMR6c/NUwJhyGSfXxWDaVKKhjEOhjZN/+a/d1W
2ffXJ8ikbEKNER502hYx+rWB7ETEfhm3YuCOOfgJltmknSzSV/henKfmD6wd7Wk1
qjPiV0jPbtY6w5HJ73+ughaWReXLWh6QpPuoWB1Hp+S2O8MtOwtst2T0V3+m8iXQ
SUEmUomZpOcUcA8fFofPzj0KT+nGOd5M/X2Vv0bEvFh1hi/XurV46nYJRU1ujauu
2LygmGN9k1PMpNURSKbk7IGx3Yj1uMNpNHYsXH1VZf77sjZNnZ3ONqGurY4ojC0t
nxKZtkH4T3km2nxSMX2J9B7DAix9GYKIvDT2i+io9Bz5jT3cjOGgLsfeeHAc+kr/
lI8Dd2LM4wdQ0/CoMBpSs2qzaAqLy6CpeDOwLiDugXJSQ+Gp3yx4WTIJgs/vWXTE
y5092x9zFnFQSgfQ4ZKrjl4xMxpwr327BnLthhgUhYAuX1TIV0+4jjFn4LsZyJ4O
uax72CE4bn9qLZvWzHys86blRO1Hmxh263ZrX8ErMchDemUZPyZaAblz63EJRGkA
4dVkzQWcVMPNWrTeOIhLcDT604EQ9y2GXmeCuLpPiVi/YWDZtutRk2pYIdcsMXLx
0aORa0kRB7peJTW2GqOopCxFOTrwhRmfUEF/2NvchXoKFYhCnfk61BacwptQFUAw
OBuko1eNNH6J28PIdiFBpYIexAAsfiIK1YD+59a5SvvBGMEDRacbvrDLRyhPOvty
d7vJxLiulVDbgvGJiqIZlhXfcek4dugdLKnGg+Z6nIM3NIxiYidSIx/cQAF+gNkv
S3OnyKSA1028gGMUQrME92h26Y+xiwFoDLNlNu7AXDcbd8WAFq6lm4WBpnsDxl99
D9g+X3Y/oLmrrh7uvOAMSQn7oboyPiy7bTindDBBtphy6pwM7T3PEoa46Ki1GnSe
p0F2HaJGk+/zJJ0u6jXGedgZ3ecXwnDFqSjNU4OP/eIRh9ITRJSt5GBrKBA3QgUm
Pvml2HYOk+Yu901eN3P8Vo9Er7SmnmIePdDWP8FLJ4r2LAqM2frMNa38DKeTrKq6
sXfKQ5Gw2DxNbZsQeraUua3aWjDVKemt+/4grTBuldGAo7ruqwdFPYCZ1r8SzOMC
3A8nvL53m3qHxghmZ9tFiXY6XtKcvBRxA/sXump4468eKXe+JD0GORnNF2q4EV8x
rzNF1I7C5LrkzXk03Xv70wcaoQW1TTbdOjNsK+St/WcBuSI7F7zZxV13uojcYyto
fKE51lIZ29S/o0KeHBOVd9mxYZRZYlhxHjZrGKjVj/CNzBzNnXAGLgVgYaWxbHvB
C4DLdAw+M9mPPPQRPdtXkfsebxGr+jTEagYIRe5AqkEotgXxxPb7bZmVADEz3Bwr
lLLjGAvdTE2Qc64OIZasuKd1HAXFr1n4L3W2i4mmDxWtptJazk0l69nSaCTsR+PZ
LOCStcUY2NJyvST7WnUHmS7q/K1TdmavWmL4X427YEI+lCpvVVirqNsvzgtBNXjx
VlUCj0NYEo1FPbD+8CqfhApULg598pcDjio3Y3wViSaQ282n5O6K5v0vNpc+G0am
2pW808Bh6VkJ+O2j8O2TQ3ag9e4JNJs+zC4rZwz/nMoA/DAc/RC3iq4rWXlScSyQ
RVjLZVaTAkxrxwI2CdyvLYqrmFUvokEwfvoRJtMoIUdUnO/8pnLan3KPZNE4firq
9QlfCsByLQUwMrG+ZyeJ5Mp/IZn0PXMpFuldgbCfnobHRHiWER7trsopqH8YDiIm
HXY1dbSuzqkSF1nagUyolJLLEWPzPJV1fH3hvC4U6SY0A4l4hGlTJRGWNrpJUNrc
UXK4V9udD8CDLVS8UdDwz8bC1R8gLMMs3UHrxSfwupZU3938h/sfQ1prBjUUm5nl
RxzybROK++qEOECEBQkkFB1TKm9X0f0WIyOdbK2Jp7eTJMJrIIO5hwB8yTXV10pw
UbubV8h4V2vkDea6Pjazmdeu/INVxAPPhy66bMhaKapSJoMWZ6wp6xCmTQ3+EwdY
C5rx6A6hsciWJssaldCXHiEOLtey2k2LY2NuS3nmm2IwuOad7MYstiJXOONyPR8q
sSvUq2lYKua4fXOn+tJt7rpm6gLa4fPF1rIY2dQRYx9PZIl7wLVED70pdngn3pJT
QGylAm1eJCP+BdMQJP2izBJb0wSpkTmjhSKhbkv4a8mHeYMuN3UM12oDDKdri4nW
6EiI1s5i/d4y1+90LTkEaFWDC3RFdE9y3uBgtpzbO5MKnZZBs/b0vJ6Zqax9VkPa
SULC0dxDarIWcfTsCf/1uSEAuwQyQn/az0Jy2ag2QYXf7P8wxiIPVVr63UQPCTZY
MMQUsCHBFwd0GdE1qRDWYZs9/HGCqQsXuBb4VWzZ693qsJ/ZN47ON3fi6e6KXZdf
qMAB5oBVe9eiSJYB/moyvxj0IOjXQTudwr4cusDFeo2dSdbKPd1w5sKZf7uk/oVD
TjWGlKzKnoWIwTiKmMvEmqdBkmAzCGquHNd3sJhuSjWohYLlDls4p3ylSjrnYY3r
qQdAuOWQQ0wMDvRn1CAp7MN8b2o0wIHRdRAlyRI7gEq91jgDK+asdBuBJBwFEHUy
TmECtLZAF7LVqSxxGRys6RLmiI9P/ncJ3/K2Elvy0I7whSkhKCza6DX/hcvug51y
qATQatA8jKd56+WVulhoq8XkCbv3Lv0lIimcQ+Or5Ex0jLhJ9HckDz+9KvHfK9AO
7sbXB5lSNSm3rZHDNgnAw+XicSEk0JZob6nr8yfRJu42mIhoNyu1ICwgMLVQ/hAB
KbVMnNI3sPMsBtUjgSiZBml0rdPM9XWUoFxnoAnjj11qGbpwqgoHSJgrMY8IPv60
nE5J6eT0zJXGQohdcB8phaUgJid2cQmFKKyi1+ABtXG/5jumMgkGev3F4ULex69U
Hm9g1IYDqP04KUD4cvpzq7m+FKxp1BHjj48QdO80INGAs4gLFTZMMFi8xBEgw3am
qq3hp+Nxd3Fr1Sb4nbFowmlKlRp/3twGlIK1JLLoip58C97FCSkgGU+QN2N6Jnxc
CBYhFX17zTOZ6QePiflngVij3D00WDBdoVVTkeMEvkg1g0RWDSlbB58pQVp4EgWA
Ccol3rNG7x8t5QOMx5HMYChkFlDXE52y15oWLNZOue+iMGzSgbIHZy1E4Mkv95a8
MeTEvRTcPw0QzPzXlxoDQtKY91dIkC6NUX5URDRbcAAhkW3f7KV2DBNmgOjS5u6R
ZO0C3IfBRYy3RYkP4ZaqjGqZEQpZw9Nq8D46PIV7kj3GkLsV7uiCX9ScuRe2V/R3
i5SgEsA+UmMOsdb8+mU7CLmUW6twimKdO+MTL8sGYt7k1Hw83ekai9Dg+b8rnt3+
mj5Lb+fXcMDV61WkHMqzyWBIg6RfYcATWmBk2cwdUXZYSwZqb1lF9kIwiz0MCXzK
j8u8/yb4Y43M/xmiI2WaO4if/57K1zNOqAxDTRsjap79+tZtly2WrkSYVxfz8UxX
cL0+wl7kqR+wxsulOkcsMf8cc4s2I4BYtmn1sRmqpH9p9cbIzqGyd6kjuLV6482Y
/7VqlknLyE6DeiucJyhGPkwIksYQbJ0jDPifhcE2LAKloiVrQoMTcubMlguRAlQ3
6iql2hbt1w+MPGTtLepHd4ZO9O7k9G4/pUmYcn43TSDsssJs0bT4BZsDCYgycb0h
+qIvMY1ozzfFEmhZxR5Mw7FxG1wtTZre6K0d1jPHUw+8+E+0HmJ9dEmAPquY2coQ
eYhrIct8fdSMpkudEj2/gpcvxjsGiKRIByGytOtMF7hXFnSAPMwvHKo+ADnbiCNy
c12UoDuQRmc3Myfk5p1HGWdcd3XnRcJRgbUw5+G/g0uwYy95mlMwbab5ilbTK0OL
HkclnHthyxNtRknBgojVl5jsMk9WLJh7y+r/5f/bjO8hlFVEFhJ+1/vxp/2+ChnX
Gbe81qhAcxNPkMrRcwKfKbCll7aZofdg5pL3pT4X6po5TjxipxeDkrNuNcnokJwk
Pc8Hstx4t/wzs0a35tPbOOiiYqc0MdMC19sjgLsW3eV/1xfnN/RW2avjZdQRCjQz
KiT3VIIcFpjj43uY+lzFWhRDJDV86rAomyOj81Qu78J/UBtY2sztpyFWZ6e3XHex
Woj7WiEruNJSyQSHycbjRb0cmQvOAgpYo1E8fe7qxgy5/0lWJx7hJk6cSjT6O3OA
TBjaVxdHrEGdIDQrMYaXtdB80y+yqvDQotAT5cRHZm5cUHkhr3Obpjxl/I9svTI2
dwLd9cCvAhdkvyU09mN57JFE7114cSBcA6jJ/myoQ6w6iQvsLJFIH3B/CNZbiUAW
cXlekyt8OBflFLzNpFNpTUePPoE251EcujkJJAlxoBO5V/NljMWJRDn8Id6/IQED
A4QskcXTTQceQ6lMDBSTNuC0AOa2K5a3cecY6SiBHsTV1OYCKEqprgT8b1RrD4hX
6NmUN+K4tIJEcdDGAnFAaNjS3S4n3Dg34dRNvbfU7VYfhsBPKMh2e5YTEpNiBduF
BST4Tpf7E0MPaQEdixtzWb9aSraIid3vYe1CKFiiQ1Y/cdwbNeZz0zQdG5gQb7Xi
z7wGxM913blW4ENquOsYVIDLOvwMSpvmjO+bloA6q75+9L7tu09i5SjR2SxQFPAy
nCQtLc3e8/gc+DeVmEcT5oUyEQKn33KBxz/Kvvw0LFh90Jr/hU8MxeBNw8KDIFDU
72LKrK1LXXJZ9AWhcqXZoHsd1EmnONuSxr3X8DHCqKzDSvkwT4bI6JP4yY5WFoql
f2n1ogYCesvbsVn39xibX/ikuJyWdFKb4OZq8H8XV2Xg5OkgElNEPPnlMOlHDzF8
wB19jr3/v0SuE+pG/C56m6yH42uI9nZNJfeVPmxaU0ru9sWY6EEfifjK014JEKFZ
4H/WVasUWjUT2eyVWPPAn2zKtX9pJLylDPhn/cx6WTIDaFO78ui5zipOoykMobLA
Nr1PEWDUbT38K51e/AREZ2w3+DzrKTlHHLo2eH/3xYk/A/kBoOpAjwyAEDuoPPzS
iRBuSJEp6mOFmNST5yaNOitIeJ1VhmBipAaDnX/U2I2EJx9wOUKCmvEkYd2J6jI3
krE+5Vq66tXH+M4tTbBSh6rSK4AcultF0Fj9hmRI9lbMla2IOj5yIhMtfePxWPtD
QSj9bl0ApUrygqntbjwmBnu6QuIlWXTaZ0tIEd9vYnTHD58SD8QbEwT/3keqh0CB
LL9K9E3gQmVuPrziFUsLZkjnUsQLSXu73QVg3qSFL6dZnf3Wjd7Trd5QKkbWKJ5Y
/QHY4/A10Wzpj95Pfqv3QYDt1/fT+MJqf4JvxPFe6aWiVFpwg64Qh/qc6+yz2gID
r6t/8SsqSfVmexYsnlX/519ThXPQNrADFiPJ3cq9iEfsnDoLKtxkqoqn1gIS4dTO
pdd/hLwYASa5bFyV5dCFfboBPpU+mEuLc3wcOYyh6LRJZZZCMHyb0ncItnmkInF9
dhJM3mgSbsrvDezFtKcxcEP4pt0JtYvwaeBSkrPA+GETwm2ACh+LozNxizJJSXr1
7ZuJ6MngKxjZIx6UxTuft1G+2tdJqBBoxTJCUbcpIFFMueU9SYwS5u4XGvcW+KiG
8EUJD32/JbmIgmjuw5hc5HPi+xKsGSx62yZLAZtUjuJbh/c7n2tJAqe3LRI4MFH+
jlMw9CtnCNViy7KMD7NNdfPCSsg73Ns4sqjWqrpYzG1/HR8xqUiJjB16UpCXDN0U
iThSd/q8/sQQ+P24yzfhg9F0nRqg7D0/bvbsEq9Fj8uuvyZEtWm2efIK2DTjylBa
B9nI+nAVnrXy5s6lbu3ywyM+kYUlA12lsZy/WNiM1pOtB7Hrn2gvep/CVmwVixRI
p5KuXODH94W9AMArvbBfszYXfT3SwvbMMKS6WgjH2ig9X5qwRkpWO56kW3RUcneI
qKy8pgKA00Z2Aw29Uj0lXhU59cM6s4YiRIWu8dU0n0Ut9qbXzSEzojp6jSnNuK52
6bf/pPiniss4yeuhD3zDIVVHknTFoCPQLOtaF1oqaeB3skjiW2XP2DILV2QaFegN
XrCx37kNVP3kFfPtetd+sleQWGicjaOJrpovKLA6jIOehPqf7VT6Mg213FRsPUah
3gN9I7ggF6hStH/uPvjRr2zBL46RYnxj1F9kYhG8P5rHRlz+siTZ9Mbrhyl44EP8
eArK5QB8MiDvFTKbiPX+nripsFT3xbQ9Lgdogkc7XZ9cN9G0dinnyC15VRWbZTDb
NBzF1t3zHgqMSKQ+oR5Kze3j7zAgFrEW01o8IBE7Vm4IgFKg0CnQyxFpRruTuINU
hQtHkMEtWHxbyDizWh3POKoa9mZvitYZCnC5ftxz7a4L/PszZxmoE7VCary16/ui
OsFtxZAHcFsd5FYClP9IvPSu3j5G72uf8fxpkLeRR+MAFEHeNS8owwSnZ8rNbFrx
7Zu3OpkVSMrV1NsQMiOrkVODtykdbPE+hJcXBlrcdVZoYv6skqdNmLTiUYJU8NB9
6a7q0gxwHMc433IbGPO69wJBD0aSkhD8oYs6o3yUdO62EkjDqnvjpLhY82LVshcd
Axoubx8B0NA8/DwmOYdVi0Bwi8NgRe2wjqufPMX/IqW8ppZrWOqvfMTfKwS3CH3S
CmwD87P7aMxAVx9yFcLsli3r+QC9FBaqoOsxJHIgIxZTUFaGnhHIVbbHywqjFKay
8Hq3U12tJIdkTnpsy1uzZ50Tpiw2KStKe6NURMigf36HwsxOL675BvWMaunJnBhF
PbB3kyT6CF3T4wQstoLsQti+6bvkAoRza2BI8r9tYisGxw+IkyN64L+66TV9h54f
FcqoKKlQUfsVTe+JDQTyd0frdwQh39uzn0rKS8gcHosu/F7Vg1UcbqIUQhLFm2k/
C8Xz70ZiI2ePRdYE0MCTRDt/3kodqnuFF3aC91Hx9pTqzEEqQGAez82Dzsq0zre0
zSDWEwccBO19g5tidjbgGUBAmX7CZgo1iHbwUZQnX1yUDwfKVDir3BdxR6TXif4i
4Ug2Ox/0DRr5FQPZ2uPyKr2TDjprQq7hv2eD6tKHhjdh6cNlwtGno6aVm9n7duI8
wjkckl3c4J1Kvp4La62JFiIGIUNFFogSdf9sSfVeDvP0nWMmNeWskOpBuBOwgMaz
mSqpxOrpJ2NXGUSCInDaG62uq+IDWIAuJrcd/4t7VPmKRPdxFyUb9I0rNCV1zp0u
4HpWTjVWrn+oMh1YVhOL7pBfDFae8B0Dp/o0K6ffu+GJdJ1SMK93GA1ChoLDFKXx
KXpPsbvLKgVO5mI4tj9k1EfNXcoAz1zaujROrkRaY+w/5xr7MHUZU0de++AU3FW/
oKnYFaynb/TICa5sxkKBonfhV77NQyRjlteOTJn8I1LfS0aZ+llcnI313gFn20/+
dTSo9Eh8FacihOqKZOu9zO3QEo0jpRznZnzWHDtkupePloAIAj90+ZhVK2dNvTS0
rlXSAQ8O/9mXj20xNMsu0zweebZBTjUoKfkDNz9FAV71xo3YcNyfXLofV8Ta1qoi
Z4p+fTTNV7jzBlJ8jJkqEdBPZX2+nhuPaBJrV5nN2XaNrsSQtXRBaNrIvuX5ryiD
tFjgpoz5YKZzmYl8eyeO8DduHPSpeesLQGMPVoplKL1qN0NXBkG41p+wKIn0IbsL
gWJs2vUP1QOBsVwDRYrOoV/r7a9f7sGWF1TBzksgIsgeVkDWabHVnh3GM2Jiu19X
uf+XCu043WwI5/wMFphaCZWcpengelD2aTKpP4M9FYVsKmevTa++O27/BsfDqpGw
S0L2lGe2ElngSrINwMqIhRNjY5SMqXfNCuMmaXEfFH41Yxx9NbMC3d2RRyyp/rwM
IHK3jD7B2EZNy6z1CkTf8y2gbNNiZA6yoN4UdGTFbDcelrs2EyYD86W2MjhOca9Q
/h0PLvFA+gGiSgEYR4JrtvC9bkWO8e0djVNruhjEdIPpjLn4N9w09v6UfiGRTXBT
qe1+ngemCUqIpBBChEFWvzVQq3ZEyUla/Htte9smc/N4w01f7d/gIoCLfPVky88h
tKkwedNiPDApV1qhcPrW9YqLvrTZWZhoRRzGR4Y8gXP0um+YTXlGj99qRS4AiKGy
06dZr52btWT9P73vdg/gUuMVxj6IbA4qj7X0Po4HJYkQzgP4Y6fBP+BnwzAfPoBi
94BO+RjAjw8DM0ZzIm2QvBe9c9h7HtLMXZbBGdlYXUbS/FThauK2zVHVDhybd1pA
m1cPJP4ZfBvbrTrcMupmnIx/bPNnrqjK9qGae4OWQLTTqdMDmB7scuiGi/1p3yi1
iXCVsJUo2SnUHZ0Ammq4vdDf+hvZfowpRANRnuAB/7HzBcXcySMILV80cXmJ4gIT
TXBZOctmYlvvAcFXdOb4QVHJKFb6re6HqIWPMHYpYUzf0LzRcbOFIAVQ4e4nYcbM
P7i1LJSMHYGKn+KSM98BwudaXQ4krZb6NeW8QIJAdijRSEFzi6XHc3cPnqFeZP81
hcfEx5Hk0R1wo4yEvJptyMRKaldHnvuKOSfZzHbtB0p7vm2yZq9qNqHVZxqcZOJr
d08Sb4sDYyi1pmaYj5Tm0i4tIaR7uWqyEA9m9DomV2A1+DjM3hEvcC7UcY5KEp6G
8/dVziSkMAwCbhgZ7BGU7+VjLj+OBIQWVkCfjKAlyhdD6hb717ZLK5n56lPPH1dS
G2Fz/L7yF5aY/5xqhe7XL3Pgfx8UafRD3qKNEZot+SxCUpXzLq2u9xF3UelBtxzk
76+NVUxlsD5DPEjrJF00DndZGIop3T04wOETWSPG4oNmHeofSqYlrqAfULk3w+Kr
saIVNpRM2wYgCliIbJ5wkuCVwc66pEKjtcRVNv3AUEZR44mIg4M3H8wpA6OvduF2
LBu6PhO0r4AMrBK6diEQ2NVINTODS2NF45jVTpYqrbB7cJLfKzMwdzuWB9sT548S
jh9WUnoM4KEZ17S3HH/rWdc2VPIsAaV2/rLaZ5u09i42lpDGirj+S+zBvk8GuGUS
viU4Mrd+JwK/I1ejPq2M1D16keItmfNMpO/m41OvKXKrZfm4WK+jLxfSCdKwfWpP
WEjN/6TG/Ld48C/NVnhsaIAMgPQTnBNcxWHICtqxWcx8ZFKg6drnHbJ7uZR0UCBL
insLktRTbvL32z0KGOqV5Aa3F3iZQ3LdAZTIYy7Tq3U79TzHn9v3cRSeZZqiaveP
6hExyqqsk15MuvZPStveoI4t9ThmnIdQHtI1sy49sgffVDuAkJvcQu39evAywmWd
xLpvI6KeHcjgTn973pjdnQKWW96gZFEVjbLnRn35RP82J+YBYbRA41BoIqURCf1g
Desh+SzaHmEzm997myLxYEZRNZ5Jg/udOC/g7MDeWSmIgvnrGLKsAGwa6gVAxr+5
NA5uefZLH8cqjvXMoXTNeFyW7qdMpgitC4aQWMooDoTCUdKmH+JZGZVq53cLP81f
AgJbrNUfxzPHvcazZxAKYj9lbSiBjJ0A/fxer9DKJxu83fMvYhZ5xwDsONtVpk+q
/rfcrxI6QLN+tFoyy4Yij3Z9dNQCAqZy1WHt3yHuPPTV6NLW4hencXuqJgkzbCCv
dx90MQMhUMUVVwO6qoztdC1TYfcheEByzwFbgDgfPMhVTgiEG1iPQvmofeO1mjZW
U5F5P1JNCALk32wrEOrhnC9m2nf9odMj+5pvuR9jHalwBo8NQoVbPotKx1hk3RVC
5MIZraS8IhZ40uvtSC/iZtzzQDs+s4PUFwlI6PN/BoNPA37o2v9G61DB+GqV/Ves
AJ7ViyMhFWFDKJEt1EBxzmD/p2O1XWgjwpzI7jH2hJIWjwAhtFzlRdKaGtz2PqWe
2/2B3rZh+ygEnB495svzAeXldQscdiMRbdwgeVUOao6PeNnnRfSRPfGiNig+ONLT
ZGI13wAm46hB+yHhVq7+6u/fevxo/Y7nXxhETfslgDWKLVRDF9S6TFciFg55xW4w
2Zni9asM5qmYRDJWftCSPWYFJP8bv+HHrFFJX+YQfuPNJkfjz9/6UXabG4sYMoz9
RnJkzk+oS3+DJ38+e/BTVZe1NFcaBQXB3OWMK9rquqywq8zjwvODJvpHOQMa6V/P
Nbes0+Ez15KX9WS8Tm8PMSM/5b6Y+FwbQqsWuht9Jkh0YjLBFUnwTcUcJfSn2chM
8p0+xxmyugZsjfB+m/zixuIjz33odn16T8awl7qVnhBobzVBNwwO9REanc2x/062
4NX2GI9w3cz/TrK42tdPd6R3XnYM+Mz8QY3W4yUWPuD240Klni76zyCl5qXAj6Ta
RWnSblhPHpXzit7P/6UH9AFg7XJ2crVQtp7pQH+Jg+6QcsfFMeDMya0lE1tuQadb
M+sQG7mJcb4lag0+Ii89vRZTMNT+O0GN3byxSei//69y/d1Ib4XS5L0hnn2wjtcU
iT3H3NfQZF12RKBZ0E4ILcDW06bWZ4YMPQoIuHPLadELNjubEO+Ee6/9MvD5+Ncn
jxlrT8xFoPujhSWfNOkzUTBDOOa/SMj7cC9U9mFcth2hFJ0VNc3Q6G90EVJyu4DN
0YWel37ja2qjQqy0k6bE4rKO8uBulp60zsSx5v9LB/RJ0CKm64oywVRO5NxqPTd/
qoKzXtfpO75qeosdAmSuO27EB6uDpBoXEMReBeFBEB8+NAy8H1ZMr4ggtwKuxukf
sphDeyPm8nzaLUSlUULt9z60s8y7JJUDvwtMqDryTlzasJQ9sAJ1IrXZYOLmIk3e
UNDiAp4UrUF1rWgdQp61CUYS659Ff7Xk/2ct/WmyaGyyirVdpSRSgkAApgffQCEl
q1oMCvcawSHJZQ//xR1T4nWunGstffj+JaoJEu3gWpW1ReOfGpmmRJqkgE5nbynr
vx0EsTqinIKNMzPGkMTCraTF08vjs2e9hhcJ3yZZ5oaLq295bzu3fN/q2BX+odDs
Jgb+wv+pAZDXbuyEckwe+AWuNBmzpD1I8NOetTo9+FDel0lJ3oH/E3J/jFHrfhvc
YEpnhljlJ4TfAqD59ss/NYkPFgIz4SVHTSaNZ62OUkkoBdPqGru6Dy4DfK6b0lam
HujUXQJnpDQkifoebK3JGn7r8u6IiFKwFswL4s4tiqq2ShSF5aSqt0cJnoAhoAg0
8TvbKsoLve3EtZHzQm9cmjWjKLTTmpPZCmM2w1fhx0oyDfJVj7vQLZgROlijJ6/f
9fgzVa7+g+HxcV5O2JZyL6IdnCaQUW3fQJMWjlJwJ0dAsSAV7KzMQgy5+yDw625D
qTJ52hIXURIvf0G97uSZZ/Cy55foymg1jMJFSMmdUn0GRna+s4/AAbFVnS8QLlyH
C/6zWL6eShBk0QHLpBVC0xymqFmuJr6fAyzSBrLsbE+4TwUbLgOIkLJZYNnAYjOm
OnNzcQPG2SFeFUFHwIPvkhXHb5SrJJ3bL2LazTdHwsz1S9FuGTKMb1jtlPVtaRFA
aHjAHztl+M5qi7MqL5MmM5EbvoqNN/nQLYjtsiRhTdHRsoZhnQ+vQuEUpgJ2C+DL
uwnAn9mKlhm1aWQV2GvVtlljXworGl0vwALIH10irV5LkgvRbyOI4JuU85MmB1QZ
g8oiP43hLSZ30tDCSQ9D14ZLDSRtNnXmcGjp2KDyxllQjYgfTZKK4YR6Peu49hdr
sKxHWYgbYxIaYX81WEBi+DxiW7qK2DFgPiHxcRjp8J6inzoDuXRAQCB/o5aOyAdt
s2dRqAUFSfo1oWo8wiUu+wqwOq3k7EX1sIU6QiFQUfATgYIBfKv0wkUmt+jHBlQz
2gbb18MHQKkdHVJF9qob1nP2Qng2oFLUI1/6CVwwPgXALejCiWHoTH4uusXL/7gq
pvhp42efioTWZGlHStCpbVOTjcPl5mM9iqQxpsVuzoq58J4kQfoD7r6tzgO9DIE5
B7Exwz+65oTbCGMS3WdLK2OR6HhYao15q89SozDXLFDCtkitt0GPQUDpcyn6V0Og
RKHoNVH+BxsuO+05iMdm07wKyU2C/G5Z/ovn9i5FZzp3rPWt9KwwWXSAC3j28vh4
g8+iCtsULsaMbNDF5j0OG7CtC7n4CWg6uunOpq34CY33kpJOMl+aJeN6Vo2m3H20
wWAFkwOKNMbK3rFy0hcjcsARP+RrxTCMLm8L2vcLDMuKGJ1yjLkw4hGQTVyCrwO4
gK8lUmpW/0gBJ868W8NtkugBH0SPENcai+9UA5xvyBvq3UNgYRrrjS0XwjXlaaZS
Mna4HJOpOF9Bn6NdeE2dhmCoPutxHk8rKPFVXkX7b60eEhaajsIDRCgK4GbULy3+
Vpn80Lg8a/dj5UOKbos9ZW9DBYrIfwQL9E2LqirlmI2N/Y/NKgG+cpI/36sDdlE7
KOPl+xIz6OaTTPRltWth8oyDTkJWWSYOvP8TsmLAoE9LIQPeGM/yaxEhQ2BoDikT
1NpXREVzJsXyU0oGchNxuxSYoCY4NDlXDtl+X2RN8PlVztgAN7nrxKRBL6n5mMT0
g3cyXyPk7BFne5rZEYkcJeTefyDPZJbDcFgGzKaAUmGCruoEQEw/JkFqOVKD8jAz
/y3F0bNoqrZv8mcRneL18uu96GHcob00deE6u9zAzXxPJtAnq+L3j1bTvxPDOX0B
cGyeGNQW735E73nHh+QXq3tQ9abem73WoWefMV/fZ+oMKYa2g9VXL5cBDao0f3RX
CdFE5MEOWBycCM+abeC8uxXnt0B3LUQDBWIozzM/U0wo3v3+n1cEikug/MRrMUTj
kXeHz/bTSv/ROHNmJen6ce6QkDTEv5KbfZx5tQAPJvHzdRwCp8wl5ihjZLnT0di6
kFuJIDzVkbo9yKNPTCLEroJN5YR5DzPYu1ATH2+a8Z/pl7b+emT4gXQl81cR2/tA
aRy/u765H5sfYksDTXYHdQRbcsu5Bz7yHwWaB/mRzC/0OVWzJ2fGOWUMxm75p1Ti
srFqkIzfw4+izavKQjNVl8MzNGXs6p7drDeIkOXmZTm49DfLNAklcE0L+7szfE9p
p1BBnQmhVX9oHNQuzAS1ZtMArd+RCjfPOY2Ki4JZVsQGLEsUOQphdj3FWt4TSvFS
RJy4QJQXCQ6fLY5MTlRRDMUaOrV18ahDDO1bLZI09R9JnAQGX79VEm4wlJEU4OXm
YQCcKtJwoIC7RXbqgVLqTRbZ8aUajxTOoFlzKqL3ZrVYpIB0t5Zl6PKxMzB6w6/9
BhZ0cR9YgQBgoGnT6gNZJ/5e5/F3s2Uba+SZIi73UPQiIEsNeY8Ssy22iczCEs8e
AjbAV13bgBjlYIzDKb7bxz66u5DZ4H3fwHwmrRgXREZ2FLCPnyhgUHNbPURrwq1S
Mz+ITtHnPYmIV1y9C0rAV1bGEp0WGvw6aUbP4hwS7bRskdSv7ZJCGH6g2uYlliok
8M8fkchPuTr75HZWGhsDVpL9acRN12KOE0yhkXpJZTByoneox6EpTew4hhdAurKC
aOvvPL5M1t1N2U/WkhUWLLpqZYgldYvbOUuE+kVP6AGDOX4hq+3EzRtBFQgjYT1T
cPYO9vU8hwJNU/lY+c4wSqy80aavy/eYKnj1pz26JQj9bQw0iL1k5Y+w63nwqtMk
jeUBuhUVaMKye/yw9bOHbDsyEileBfKEbiYMzCwhAg5xbhuT+dTvQ3gVP6mmMdEM
0L9ZjVQAgnb93E2ld9v4JPRQ3zsnBe5iv8HgNBkiHh4b1FycYAnNfnFozA1tX2bv
g28atQjT73+SAxTQ3eo+OPVy/exqTCK2BNKLoE4UU1Igu0Wagix0Lnqrlx2fk5r5
nKOiJv4zD6aWsdXP+Sjc9Jdxa5o4pihTaIJnMBCH589RyW61SXr/h1DVze29RJr6
FdRuqU0oM7olFczt2otwCCF1ndmI5ekMpNhz+0vOcLqQWygEfPud52Fndbs1+rIG
8dwLs//beVvVqdKGXKNryk1rqfUDak/R36qMLrhx54CQ7xncoJbiGlMtnKDVwIjx
VFKnWNgmc5clL1NDdmauRK94CXmAQzFg2Zkrgd7rNDZ4q3RJFUEcnQgCutQqjNBH
3JMAG289ePMlM03I39iFrXaj62mjQNkjCDF9Jy+TwlA6gzOwFEsWyLBjekOED5u3
zIUBzPT/9a6hTM/M/GJo48Zr9be0GD5uoI7xJqdM7/xAN7oSlSD4fZjSQTVeN2hI
EfxbrsGV8qD9Xyb/VvBqHxKaobmQaGkUE0LBvla0lgJbi+4rzHrDK91i4RHBopky
wMVe7fq6EB4PvrY8fHYneHYtuQ66ZvVhtgVKOvzt+px+v3LUMGSmivYMyIr93YU6
ZPEjtopnfwlI6/JupsOvhIM0pypai4b5PXvdCoIhhbnqixri6dwL5JQySc3XFf8C
iZJWl3a3NJw2GMpqAzqk4BWCiDDnGamwkfRQkof7QzZ347DwvzEhkkztm5cXq/Lb
G02MjtIlgwbyB9S2hsUx++0zGwypPZYyEOh7Ot+NEE3kmTAzG540adCpWpThvoZX
IPUV4VzcCFie++7gQcEZmFqPebgsNgUm03sRE9oT8fJJ2ZoUIsUyS2QAABCTDrgA
JRtG45SzCjpduyFdnzkaHXYBI/3gEagd5HrHCaxIIUfXJl0F5zN+syVMgIDaR+Oa
mgarbJVmLBpkyAeK+DNJ1PJkOCHaMB7q9R9/o/sG6Tg1GoaXY9hLZP0U58hJFOAz
7IySMNnH3i3Q/k+7SeMCvKgmHG5FP5wwsg4MTAaD8krGkPJdwN0HlMOLqPFALhoe
UXylDvsklpYuCxHmIeTxPfcXnXCHn2Caj5tOaT4M6ceMi9fxWnQKDloZOtvFcX8i
BxFvin+JuW3UjdkI9RyZ5V0LHNFAkUYj/1XCxIeMAorjM+kjPFN/AVuqSiazxZnA
bhEn8nqCxT0Buh1qzVeqV9vP8aZXuICV4DFaxNf+d/m6MripxHASUuiJ7L0fQTJw
tDPHlxneEiFrllhBb/PFg9gS9tTdlCTWy8gNU/6DbPjlAv2XUh5vi9TJgXP8SVvM
ddPv17eictTfTLaA7c+OGwg+rGH4KvHYOCbfRJT9mNnTNJlVyZw6fKthSRViaz9B
t3eoCxpOI8PrYCw3kjoWmpKX0WKA+iCUYotShvKIeLQS6VDy5xZOG9FF+P5OHtNE
22g/sdG7+npDH/790IeLw94kOrBJy/EHniD/t/0EOiIf4hhZcPXF+GEs/dOneNek
BD+tAbTqx1kQjZTMTvXpc6Yc/biKHnybbm937l5rI06kG2g+8HTfPP6PLCpqVwtD
sG0EJ7yOr268wH63PECznplauEdMbLjnTu0HxSEoYB2q5Dll8/mjKVHcL41Abo76
WGqod8e3vfUzFnLyEy3NsjDnxvCNQyGHNxSMtLl72chhxptzVYERf9wBxztQhoo5
YDJd7mJLV4rRXBEZylbj3zAt8Eioyx1jbGcxpaDfPW1gsbDytmFE7E6XlziGauez
9kfrk/PE6KkWbPnMBeYpxeqQZjGLRND2qlpOkZce3P3z2K360C76pjNX/QqWxIlO
cCuZdOH8byRm9LTaHLibtPE+1TbHxZpojJ3BMTEAGJb35Tyd+eH3PtuBqmtzMifY
GpiSWZ+oE/v4gW4La9E161xDtvLApoHyzjR+dYlrePSQBmWQHM9g7GPu3uZ8xRmv
WgodkVUP5wrVv2gbJxRbtOFmO9APRe8pOkXBw5jLEX3h9j8x5Fzepv6UzUIIH+eM
KI8+cKgXt7ec95z9Nnn4eeG+Ye57lviC/LSywUCKLANjayTNAOq3upygHf+lhp0/
vUZsnr0k8JJy+iCFSLfhpr0LBuV9n0eQHLt9hjhEL9v+sm7J+ZrSwTIoEcPnAdPx
I/Z+3aKLLdQMUeHAdXVkVhXBauxwpm0yPca919vdwvwyPJ2Q54A4POb5Rds/3hJ0
Lhq/6W+MOSpEMuw8slB2CCxq6BLMjup8HLAp6M+5rxwNfbGG1GYZuCNfuLLHZ0CJ
tkRRo/ngXtdkijX8gXoJ5tp6HmmoJW+lNe12snoNMacbZx5wKchmTSAQBAFcRdtI
QwBuoZCxdi5v9Ksmm21XqEqbymhfCslqDoUmyNQhCrRaS+T1IjnGURn3fI/K0RH5
2MEYsH5T+bMGSQWxuv2qc++1H5Qfq3k1p7sUETvCCtmBelysbFFpcHD5k+pRd5zJ
Adb02HS++cDQQIrgB6YLmmn0pan0kG++zfAdObPCaod6fjtuFhOsMn82R85AOW/a
aEQtutI1V41OpL51RAdjYrGtbj90JhoELnvD1rD+mpf2n/sarxMsd10whABj/CLw
BK5sChxwns4AtzKLEE6nMaEixBsAbtQt+ZzcjtPenPAZDHUruw8dh2zP3hrxbQrE
kzjoMfddXFY4rf5jkiuwQIei21ndEd3h3Ch1w4uos7WyE/Sewm0E8aEyvL03CZLU
YVIXkAX1SNZeZq/x8NcyqJ6RuZ6PZXyIc3nkiYO2Bp3K0UM4KP6xZ4lI1lIpT2QE
jE24rusLI6oYW56hsUxyxgZkVBMZW/OkiOZeU+/j4Cz2t47Df9WgSTOCG4z187+t
7RIgWeyeLIu6lhBSZ2zVZaTHZY+bIyrEfW21svGJAQYWGke2FL7P6x0TOy7j0Ke9
5G4CEoMn7qXny2Cpfb74qsN9ffyl5SwcY+zkqZ05/sstnYr69rFPSJ0ZJkr9BD/O
tg83A8ussc5RRRyazv4wOYLgY6/DS2vRCee5JGxXf3f+EsuBANxSwUvdDx+418+D
oleksG8ymKcyUiEi2PUjywgPVMnHfWyPrRrlVrN1c9cMuMVF+EVNUL8twcMbFLeg
hnKwf29uP8evLSDlnR3LsidrhHHH9p1dNhIlguF9D/7jaLD4JHrR85eQ6OKFjwtD
9PPQ+FfiTXnbvp93U7NPUEvM+D32aXkjPjXTinsonyV2Cr5690XsV74rRZH6/o5Q
qcsN7LMz/c52bRMlq35/K9YpiCOFEWhhatC+wVBF9xJnj8x1N6A2NWowtqPcIn3U
4UIp7lgt3ilOrQdVjkBSuXHCZvbzuxMtaW5JmPaX0NbNmSIY4vH3rtbemr0Dnpsl
1+tS001byvt0ThiJk5seScYBxZhdwWh5cu2wE3iIM2H3QKbqyVyf4bbgTe6MIcA9
Dy1mGzHPShd2oITg80AT9W5baFN+RFS1B+6aeo0iQEjrDEB0cJCPsI31WzNHu+ZU
hYlDyJweRifDqoMJFnOxA4ATsB7soy+TlTmfbwbIKfjgoFtS9o6go78uHwSA+srL
semxqW0Nh+11QYo9y6+wu1KzG0ZX/sYVIMUpSAcXH48YQgGAijsQ3pdJCcE15Axf
aHu4vZ+sWm6034U9rm6ot60bicxULv6Cn7PEtahtNlW7pyHrIFATTDJ3GXRnVLUH
IhD4RYZk2tFFDViFT4KKGhEm9c7EtjVnzWe4/JkjWRtDZ1Mo+VtoczARWfGoXg7N
leDRnzXIU/MA8+pf5HE5tPjKkvLZpCZzOVhxk3SnS03ux5L4SVScRP6LmyXp6yZT
najdFi12DqWD3u9ChRjavDQKUPx4ccFerpVd+gTvy5mn42Vw+R7fZybktuDwJ1xx
MAdmU41Q3W7rNFxzUvFf7NUtOW2N2dP0uS7ZjPxoyU2gxowCJjxURb7+znQBDVg+
Wr+PmnXBZ4gMuYjKFMqP5PtcPVJRlt4gvxYGSv7bxxLPLu3EeEB3xU6Bkfn01jrk
lC86QZbrN5McNIY4AX9l5AQ/GdleUhylmv8qMkc49DCoeQUmKceyyzzoIalrWtOi
TyxeQcS8TSR/5DsknT8okoW13hsDSBfzauTxNz8f1frj4kgeCkAFAI4gG9cnu/cN
pud8yGIem7sks/C19z4mHCYN+4brfcGJgs6C4R9fEdveq5QxVqPKU0SIh5/WZQPK
N8NXMQvj4TuZ4RQldw8W1BMQ9TppL0vfWoIw48cglzffYd1lCuOmgGJ84GMS5Uxz
dU3jcnRb5VP0B5SararX/gxM8ZuQdjV/yIVCRmOL505gqNfHVU597rCNdhwyYqW6
INNyzOitw/wstlJWvDu0/g5LnJlgLvO3ufw8vUTpkvIQ8/cmYnaI22RIdW5R40/o
gHKK6lY2TbWipZ5uawqNdH1DiXOE+MHFRQCHzYbBJxLkEqYlsKc6KLCR6PH4BAyz
W3G74pdcDz80wTjUH/mSg0zQ/Rf2d/4y/99RoTktfXOzwcEZbEGcVRvEiVeFBL/8
dznw3pZnvg/njGXIf8Cwig2zlQDv+lHb+QGcEfk2jt3n+J2o7b30NGvLdh/VXz1p
cAQ3AGxiy6ca1lWJ4YFPBNreudiOOoJjsBnCEvw170vOIr0JkDqgCoMp8nEI8dvV
booDVXWD3ndNf6NaUNtVib0BIQ/n34HY0waP9KetuV8OWOFzSKulaJ27UqVEBFaD
dzq3uhsSM1tjL5iGqp4GXWj6Ak2Ux1B+qRXoRYUSDdZqBZuNastCDWgObxQvBYnb
/xf0AjviVa0lFUxUkfptuVR0glm7KV9q7VPSmzytKKPA9zkxyI94sqzX2Ya/9isF
t2FL8bIo/U9FMfZqGPn5qwcZ6goop+oJditZqKw03iN7wPTRXwOf8L2LY4AzfkWc
H4rzNVtNQM6LjzMVs0JgWcifiVUjTS+9HiU4okng0O/WUMWiNzr+v3zZO7+RL6vc
czitsSPAl7m7DiU2wFivUYHarFtfRSd8zTzFbMrqSTQ7Q+c7D9kYw31fPuAQUQNp
Mp0T9pnqnv5mnmnxyv/skW6kPH05M0Lbu4i7qXLsQoe7rHV8UKudk2fTIrst4PaZ
eg0bhxiqPjb8mfOp/v6jy5BUWbiSbhBlDgk7mDPPJeglHfvLW0+zhL2UtycluyWe
YSK/h2x1VKamiDpBSt356YwaKFpQXFNkv4Vh/66MhwvxvQow99Py6abe9wgVZ3UV
h46TIJdcATm/dGytbS3n03M1XjwmYda4tE87QiUdJKQFKr4oY5wgJh/yQNoiva7P
7u4ggNeojt/UCdrTEJOAoTKSgJ6exOzTfrkSbLOzWoGW8vV4tvyadCvAo7fxOyWE
R2l6SyT9gAkijs7e7y9x5BHRrfHpde7swd0RsG4FrLvihvzGkUPASKEk6CfWz8tV
xRaq4xsXI0zh0+dpiiktYwmxqMilfeFC0Fr+QUSIuPw82dYymJAKrVztz9RmMPAm
CoQ/AHAk55nDsCQbo1w3SY37Ibd0csUnRGITkpUb/xFc+Z2XQfvIyA1qDTS8lH8Q
uzhsKP1wrqSAQ+7p70kPogz54U7CnGJ9M0MPSaqK/nIJTnXQCAL4EzaLvuvz+WtU
4ncNujNJEuOZ2lU8KcBBLdkX44yMx/Cn09tnp4syVDrkx3cjt8HUo9T22Zy1yUSg
/g602EihkqH2MB+YN/Jz23OM4z5aP8a+FdVL2cllCi/gKTYhXYQ3OYxl63HvCvWB
1x+GnWYfSk3Y/189fV9k3uqWE35x4hTlmo/GD4105ZqgLaHlZ0HleLeeFNCIz/D1
pfQ4cfzXwXZCambTG8yCwetAh7daWmsHhJ993UbMz29cx0Nvz04AzuEm+tJUqoUE
f++LpMTkyISQiwVVZfxKCatAMf9OYvF4DLi1Xk1dr8Rn+bxHJ3Occwt5+wXCEOih
TUERUuar0a2dh1494Fzz9JaLtPXTd8z2QuWSIqo8hw4bem6VFDwdsIRADuOUL+z/
repoOadOULVmsXf9Wdr0XdvGMCcBfPI/E780Ql9A2q9kpLJYocVqzcfdhU1ET8D+
Xjd9L3pxD+H+pwtJ4w0mDZR49NIT7aDPcgflnLnX3pWyFS8TgQ2k+vqfH3xSTRkw
01lYy7CKmBULgoHpLsP0G+LmHOcexUzsPKKF3apVX31uSJqT/JndCcZeRVX0QNqn
lE2msv2Jp/PrOCLAtIHTWJKcEAlusiBR+56gf9zgSgbuDIu4LmxYo8LMLy/9jrl+
vtwsp+eKZE5aTWbOWX9MBZddgKqNublf0vU4Pn7++dtmsmlDnt0oTt1GYoiN/Mqy
Xx666h3TgGIAM3kHgvIEKkcLSG3vpoaQ6EVuZWdgSbBpkMikgmNYt42qD6+ErQ0v
02NGENGFahwbXe8l747K2ZJRZTJC/R3MRq3tE3F8YyW2MyrRxLvH8eprBfCf5TGh
FwKTfuo29DialSp8NN5pJtSwj9RP0AL0Oeyydu5qH0XFwwArizZUDXu9PgUqQDOY
fq7Q18IpCUTJRYxIaBRzW5USvI1lNYXCDYUGpduRujDILrLvmrr5dj7sH6A01hdJ
X5aGNSVPez/9j6yNoCd8WSd1b4Dm2/BqP5igXk5VXocCaDa3rLrfA33d27OVJhsa
pmID/TNqc2ffEdrUHIyCrMwhU/uUVQ5dRTVbxk4sx5M2okSn+THdzpmPovxkIxUo
STJMFKNrA881/Cfc37KrhuxzMvNcqh4903AdkgHSgkIlo3Xb4UQprtBRyfRSgG7S
vTE+t291J5EZXGEi+0F7WmU6m+jsbj5Ge6iYbQvhmbIgPFxLRFbk8eZsE+76Z02j
TH4hTIc0YEj6/+mO1ajo3n/QBwXTDa2jW2bvTpiGgIyqCVqkr9rc9xAQWYGdlxsc
yhWJrbWkHtA0YTbP5CZttgjQ5vyeiFwzkLjRjJjZCrcsFwFA/u1Cjzo9b80Ku94F
Lmxc4Jea/6ByUEGI4hU0ik/blneHLZD/b1fKuNFglyg6U/Ds+qbMxzJmYiKnKmNq
lBJzpdsFMx10UyTPKN4SRtyEeGcxGpFmxvf15NJLK4BVN5jeFupf1SvqezlOp09Y
5OvybR15+WkfLKCacXgrmRGwFFCr4avdW+iBCUC6NgSkrc9pRk0Y4l6HBScTYavA
+YdQ4feh5grqXLNPkQFHeP1+e+CEPJQ77/z/6B52A4Q02zgxVRQBPEh8Hktm58kz
b6h2qRooxnuz6NJvxSw9n3K+Bog0kgZD68Op6cGRwPJsIuTbxmefv0Q3YTpwpr50
Adh1smcFglmPDSR6b+dpH8CYSl8iCKYR0jmu0QqfNgfKOtgiHLhOcDWzokof2oEM
lh4Xl55/34Lb3qq4TG6IbFJ8jppdzAQ4wtqG8c51XDojbcSq5FWAcuMs+pyFXjfl
tlN6HcWHYz3r6BNdGGdm2ka5npAcvfGzCLSM6dHGuJlMXdkhRUoIU/YLAA4NV5+P
YXMQfHrRW5zpa4N0Bb6M8FESdU5WSYahQHutvUuCqyTXpVIfZNn0T716e/8fFELb
MTXwvWGeHDaFvUbrYD1RCzbza10B0tjko0NTDEc3+XGY0prnF5W3DsuY25Z9qWcR
rgE0IlBPHANPAz0y/j5tnjgm7gS/LG7U1OvWdyfgklEhCmLlU4G3e4DXIU/vflYy
YdnH4qWpmIWFgIvYMEn9cM2/4OJ4fKikBo/F+0/4p/p7rNiB6AAqeI4lWsNG4ou3
nSIbbvRtsb8GhF2X2Pe5nkSJCvOeeqnWW7RFwYNqa72lnWhSwYGFj0YS28+J0BmR
U2I4VfOYZxJbR5ixEHSGjRwoaaOcBP4dONJUTNhY5nZrIqY6BOUvKHlPx1nwWMq/
9sFwa/gFyYZ8MYE/lafazK8dRKYfQSAFL3xNX1/U3tL6AqLngIspuaJBLKjGCuLH
XLhMtY2HRFEFUb5tiyHtdQqvpAE7/c9SdWm7wBr6/MiWJZOBxiAX4wtQryAvges7
Hz37m7gvMwbYWPMCwHelSREr8czcNePJakiCYQqhzvmiwrBVWOwbeQpMnkgZrJQy
nGSJCz0UgOgbb7E7/dx5zL40XWKSraU+nrqj2hZPLN5olv3P9zuk5WIoogrcq/IW
JcA8I7favDFpoILQOKYfVA6QkEvn8PWSA2zqX8nBiXxHG3Wy+ZTnF475FYIigkm4
PdBNlGkQ0jTJq4QqJfQpGwW1XVT3TKjwiGIr2Daen7wmnG5bBQC7NNBkacUdxkmC
CnNJ+ttmg+b47bb40DOUh4vXVXIB0k0ZWbdKyRZTjrKufO7TRAQkjZGeRwBq68BM
u+KoKu+Pjg7AFhf+3pogI0izEVxUFLc0b4E8a52Q70FdB5QS6vGRgenrxf77q3vZ
pbptsF+wjldd04o4bXRFf7W8i3wK9MGFtIKRuoz1IVE9kk5JmtZSNmH4gPoAzvg3
6FxhRHGAaDrD8w6QMROdgwvIh6ElefUAv0exXSLQBw6UMCUiFpLDm2WtI2AbodUY
8+Ur1TTNQx268OnPUB27JCGFmAMC6LyO4Sya28ZzROwpGqt8GvfwER6M4eGP5zGf
E+cQHuqk1nK6nKIM67naG1LwzamG83HtGhP0AycxpLhdW42g/OS1nmMkPR/yFcfy
l/wrc5kauq5Qorw534b61S/EHFJOnesuaVcbwNxJZ6U1jQydZltp+iO/KN/WIXzq
4DcYTnwB0PldeTi3e7uw4fszp4cGNDSYmMvUx4UeD4TThBrzTxGjcXsjFB0w1GTV
pNiE41DcUfgbITf8dfGoWhI7lZ1uepo0XGJbU/mqw8JLQfrVC16j0VTaDS79VlF2
0OjlPmHKeNSFNzGTNpz4P2EQEh0sYb++8LWeiiHSD3FyBkRzyz15lteDKRGSAk1a
//dMHDjXZItcWrk14OCN9UmeGTHv36fj5KYoLBuQTdRhY3Nw3rm1rb3eCBG9ReW/
yEOw028StZ7RidYd3KveWcG0pWBkoxmn970F24RyxMg2CPGRA5t7RVluqyAI7DSI
jZXEL40hw0pV5HF4F+JvAqWURta0aUUl4/42ey0MvEy/JCKFicrOJoU2s73DiiGF
zet/JmkHMPzOxFulsJXpLqmp2WLUMNarsT3Tma9CmnZO1YVslRbOeXe+9CmMzTij
Ok/3kB2s/64pk720rRpv/ePmhloBNvnkHcTAMwruobOcw3qARWTFQlyJ43QLBhSW
SycH4dN4CkOI+nkjKnwU/4f/2u/YMzGqQnrbOjYnU4iBLqBFSwTz7upKAHL8sx1s
a79vZQTiiV/CiRcPPN4o14YNyub/7Vm8YXKneZYmPbtUGWkoC7lsU/uKsUNqsJws
lr+811ckLASEuLR5XEl5ZHDceiUTU3LXxBWUoKpFu+RnTz4p/8oFWaK35LuUpTBn
n6lKh066+QZ/qgwRMjcIqvpkNVxlcbdi/XDF5rZxZ/mwyuCrsH8suMH62MnjlvK3
+i+3YUpPaZIUBlHc9bRhCLbqTmvTjRCOo/yPb2UEWuRuXFiRvrowctuKwTofXEAh
uLS7Q/ePq0+QRR/c7MyLqccrHtcmm5sfyTeZtoDLJLC5hTS6/qneLUUIaQmku13Q
2yV+FP1RAAxyCA/LEj43/kSyuj7hClonumqOIuxrWX/PhNjxxqdcY/4/xtmK88Px
D64Q9utNaLjdMu5dRx9q5eRMRP9gmmF1czL/kl99aJX/LylhIvyr6LllnuZoZzJd
AAR1WZuMTB7clHMhI4xaodJkb2JGw7xgFJbsNedlWEkYyi7H8z4+gLBC2kdLwLr4
AO7KgPOPkaedvvCzUyg1F1dXZp5Dhrtr8DdS25to0YQTgZisAkBCPind/HYM5wQv
iwgWtXq/+MNWwqMJyQXkRq+dCkybhriQ5qjg1zvc3/7X9q1ph7xi518z6+OD6oTn
TMcokY2KK7p3kWUOfypvt47zMrkqhMMaCR0UKq3QSqhlJIOq0tz67S15EAe2wP0T
e1SwDKvNCIpbmng6XAMd1ME2wyKVrC/FeBUy6Vynxbb0Gnyi/ZAIBBG/ki3IZPuB
mV67gi/Kc7JnxveTmRFsqIIu/1nC3aqEP4R5Jh60QYGpbxdruKPkccrrIUZsJG05
gdf2quOLtFaYyAosVwkWlpVQujMgEpg/jcpWeftaMGJ6qOCwgr09KuZyLsJm2s57
dFCxQ5ivaQT0yYW9Oql2DPRuoIblJHcM8L0cpDZ4fDhgtntYZA6qJirm6K51gw0N
a27O7H/DX9uNQLXbk+vR0szSJ4HN0anGTcn1VDkxpGgqJmGndDiYr6egIOK1GE6/
WlBlObVSglX2xbFYOrptFI+m3dQq4kcBFZMJSeB/61xthS6AEiMw2XkWwdXesQN5
wixvYF4vMyg6k7WIqvimWIow1AK/nUSMOTEJxP3T/kSbV2FI/guo8K+eDYgA4+Zo
JPEuS02kYcpDddpzRQL6TG3ZzQzhHew/C2JOHqpMBPUGJPndKoJfejrT2VxUyLEb
TJRdbAA6CukwFQXqLr64qFlnaPbd34QHzmXKvdSzTq8jM2xtmGfBxjmJBaDbp+yl
kUcKZKTYuuZoX5NVIanWnNlCOthZGqYd4flfsdksYOx9OjjDo/on4jha2xdWigXV
vtpwgre4Dm5E95oA4g1+shmkzW5woho001vX2TjN9Go4Xs57PX/96aSLVEDJFcuR
N4F93FvBacaZr9nqNuQoTGyqU7aqzhrMPW8Tfn1LLzv5IIMCt1gmIdLcW1SYFTFO
dkEE0OUGGfRfNpoPHQHbdiCyYv6E01sZ9dLEU5IFwDKMYmNaceImmDCbvHUtJXce
n/gXu3L5weug8lhuMxeoLP3WxPknqgOfUP1PyCkQGyNdcFKNPLjweax6fOuxl4xI
3CeSm+Xjd0tUuPKIdWC1QGDNQjBis7xO0Ge1g511z59h39Jsk/+efYQ4JyNnrtxd
5rWkMUz/9tqpgOFBlWwoe+4J9PyxH+H/1A6704Tmmhgikdn73SzyIBe5gIr3iRcT
gGsHj+igAAujX8N1hg4CxHUk5gWzum8++LAzPa+VYITYagh3StNmmk30onU9NpsC
tZKiIyf8f5yn6UZ2xBrUpDYZZoyzFuAqao3XICwKPuETV2r19HKCN1s+nnKkhxrN
Qqg0XV1WRPas43EYA6QxjMhp55qjoBDNYn+9uImbhschZjyGyj7JMTNETEz63bP5
5u7X1h+DTOlJhbUNq7lkWged01ne0SBh4fmNjBnz3bzDJHZU0/6opbQIz+ikPKCf
04he1MjO80RZ3Y8HfSU3at3LrMh33zo9jnyBwl7Ei4z36WrxnlWFD7vL6QqfT/LI
3Xc+lmiQ1ADyd/5im9OV9Dc1iwYE1xRP93UO2UP5YsvADQRfBob5tUCAAVjaCNj7
c87aCDbRLjWzWEJWO9PG+XzbIwanZmda40de0p/CaQqM6Cq3nIR0xndGJxeU5nhz
AVjFMgRFxtBVYXXzvRUUHLBDif2IOBasdlmVkvZvCVDM565qZfHMtlSbp+GdKcsB
1KN/wvi1vj32x6w5dl6zex04cvqgKV4IRLuKjDH5BoO5GMVSbcVchs8zWdbvDYy/
bG3N+2bmcKwNMbg+hBX3Zfc3etrF+S0XWEH//53ks4uIR0WoKty+gLpjgrDgtL98
DtKj5M7kCQzLvjcub3PSucmv/sFz5YdvT3YMJTCHzhHprGeSfPWxKSlREEfwFg8n
RMYBWgraBHYI4L2PxRll6ZeYcrUMzCtGDZ1fjL/u3hn+CC+gbGIpQyLXorsZKz4p
aHOciTQ8QFWsxywHgrshEQfGT70v1QZC8ifVLOZRqZRrvW0MnOBy/2Zrt17/hqC6
KHY+ZwMVgSnKrwehMvWHd+N3uXvroLMZ2oWsLiEElOByy2pjoCbuBf1n3H7jx2b/
LX/NzBxvMIJi+ZTZ+ab81oIq9g+FAXGZ1GeIz4c88MNFnoO6dMtbeM5aCT3hF1pQ
LC6CNoTHKCED2ymQioj7dFpSW9fWubYkDNZO+pxK1HRPZtqzageK3/0JkNRFEQ17
6l1Nex4R89ZevZO16yDli3p3zZ5H+i6RT6QAXuL//wkIQtIALY2pa2cwhbEheVtv
7VlmZuYDWQcOxdBeaJezY6RYUbwMitFadITsmSE8GreepFTTjGy8DRVh6r6/TM6M
smy/k/H9ITw1BvTbeH5jcDT6CtxFiHUkBVCp0HSGvgqLJI8XiKIL/xIKxK91b330
Teogmpf/OspGXSQH4rB/zlOSOybE0scFOiLg3vekwptXlc+WMD5lNQNb+BB2hcFH
+134CbzGEZwbB2fifET+8SK89w36UA2tcBML/ZPR2nObpkBVKgbaGeXnCnoVF7Aj
NB3jtE7MG3vfWQ4A4hMoC+2dNyCsaW6hcDRlSgoIQx1XyV8XNlMdbVQEnjtUjAMR
VEItTobsAjywuu40psGXsseG5JEkzMb0CLysdfnVGHSMcyRufOXcWhill+/3bE7/
7thz8OZiDKob7VlhPHLLkPNPLcOr1NcEWunfc1El0AULG4MzG33aYvk6gWTSMD+/
E+bYb5LHj8mRJKQ3iE14zhYXL44kOmJbD6Q68jSZr42FqSwznJHLeIzPsI5SvXrn
lsdpj+CFSKfvtYq2aUPNF+JZzRW2A3Ykz6LHx801f3zOGvjFJlUjWHX1ir8w8jZY
fF2mkjcQmEU3BYUz9YK9K8+ROJk79vrXrL72q/6ou54NiNWqJ33m96S0Nsn9WFms
hIkOlqyl//fxrgCYQWJga9fozYXwk9AX9BSX6isjDZXkJv+3yiIxn+ILZ83wjl7f
tsa+j5v/GmPd74O84zbicj8M12fVWn9eilmLrA+w0gzAsyNXFeO2YKvYHietYwj9
EHI9COUN6XVpBKK/u7NIDmuD4cXy09F9i8kJvM6Cq++ThP1hPjyZJQz/OI/X49Lq
piVgCfAiPNj8bAdknZFYd0WfYYtJlg0hRtTvUQoT+oXMstAoZAPD9BEeVpctCemT
suTr8yg+bXGJelh8TOvXdmclogdk/rzi7CZyD/9WmpjKbMPeSqS9xr48i3OR2kiV
0auI9cZUiBTLGKqV/goHRD23WYc1Oyo0EVUdUp18hCEBsSzsTuY3xTpI/IMW4QeZ
eFWww/m2ph8vyskfF6bn3wfop2Lpn4E9VcW8LyULqLWB0DDeJdWx0syEMWoOmwoO
EpDN6iO/z9SHwqD5P69+CokMmgAxtKaqq4hK7tOy8rjY9vXwKLiJ3MpBG7GJ76H1
Ad2/8X23ILf0j+F37azV4nnpdopQYQl25KOx6GHhahBOsuPcDRCEouST89/pqLF4
J06BK5sg26lWPZwJRwpFEqEBbvVmpTKVtyskmAJX1TTWGOmmkgknTI+Uw9uZmqk8
1I/kfyuLuUkGzV3CfzNXrm+TLZsn7brsybz5uBCPaTIIyEG36BgkPz5IUkeHha/R
KbWTFpLK07/94I2cCkB9N3UZ3BMV2CyRERNmTpyfjH7EVunrpRTUENmPeENq1qeM
DESOQKpS65HRNyn2uiJ7ft6GHXUWo3ulEo+EltnwytyByJRAx3LcpsJWYe3Vanfe
RuXj3FLe88bjgtDyYExDn/vXOmofNMrBGCMrehtslA/Gb19J0VoRcU7nEc8D2IEt
7tvjh/5OaZVwiPmn26PvzLeY8S+Zt0MZdBnwUtupZ7R+PSWGDGxO/SkM8HNykNgs
q6ecdTs/G8TfNm78tn4R+2qHB/CQlrtUZA4whcaI43o/1c1nf5KW3VQlSvVdNJ/L
Tew4AOUDQ5uN8dwFXD7pI5ha98WT9F8mu0V+PmgHChjJ5pZ0PtOXn+DteLCJ0sMh
EtyphWCi+6zQeDSIVAfZXzTuMYutd9W55Rs3C1zxypXAPxMYqomH73rRMrhtOmr/
UG/NRCIPMUtlCQcaxNYJUZREduMVtiWjlZHwfX1jTvl27a0L6zT1So1+CCu7ESSF
iAOjRxIOiY2LLv9is7mr7FNoX5AlWrxim3hcLlHQIbkLWOK9ZokpRTLEgIWWwap1
dg2Q1ieepLHrnWuX+n+0HOZ2m/H7gQrei7M5vRBK/89G0cgYxQajCcSl5fdqFs0n
cxbDx3/LA0aE0Mb1d7BAruyRqSr5Op7S7h1UFnUyAsGuhClqRNkKvyy0uFHO021g
J+HAj+qGidygcLY8zboGLLfIP+gsYK6I+NeKQBNSZhUGTh5L2WkbM/0l4YYwwoIX
P04VA8g4UjjQxxFAS6fgkdHFeWQbOxVKGNxt0RWxDxGITPqoonBweV/ny92obTNN
rh0Ov045uE/NcJLv/E7TmQPhjnUD3qju07KTUXtAw5c+UNF3ZCWjLqbx1nlmLQih
xuMYsY3E9hTg1dfq5//bPTXHSs+gaOQxzd9ZId3RcjQ9ZaN3WxFfbHJEhhTy6klS
BXai81cFiYKWWoniS4p2HLGpwEyAq1/qUIO22CXSJoTcEhQHgrdrP7UDc2KewGE3
SU83hmiJTkVMU9uh2+3vWAS/ZPCs07fYIu4yPcgkAYE60xk51dEsApKnJcRSCSCa
21w6l4pzKv+6y2/PQWslPvNOCXLX+TlXe+ao7JImq8a8k803we9beH7oDTLAubk+
4HJiP8sQVBj17KRa7HKX8LFeyLqJGyqM/o4kwzv+pAO0kPISnNXUdq742PBpUSCd
K2C+xppVzecOHtZloXTG6YfbCZh8x05fXWnBq0bNgmeBGkgACdYfER9rItgqZWtX
Zj6GKde9mZ1BWxUUMU0HCHqUFn6bc8h4LrucoW2mRto5tNXVuK6BiJIRJqN7pRX4
3bUs0aVe96D5QSpk3USq+J2o9XW4OpHKyGffg5NnsP2QQSFsQydc98lUrs6KXRku
0AzoC1sVgU8xdwbJHLySIN+IkB0ZQsbWCdTk+Vs7EygcGxZ6vDx6u7+PN9lyRZ1O
VoipB5qGtAgbqs3SkHReAumIa0aJwobLE1JAMqbsLUkoaDhTjUGQlO8F9npf/8VP
z480r8Xx/i/OkIT6FhRDz7o1idZShXB9B47VOqZPN4ApW+IEvnCexzoLhQwGjNVJ
qwhBr7AEM6AqsNsiAXJNxlYglB1L74yIL169/rQuCgcCzUNp65UHmRRbIAf1kyw2
epZNIHYX9LOKx4EYX83ZN+ZXyjo+rPNe+cxDANBXyxmdOkG/oy6quOclhFh3v/Tm
gRTeOw1AzRzG5BwnachhXhws18gmXG5XbmQu7L+zSBFQa+bJoc+3MycxFJFWT/6f
0W3ANJlC3BmN4t0W1ShzEh4EysMtu5fWLulGNOzmAMMFpoxogqNzLxoNr1LB7SSJ
jjgh8akcR2HHZWufczP+SKD5ohyIYhm92suX8R1CDy1SkUNshqrolkowWNC+FUou
PQbbio/jDcPho5gs6Fa+uXGAGMtwKbN8UXsJ06f4qvj3U2ciQA9PuXP0LE/+av3L
d52NLqGVBkmyO2LVYBdoxSBilAM69OsAMAaFJeNhULLo+K62QOsRZdx/HH9T1ZIC
BjUbaDfMj55t/Erk6v/9hPftKPzRVu7kkmmVqmDLEgLMiepbkWC2+iEnLReWsvSt
bjQRixoHBiTpa8A9APy/nAe+WL5nf7UwvBSEvbt6ntoXsapEX41uibCKaOphW3dO
FYyMsttRlnqnoY31sl0we2OE2ClTZVQzFQjvfLMp1rWOWz94KJxNOWutD38kUDBc
A/T42Lh4Rb9mAN5RHeEaCd4WenD6eXF5eFohoaZiTwPb83qCmlzWuZe/DKPK7YLm
emoljMtMUDe5Q660uYpOu96NkH1Qu9fKRNSGHGcIgSGtqP1xzGq9w7TaLumeobyb
/WRaOpZpLrrkVT/4sbYyid+Uocs1wcR5ByPYBI4XmSL0wu2R0YGk5d7tThdXyH+E
bEgfoYgd8cYufuzGO0SmzmjKc7vnlX8JqYPk+NfGehnk/OTdmLCc6WPDQfu/dfrA
dB6lIPNgscSlgxUdA3v4tjvirD0jDslmRFAHO8qSBMdX4hCcu+KjGBMCRB4TKW7u
vXRUgyC3if1Ywc66qjD8UkBgz4f+ZUXayLNctXJDr6LZCA/6HTF2LkPjx0O5jvK/
bu6Mmjx7KJmEyOLYkv0wYKiLpBvA3h1E+kZziQ9fHRoo2gIBZarXJNJRXeMiojJF
FixPh3OvRi5tP7l/t0yEIcv/ykIa0mVO/FnzS/dH5uOd6ON+MWNOQn+t80rond8g
9/XTq74ylJr0mWIfI8IlJIJXhY3rb51m6G9CQM+X20Y8iUPrbMCn1sjPSBYntCCp
alQBVf6i9guxRuIH8v/n1uOAQXgOc08MBFX56/Cy1VaROZAaAOR2UoTqbNVlX3uZ
3Um2bgRPl4glreFhZl/1hnix4waEuG5nCXcSVUt1Vf8YjwYAfrtvEVvOLGx/0rjS
SQGLvLITzJybv+9pTMfWGpV156tgu1jANX9hdAFwBsaDumgxc05J1g9RZygwvUSe
VfvoIq90+NTRa5YVYrwOFbS/FEFwrBoxHA70E2L9VVnLsRwervb4MvbDKfLB+xwH
MlRIHgxFQItchP2dcbu1FinvC3rB2ZEBdAh9i4J3ZCv/bEqwI5wLk05vzFYkYP0Q
/XKDOx11JKUubnl8sQRCvkC8dhT/xxrkG5YONF4uXWWq4d+mfbiW8M3Zc6QHWQz8
AgHWgZdg2MgT+4xZ8xGgz82Y/ccKUh+NpAZ4c7J+906sjQVqR4Q3DvVXs8Ovrc0T
16/90MQHyM1NDdrWXKKl/+5z7NwLkcAx8vRDGMpZSFD4ePPOOxi6LQeq9ge0/c0o
jbMHoK1wpohknexY3TfKYIvPzMYp3Ayoi0ZWqe5xFWnNBD5sVUvc86LdBFGFEanL
ZVsUnuiRg02Gx8CIJ1c10VanPaSJ87h0FN+pXP9YPqINC9jHc7pjvVJK7f6iV3fs
yYHespI4ZeaAAEwYCgk3lk2mPvbCFD55svnpnDNVm+ZkX3LIL/z776b7dvMRz3Et
H1lR328iZ/27eYmeWIF3OK6l/dMbOc9DTNya+7Mi4gmzs6RqbXA+Rtivv4UnAZbT
D+7Dh6LdTzK9qg+NEVUivxRLGjYL5dQbjEB0f201qWlz7f0GueVRIUsRaR7oYHdt
BswbabXyILWj4/Pg5vRS+8BiWL98DdfiQqeiO/JkGywW3Ag8AXycb7bfJTO++Kby
GPo/5t/c5Tj4iQNXNdNdE74k/NX1KHgtDtXHJin71vEJ45Dq8Ey2QSGiS/mMdx3S
BCG6cvVzZu7dfnpt73VgwiZk6rE4AbyeOkD7CuhBDdYeqZHvDrrmI8eBk8zEEk44
U0wHo7oqIKy+gdZLHmdWDVPiPp6psQmty2Dcv2E0s1j5fUAz/9CHCCJjWdaO0XPr
S5xipwdVJFwVAap4t/ilKhQ+10nrkOl7R/S2ABnkhlGBm/YIsFaUjlFZm2eweddJ
X2ge9GaEKl1db2z8UnTV6GtwqGNc+XMyOcIiTG+zUzCPXAn+s1YRENAKwlU6v0o+
xgcnH2RY227oDmlWA0oDeFLt69MXNlea0ur4b1df+um3u9RUK9mr+Cn8I5TDQkqw
esrlGUaHMZj9dWmLEBzkaU5Ipo9fqQ8AA+ZAhYiqAiZ4+hcNc7WErk0NDq1eZiBM
YSQltMJfIpeSQ3neyftLkoWTZ8C4Z1MYsGmBvpxbHciVvfRsClxYr0nEFkGyywhy
s9Odm2LfvKCezeLJzhNVjLunDBGNsulL8sh3fb1G+7c18kt31J3X5g2C6CxkRNyg
wr+/BV0CiuBbs1+AZsDm3KEa/KYAV45bjAqWNcuAVlMQ6F5DR08IJgOTwH/SrkHs
NCegQ3y9431p5j0MpUNZksbZ+/xjNX5Mo7v2DJfV7mM81Ie7ukXslC1rE2ntl1a5
lso1q4mTk+l9Zi63PlC7Do54adDefEqJsrlVI9LkFNfSDm4VK5OrZnC0chFMdb7m
c2qCUBEx1mJxCZU5N/zwj77Z1CQaEoiBKPJhRU7GEXN1GqZjmnExONQv8q83aPZT
wpO9rchbtKyJyrHdPZvL7LSjdFotEKLZUO+ruYmI661NYLAM4aCuks3oaHztm19m
Dz4T5Qg7IOPFZQ0XdOUQ0tdKGbQqdbmmd8nUrTOM+t5AmO9zER17Srzr19tNzZK0
b0MT+28suAyGP4QzEHqowTor1Hg8iPFo6lPzC0R6hNQR4nYIzbYUnHIoy1D3mtUn
dm4eS+RDiN0kWbmDmrWdH4jPMxI7UdvkNpTVJU9mvIeZdK523wHQyvtv9q1+OT//
Vs5bugQOUE5QqhmwUYUKk5SuiKPm6qRSncBIEbzqhZ3ZYjhLuszWeMlpRHa4elZA
yUw9Rtkfcd28BrhAKn2u72kt/a11dsH63rd9Fgag3Z6bKu/8eBNMlsyijqLQMtzZ
tNMhHgw//SQcZAiGsFw67IxFmjlTVzWvkrOmeWM7SlrAZhdrh1Qqb9gZeojLp83P
A3IE8nxlG3gVpuRhIVp1xNq+qVMkWrraWYYz4oE8uKGDZSZtXjLZTED3dHBa1nSi
vGvRkB7z7aHbfnNcM2GO5E6Gfy91bh3UwkO37bXKnRtsGd/GQmyV6qsBI6iR0M6M
UlNUK0oZJuLvH122oUbZEfxhStSfWOsWHQnkGhLdNGMRUa7PNRk56guEj+q26mbg
eIWEVqkI1mPAZB7lOVyp/jeM+qhS8B1CV4AVaYtgjN+0gNzaiqr/KPSWfXgKPT/B
p9wQF2twvMGvFSWD6CcJYIxpRBqiOlaQuV8WtMHdjfcZemEaPpshe798uYfNn5oG
nryxs/wHAe/Xo5YzWE8zLHD/FHtHjOItbDnGarnQrgbvXVFO+M36TwKLlskJt9hw
W+6cQJsUBBP23KPNbiAapQDExFxgnfR1lp8y5xkuNl0MY3OGfEUAngWFLwl+FwKX
Cb6jBV//ZXNc4LmjcjK3Xq5ndRaYPfsbFLxdPyZMPPrTihTjLG7FOUYCiYy2Oa5s
GIVV9AxDvpQoQoXT+gagGnHX6q28ZRnLO8o/o76U7LpikRDyIar5IQjmqeviezXp
AbGyUcZKv14X127Pntqjd1gZvLCD5N6Hm7qAJ3hEvAqR29Tigg9+iuh0Hw/oquW4
12MLZS1WHIzaqgAW2laCwZc88VLkswqkxoqVEPijV14mi6lK0wc9oTaLgpykO1CF
yiITB/ekfl9MYBf6Q2GBd8WasqzVo6p9BLKNlwoDNK8R0DRiQOm9tTFfcVa4/PUf
kFlsM5pqrBiXk6CviVMYEwYV/lU/x0p5NpZ1AX7jxkd/NTiavyVfdHMh+9Rs4eVX
ySaBzExxvWiPJWqMZb80jP0puh2V7q0qeFIxn/a3q1yaSoZ4ZrRbDlSmZwo81ByN
Gg8KLhTCmLEIwfMEi2X6Meshh+cWsxfLI1o2yvf4OzLIndSGJLVdV+Y9fZy8EdRK
YuSRORdSDM7oCJH5XEeNq36mE2XvbNXdXvRe7eUv+Cg3ONnNjnT1PO0AtY/qpn84
ekIcvYy0ymejB71jdstWB7wkYm4e4L/tdrxTWQwbIsmqZly8b9H+g7tmLFVIIdyt
WN3m22YQbqzihVhPdlPkUYR1gLwTAqztsiP2iCQ45fgfQJu7JpZ3at2yPfZqWrSw
5QGVEoVDTEBdXj+nTq6GFvpE3M0sqjAlvtRkFtSatyBhRm/CMCwD3MHbL8M5V1T5
x7HVb9C7Cv1mVMLqknLMBH2WYlWi2AWReb9R6ER9BOjrO7op3NccVbqVhp4JpI7+
yHKIGTbZ2sZJRVcbptwJBaAiuVUTGKbUSA6K0CQrOfzthmTb9DmZ2E/H/JaRACKD
px/kZCZi9cv41lLOhEW+o6db7BZMu+O0CCTjrCqHh/xsnlVMPHzJn69THO1PoJYg
e9dYA7DDkY2KiBGlMONoRCl+v2TdtsTGGLIoobFHe1topjuiVzgLbnHbVqLd/mxw
sszFKb1DePvM8P7xFFKXL+Uzrr9r6+sd2atLpeIpiGwPyVHSB7ITTmZ5VRwDGp08
z9SZZStrfvcNJhVst5zjT9IQhQsoB+C/19aW8mnBQ8lLXQ1pBFrJ3BXRvUcmMNGB
AVh9WmFomdAksA4g4sKt3qqIUKPitEz6jM5dQK+lEbdeQHB2nhiVIkROwkakSaVP
loEvZyH4XOOTBzzurxGYQ2MVUab0h6KCDHV8qf5O/eQU7Pij+cuSSgZlfYuhYpXj
eo9UlmK0rur1mIQuRVLvhpXs9HxpYgl7odyM6ZscGCfGil7rsf7FGgmHIhf2p5Yn
F3x90IiS/ETE/3z1A5ChVXnC6iaxyK3MSG2lzBliiRjMPy6t//BymdnheC/2zkcn
OOYPaM9deCEeXvr/x32c7tTjMp163cfSda+N8SsfBHBOsuU/teMgR9can9JLc7NZ
lKaJOX4qc3m+CJh0YML0oNF61dmI+D5YKGukP9rLVSWEK1SQSqzqTyhSIv/weKso
cFeJAM/7CA3Js2h6w0hVE07/xGqtiTg8wZVLWsqqa+LbkQhcckweMdkjw7yGMekU
OjpzTxShYATDlBTZ05r39TFK1WCtRzLz+4ESQ+HjH3M2jFR+vWd8KUNPalXlN/6S
OR3PhMAjtwYoQA0mJVxojDgyQVBaAl7lSL8l9aR6iULWWvg3YFS5219DxlRirwJg
mfBtlIU1uPbkvCOcYcRHooUj0X5dt8AAagCk7ytq0VQPqRCxnAm/HECgL/bpP1Y5
w7pz0yTLdbf6egH3mi9TFgmdycPFaAlFW/j69EBJxJrBvgYE4roEk5EgHQiKPqHS
gKWjb93c4O3i4t6OrXJO81g21UyLbXEgNcVoka8KF38U4shFw8/5yG53GXP4JukA
MfuJfRswUag4FsFrdBLs7ZBx78ynGigSL6AAdktVku08vtqtmbQn+YhNMa/aif3J
P+s1SGltZDGQq8kYrC+qh+ENbozwXiXF6gnYpeYM4tBIRu0nnKoQXQydVEpo79ID
B1iY0LDDoWQJO0vu1VH4/heE3Ym3Dr9SJ/g6KM4yDJAFxWJRvLl/fDnJdcwSrwD6
iyD2ZoPD3p4uXu9Nf+TX5uv7Sq12suJP3oSSoJW66uyyYG5huTH6Gzcw5coroJrM
6brvQgxTCPfDA2cDv9BnbR9yUsHFditjBxPEiJ07P7ki4P0IhsrNTn2sIJBULjZY
GZ/6Ca7GxYe29a2vDND5dCSYqAASeUNdOhnH7QbRTMg8aEpU4FdjJ52Fy+m29aWO
EOywMjN1jq6lwmqVeUi5Co66NT0ENXzrDMNLcposrPLPjDdwGul2DGmd2nH7EVET
2E47hVxBAgILrJhnwvPmaUE/oe898oH68dlgnjhHZESWNnJpDRQCO+gdjyXSV3xH
vjwepuv5TkIWztFP/Q4hO3llgQ0qM+R62p0LRvLgqXktTy96XXotQnGRetoN7TtQ
PjNb8Vvmpy33rIpqv7MHrY8OQO4lVFFxbvF2f4e82lLf1nmdpNSHZ2DIOQd+7Bu+
T8kOh04jd16G6xdOyxdLH7QqnIB4pZPlF0PFfcrb8+rqoKHy76IxeMIjn0IIvrLi
tEL7QNAyk+nOL4BFLTq+sFZv2iCVZ1CcvcLzt9qTr6aitUNUbBR5K3t/a9cPEwI9
oeE4vubcxhzQxh7537chkmTp3M1PSNjn5BEdAA/UzvRlnQCH7fxmXZo45EyDKRES
qqRzloEArbZ4SxN5vlBz+JCB0JRx2zUwZaXtqr2MysIwC4pFxT+u8FLFCHAF16Bh
xuYjwFyK2C07Itbnxdhu2cdNhzkzsVDcWysZx6Ot4Y7vyQR4JkYQFbEQh8AiwrWi
KfGp2g0xzBJtjNXc3jYb7RiscWU39SP/BdVVy+rgURnGm8gYhX6NlTjx/ZJ1+0sJ
7bSkCuwv0Ppx8pXFwRV5Ud7akRzl5KkgK3Ji7W/JkXO1WVbnxUtBPbitxsyhyYEK
zdh/Tk52/CE/InikurH970fy10sX4rUyz5YLzDTamdMlQHokMmyWPmboHZn5jQyB
sD6xOTmaATchD8zGfE8Cmpd7ePwDGHx+T0cYSuGnM1bQfZMFFDN0LY5F786PcBdp
5jTRj5Fbv5CZcdaRc3lTLH+3vX/N1fmmWvgM0Iq/+PPd9uMK7oZdf1fkyb+s72Xe
zUFbS7jfkD+C3+2DIy5Vm8+2Fq8ZCx0XE+tRLWTz2IHabUPdQZxZJiN1YPgSqcrJ
Gg16O1jD7H5RnXcAGBUeg1TX/0PvE1R/LeLDGxFHpozT6UjFrBLsj7bwI+F0uN59
VCe3EWVbX97VyPD73gEnKueNKSj8G9IMdNggGY/nFdo/U9YOVc2VGoKmRv6RktEo
AZZ12LNpgVhwWdIkatA/TGLbAxkXl7HaBb6BLJd97yn5+b89HtF3KVkJNNCA8erG
qg99YOY737VGdyk8CZt/NgYkvilJBM8eixzpS+HlHKisYHhbOMzOiEHzGdKt0BNX
oVNKWJg4/iY5C3lcCyiz8iPfSgAagMWPel0MMklPfwNLSPV8P7Qng578bxs5Zu6q
o4QOhO/VT3ZaanNpUVOIthmB0Cq2lhztENShYRTajnSlzHUxMBrvpAf7Of4iiqXx
WK9u2AUNPJOIA0rJQpmoTFZk6eH4qUrlph7sy3h/IlCH1rLO3iqetUqj8Kc+7yov
3Ool5laOPHqbhQWh2yKrpFFBNguAYnSrYOtYd/M6RkAyoB19zUiU62lg6tNP4VT4
qFOGGPle+bogvjji0+7pfpXV4Nfq9S6IaiKN/XqWl9ZbwpwENidF1o+7HHNSV7M1
Cu1367rXEmrz4QRgLzz01ZoawehRut7mGf6Wv7zK8s0j+WuEMaF0zOPVRQxOJWLl
sSSV9U55/DN8JgNUjFUblwHO5tTetBohx+6w/viTm7OhhU9j+SHvw2QGAZvDGR+O
GTbKiD/zgYc/g5e+k7l3wPEVrsp4Hgz98p2t62Rkyv072kfz0age6pNOmbus+uoy
kmpzUiRGiccufaj4UTURw03rds62CGJVD2Bbs+eGVQMVGhlsc4WVuMt2T8nk07Dg
SHYRxNTcC6ACrODzbNBpjU/uXAvK0wEUOd6d9W4ihom9DX+dX8m3/35eTAgOQmL+
Ip80DD8l8mmhd9MBI0PLdKi9EHnTXI4A6AXET7Ai+cYmCL3YWWJvWLbNB1jzxg+K
FMtiCZvSmkPn6/55rzdHy+7BRI0VHjG8gMoEoJhy5BsaAAZR1JhyUnbsMTkAAgcy
DvR4cXvibrE1PVTCiyr2+VH27rsyyS72kV2vmwaPiqUe6PvbVMSrY0qqy5C7kiZj
2GiTWTK3rE32pnRZx6WIzqvDfmlOcJgTtwWjpWAPDi+Ybmi5OgCdYAwLT92OfKfm
WjiBHdUrV9fDDM19Z/ZJ2ajtl2dIAtIt09CbZ89sHLusNXP8WLJfh2afpponD8PZ
63NmVL+FAtapwcQ3o5JELxg4rS6W6/VVGDRQPLvQxTpvAgz05XbWaDtK07vL1A41
f5/4+0b+zhDdvgz0pylhuGyWhWP4C+6CJVwox1l5q/P+pfiBL4LgJpPKPycfjpp8
4kGLxEVk6RrHoMjkzkB/jfufoMwgIHva1MpZtwxoTNZhjS9p8LErzhJO+NxNmPM+
qpudRbMNt4cHHJ9Hxl/4AfplYmlcKEjJIyGXKFm7BIqLQN+knqOypFaQiCxBPjak
hQesXTvnoHvVGE8WCcKIWNuuMphayUgqAz6qW6K6gD0zYjq3qEyqduncBoETdcnX
kA+p/FbVFfGbW13CP8Z7gXwm8GcWLwILD5lzov8C8NEh3FbpuHR2ZukuXjwYK8/6
gaTGORTLTqU56/9jaeBduN93HTieAzVLDx3aj74WckVXIDSIS0UOG625kmWjEABh
BHIsVC95cxUbDFddvCGFjE+Ye469EqxuN/PYx6627YH0qV5iJiXfRFiEn3oazIA+
Yq/lcuQw2O9v7hbW4cb7Wj21wlzrLPLkM8qpGLsQH1mnNOltukJ7+RLkMYgYwZt2
nUJUoGIZGTdqNBJr3AQde/Di2QYYRBFt1akQE3mYUdPQN0Ct/CMnbzaIwNiVHp8U
rHYP/Hezw6+gqR3lpNx6gChIDhwzqBxWrksclOueSiM+wOXBhdR+ax9YyUqQrdNV
ictMbEreFFXUAGi9FmJ3y9XCmCsHDNlezA663udGol/sr3YOl0+O2/HdYoqbhKRu
VB4soa4w7tScR363LWm6s0mEWp0yCmZCGou4lkDdO1PIUXKaEcl1UgwdhCXWn5Bq
IGNEx65k4xIxq2oE5S9oIu9lfsNYMB+BmDF4Z+46g0InOI0rpiyvcb+twZQmPdke
QMjst4LwPmI7SJF7qdLYx8qXDHmEOQgNCDS1+i0vTT8NIpxvHwJFBIpB7ayYA7Qt
jpfwQDFEDoJjswbB/ZXzp3bpgc3OgbV5rXTrOx0o+T46+D8RsVrHtWj2e69J3IN+
rV2dAiIL4Rep8RcA3ta3yeKr2Q0bS7HahtQdu7I3B9Jm/LI95Q13gVE+fj42hPI/
GXFL59BAy1DfZxqwqCdHSDTH0i9NjTpDK9s1GWwsKvl9GcKojabYh4DkKOB4j3Uw
VYFDDULJxFte9TrEVkdQ8r/zTiyFkdkPDzwtAL6TfC3DmXsDTkJSXqRMssn385Mn
vAoyoOmnhfIw2Z5PGLAPB4ZZq7ByI+/OGG83exerKUpkK7it1MTJKQwTyaPvRxCX
pSUgxwslA6x7p/MEiSQot1t2sQ8e8/ltmzhIgae6HEvdVcWN+HlbX/uRtCbXlVQU
ijC6fiXMX0Zhqstp4FaRynDY7Hj+2NmKcFwu7F8nV2r6bMJlXNMSt+okXAiDl5Cq
LXB6ot5LMwT/Hgc8iNHwVL18fq7+WZuuWTkdtFaFdo2ZLY+nHZvGgOeQWRAGkeEN
RJDkm4ddfIhD6Wp2D6GXF6eWSIKPTPjWvqU0zFGeE66EFbsAoi02EV9CHPp6KzrC
JT2o8bMEQuXz/60nUstZmV4aKVVVnC1o6Y5GMFRhV5664Yc9bjuEnsDCnELCaGRA
PLNYwEEBJ16r6UYCs2fl2A0SzEowe3mKCuOgZIysCpHY3EI+SSmLIOEZE9Iid859
c+qlbLHwbI90fQ6VT6VPAgyZjyN7ECMO5sMQ2hlwU4ntkh3KG7rNBbgXobnmk5E3
8756aeLXIFIpqnA4v398BRoKswhR1Nmh46y4pPKIzXyyNb6twrvXw14440PJRdjo
0nq0dPnesw2MO4lpGPjqqe1WwjBwKfeGzhTfQosxU+vquLlTCt3nkVSFHy0fI0oY
En+pNSGpNQNK5BYIfkV9CAdRrLU2+fp2fy9yfhx9X9exEWH4xBCb5pBGRzYVQkG6
5OryWDKkPs+ZBNfHWNKOPi6i73w/xarfklF5dD4CDRfSOqRtgXnVMyydmMfjqZ6s
vFuCBkx9Myu8/FKt5NpaTO0PpKHWwtu2WsXwV2SMmOy8k/q3ub9Z+eRXrD4Ni8iq
y7dPEKO/kYESn18SlV0PRKN/x4rRq6lnAwx5G8sX7SaNZxWCu9qcOY3b9vIvxX8q
pB0C5zRQrntgtPP2oyY+8HvOtBQJa/7x6Y98o6jHoekc2JFb6wM4IX2hydiEgcOx
osy1iEXOOTUTM496/8ooPz5xug9z+Zx+kB7H4NC//VR1amB3KPbx73h22ewhueTb
sHFpz9hMcWY/v1xlv8dQa+OGos96q3K1bcmmz4uForooMKYGlBLw2H8iiyOCHYE9
KBN9LLqbzU6vQHvcdZXWcu18GNBRiKRQVVN+R/ZkpTmbTkrxQFoPQF9k8tw9RsDh
QNFwlafNyyc9rrgEBqwSGdERLIQMvfftE+cuBSQx7KVbjyqnPQm0TFQof4waj1sD
UyV/x4MQuMM7KmepYQjh/F3Rkx4cjBxpRk1rZi84CDM6kLezzIXohwCGND1ueRc4
tF4r4Rwx5jP0V5rrdrYgS1RCKs3REwIm7m6FZQ6mTK4NdtXXkIIUATT3wST+JoPz
6AP+RYtcMrB01TB1XWsgGejpuX1P7kAGMMn13SK3nz7J/LgeWygC+JDsc+ff1lc8
rVVa7UrMolJ30zYEChhBPjebKIb4XmfH6MbTxd6M27urvaZCdXw1SlHhsDnTAUMC
M7/W30IDsNGronkFEmJZQ6alDdYnCk9IoIWtH8BnDsECbTJkV4NnuNj9mE8tpPwD
mA/oKVRsD2r4rgu7+Lxvw7Sit+vJNiwkRzD/F1mzyZLhw/cogzBYlGYKHlFWeBfg
BmyafwlX9WemGXlXuaQr4Dk+OSpApR8ee80UC9+7YDemuNpzEKjT/gLGKcPjQJzH
tL3BKYLzdeH/ECUYxKP/Zp72BVhFVC/n6klf9sZMPX15X9JfQ29cQN0HJdNNPc99
oQCNK2/KCBiGp8OSP15hcL6+lpn1UHrWevayORc2JBVwnPIHWmxYcYusaAMW1I/F
b7BzJuaNwH9x54Y7qePaEuIOTOzV9FpePyXmqV3ccsG2HXBnCleqndh6B8MFsSXk
qgtpWgHu53lZOhkQW1DmLPWumUg3HvNyn3sdH+SVDB/fYBp0OOCqNmTdvBE0nTsJ
xAsCzarAs9K3tAbhspnzvEymSYF47StvHCDQOKAVY2GVxo75pChZTSan3D0FKhTG
Y+8sSaU8h6YWFnDtUe/g5skYVOAq/ei0OFNm8cgUYout/wbqXKi7TqY1jKDOivCo
D3cW/5VtJ+Z65bMJZcTgef2NBjZi0nto48RLUarPRqRBF6Y6DlNHC5gTcd171hbO
46iZJVL+s4OesHsF8JV2V8SaQHd7T8aKG1VdQL94N2woR1vy8zCyps8323fB9WiX
3iG8ySftsOhjIKtS4bAXjlDtEyb39940GH08huxCoY+59dpegx+NaFQyFi3BDt7G
T2RXv+GMqmXzEbtjTDv6kXukQTJ+I71cDm9cY6jWNdmyxYfOhYVtrgXv06LZcTxa
72Nzi6QMVJ7G1s6IZI6qZ27BPKwpKcfRGZ0yFCEZZswseGIvfNjdXXOjlZnkh63i
bD3jj3QC51NoIbp35L5ZdI0N2IN9RPzm2t3igmBnoIL/lEuedGAMn9uD/1Qd0bDq
g48y6l5yBQTFbPPvZDiZ7EVLngHJ6ufx8/irpr/swhexGNSQgpK9GwJEJOa1lWhW
mD/jxnJj0tYzRzuFP3XSSTPu47L7yhmZwR46fSMdlP3ibq+uCVex1fShIeEFOFXB
DjWKcM4h3y0kBGPnOTNMe/a4rOq2LeeNJ6nt3eszurTma2G5iT2s6sp2KDCbP95/
RJePXTT20yNkkzr5IvVqHFZ9OEhRp7DKGyXJI7npDL65PRolDDvIPQiLt7PKVULf
8DPNVXuqhuY+e17ivlFRdm/XPapNR2uRid9bUZB7Bb8VGu8MSdNWbxaP8FzPWk/S
qgsEhO1LCUBluIsrvWtuWtLB7Kjh7GIMgIppbKBHTrS1Cz4z8mhy3r2Pp7qjsOFH
+wyxcEW9Ip/Av9z/UD28mbv7q40ztRlMdtnK9NpMe1aSs2zPXOCrMBkwZI7XBbYv
Q3NMTK+UGSJQbkWeh7h4Jv6cF9xGYzMWiG3IWMLBbUa21QVDj1I773zrRZ5XudYU
6zoigtIP5Va1p7KVcUyeHpyqJuCdFCXvAQc7Se+LCmJBaGvtKY5dOUx3FMR580Ol
2fiYyvOfkJ9wIFbD1OulZf1K7OYp45wE8GEbfAO7rMyp2NyrrjlOXO8rvulcSUz/
aLs1Y4qdQBge/UlHgfrsadJWCAd1b4RVtYeFDoyz0vufbpSi8WGSzzP/FA0TtjP1
YMVjl+55BoHFb5bdUnaaaJxq9m0ru8pki3Ph2vMCYXkz+u5wbI6Nnu5oGME/U0tF
N9WMisnrCp8gBJTZaQZ6KxIOtiWKubnrdrVjKfLcVBJFel/N8Rs5Mb1RnSAMSX9J
6Rcpce+EDLJZmaSppMIASa7pCZG9RQXzNPteT0BL3jq15I/kJrY4+QT2KsXQfD0U
3RpE8a+WRLT14qd5NfvQNjnl/fubbpUOb9Cj4OQ0ex0fkAuabgi6ePv06oYREtkL
O3TGJ2q0jKN4dXKRL7N0HTkdJwAvR0b4Jbgvca/ilza/vjcSv7qtUJA2Bc8K2BMN
jynsRvnIIh7lfxaCmsPFvboPorhUIZGt/524tVBxazD3dKKZbqizatKusa6JkNHB
oaewDAi6XVo+xOz0HeosAUMxVAFq9sCId7ttxu2wxu4E7mLuKsuN5K7jPfoBbcXK
adr9AzoCWaAy6UPMavcyuh+qdRMUgc9yj7Oa8SOrEyuvkDd0Zm03ov65eKhczVQI
lw36P+wm/V8NGEkKC4ir5h9HX/xQ7nwRv6NonIxEPnhiDZ9JygVy/Bw8Lz1oC4Jd
HsWYClifNokbXslPCsR2M2QP1h3M7mwyJWqoACCUMooxEAE9K14OXxxM9sUdGhF4
YDeZnrr27+dcHUldsv3ocWJWfF40YE3SfjYAIuFTn8U8TBYcqdt9epU4CajFJdto
wPPh/KTCmbFIXathduhHs2/j3hhiseb1UFJ5iaHvoGqZMYxNNG9E4aYt9cUS/EV8
zdUpQGcBB598u8QJvnnFrbQ3hxgI7zKU7czE5Q9DmHZTA+BSFlC1Lifa/sazeH1s
a1C/F/I631VaMRRgo3QiUKQ5SQMJDcgcQj9xOymiI+7e7D5+ZqAEjtqcshKHg79X
OhYt3xmasQDa/HD8v/IQUOKYPLujBNRDlFoYfv+0WvI+AoFm8qg7Tw84cY+MhEvF
sQiIxkZsCYq9tXcw86kbDSkuOfz6Pd+L2j0hwlbKDkI+d8cB8cHmgBC/cgh017BJ
sc+92aO5H6hbmyaza8wjQCNhZvEGWBVKQ6LnrtmmEH8hGcW4WzdHMLk/7vXpKYbr
pfhaJylZ+9Xhsd5sPgpp7M0AlWObkMg3n4OY6ODKmUt5A9U7C+F6aPTx2qZHZs0+
3cyqBO3KRxiUc15vezK1h04HLNG4s+1Em9YHYehb6BorZZwiEiJtXlSKWoVUIKWl
RQETH6pLcE1fRhPXx8XFUCBjMdrTmTH9wbGI0PB3Qyj0u2XRdLOTvy2gZVmX688b
n8UE+7277vimVyM1oCHgUGEmwNFZihUKirLWInj95RBnTI1lF0hh/wB7V69ZMm/q
9Yqur6vyCbbI3k3zQ74RbM+hmGhBAwLh6RHf9TZAFqbW8m0njB4d4ycYDy6TbmM+
j6mwWSGstySkeknGMvgPFK0a8e5UAjrlRwRDI7J7bkJ/UymNeIMj10cBoCvoPF4I
dc/e8VxBfxz/g3SbIkc/zM1Ei7NSgWlQdMzwCUwVc39OxV0k1Sj57qA1n8ODhgri
hgDgvT0+vyemDyiWk/5cEfz0DJL5mVIZeB8DmmA+kq7gkuHeiIRLtlBUa0tiUOCP
oTnxd8yZoHurBlHen4tXY2hj8IlJOO1bNNNGJ+qiBbT2nfhtxbA25e+OWf/voGzu
Kaq0raifnC7PMyXXdfC3wRg1jMgFzvZ5BgSt6xzL0L19L2RVajRhI4z8Tm49GbJk
6b4FYbVBXMiLEBKtUL1B/mtYSU31mloR/MK5W6dGpdXaAQ69tXVBoBZ6pVvJlyNb
uV9uJ/cbpwo/nSHMpCOiuLl3rGAKJreJ6dILQdcnsbUFO4aHwghsGysvLWXpw2w4
7k7ucdEHRaQmAEtLipwocufG4igo+cLlmxYPTSkRTgyGI8rNREmqKyBCOb9ufa1x
/u2DFwkcxQPHPSgwd684wKSST+C9gXehNC/kqfVqdV637a0USafq/YlYrdQw1XYB
37CSRTFZGkeXogIYlNvz2gY43MRrG1aG2E8OnGcduxS3sP0cHsgAwt7HRMcmBLa7
6YOj5wIcPms4gq+7JyWivz36l+Qa2ef5X7mTzpHWdw6f0J40nCXnv302AubVLV59
LQXcn6t/vZMsS7LeD3D6nz+xub0bWoGZDhWpB0whwL2SqNlspEyfuHdiiID2oacy
ty9mOVECYvdu1cvvQK7u6N6EwlnzpJq7lMlNKNrAlnqAS8CEvcaSng8zRON306tX
VZu9kUQx/Nc2tWvpONNpoFF5jfcNWmbIxmerfMJamhektzrecc8GhceQaXrWtI7R
N+HzU8xiaUsPwnO1Qy8nPjcGoTi06hKPx3SSmWBlsGD9mHCbwZ1NPI+kemcHgkSo
lJAUPc6dh4v2eyghiqC9Z2Xc3Oi7/9A8uqr5JWp/l+0ArBdSLIxycy01RyX2s1et
FnBo2djuz5QUK0zY59qthEAPQgqoIzCAhlgKIJwYS1Py3eO9gEPj6mdHRbjHUsI0
EKiZp5vAF5szd5UCXC1XCLZonc6U/wuw2UT8DgN/bfsY/4V5Daba2wBhNTLewTcx
4XHEjQ0bWf+NeKI0UYNC0vlw1e41yQBZOFbKlxrQxELMeTGJsjVVZDp11bMq/KGO
GLSuKfUI5TkI1Nl8W7yxt3s9OPT8+fQvhk0FYrHwP40O03Bdk/rw6fhMXVgjVYGQ
pHZ1MUW8OXDcwF9qJVJaVlz8fqP7XyOvH4+f9EhAwCIyZFuvlNFqg4FV3zRsVptp
JMTMS1QW8+TqI4m7mdx3nUJ06SZxpzgfMvhMpaDR4zcOUpx3YhEJ8Ka5SKxMLYqY
Ioljhu0MWFOPdfE5O0VNXUhHxvIvSeuF1dsNhHzGnQvPDhldJiN+C3FnXEA6w4Z3
V18h44362B+QiufEd2k/+/8G3wFEl/yLTxSOsuJnQjJjSYlPTy93Zz3/KRqVWzzL
gDk8USNqlD7fXYBOhwl+9GScn28DzEjZJUWvEdwpM1NiJyVHcKgj4spQU6gAksNE
cfM1MsToOJm/17NEV3X2ur3fOCXE9NQdC5ylhMKQK6u5qq/XKOV3p7Fk/rmL9n0k
CNLJ3BKnzqqpeQ+1K9eSqhko6868nPjUt2GxxzdKeEX+dGTXpTNB++fSgzfA1p5F
cNqfZBygJLAGE4Q8fH+aax18J9DPb/fpng0pEb3MxU+0vuOEdbd5CnvAh8bZsU6V
8OcBp2KgzYfES6MKszT2i+cmFWHTVLpUZcZrenSZk5pyXYtIUSTIkt4rIfUZbeIi
iHJmxU3mzjYc1Ey9CC90iYqIBvEQElZsMeiOn+to97/avqAux7ADtYZLt06pDsd4
RdtfuzP6Tohpn51tReNDlV53gS0v48UICfBi8Zz4YjsYCRD4r44Xfph7o2nDZdJi
2bMSmxID7BdmFFMSog7EqyUmxfLm9p30p7WgoN91PhUhcBi/qZsJG5OnekPLDzJB
KA37XwOXz3WRdwpM/LEC0TKym3fvusYGDqM2FeJuqc+tZTpXjG4Fekg8iW/31AFP
7M+Dbh/d1qbQS8jjYYBebKjNsEiq12yhrlVgj5roym72enahxMAFPJnNqqg8DyyM
VE7Zw0KlrXY/GSfa8SE68VRIx4PPKKuPXQxJEE2k8vs9AkfkwjHB0Lmebpwxr980
DkbdfkMvuPkbszkZ8BGsiGnGcyRPc4REfsZwJWic6KmFwsljy6ZZmMv51536z7Ah
FxY55D4FaFy64kiiFnqMAPsSVWYZoJOj+uoESTl2X4khIA/zwky/r63pUIBusLzK
4h2jryUhwojK2Ahfh2G/Yl8DkHES6EEBulPcef1K3kTlE26863guChxJTkSEvkjt
2vxh16sHNcs1iDUz6eFHP/ACpEb2Bx04RWZiiI6Zw/srbZuZ9K9RXWUrRlgUDVXW
ju6LfvjV3lxig6Hnbntj16DrQBUxuXIh7wacM1MJoVbRRLjDIrSx6R/VAz25Ch66
ZIqCl+42F7qWUXXUkbOqPQOAoqblP1xJzJxKLs1kuAeRBGeNb5nnp0JbGV+37mSL
a2RFDl3Rf5iBVj6UkM3n2WY9seaV31v7PDC22kkOB0fH5cybZHA/pmhbcda0oSVQ
JbUVeqa+NHqwh7uWqosOU/qnR2K6ryEjOGrLYYg8UYoPnoawmbBKeYeVQa6a6+mH
MYBL5O7RySxleRwguJdsR8sh9fahJWVhQ8lsqCHix9O5u3SnCCYRseTHUfRFPDNm
96eETJM5tGJlNxxGB0JU+z2UUXW5RsqpwihLBBmcahOfjILinGHs3aR+jt+uPEgP
fF2r5K4JVSGONnPYvennuzxy/UDHAa2HKSKO0eISdb2p+wlzazd/A4fyFcS3pGIC
I/FET4lAL2HgSwXsfaOLSfMmVRQw3/Zj/YE0Cuhtr7axMw2UyMWxe+ApsyuHA1z8
V1/oTqhmBmpW6HNFOGjWLaa4GtGuhf6zPetEvNymsskFfCXo6iU1XLO2bSk2MPwD
z29jVl8Jk3HrhFOTJmkyFS+DaDx68Sv4Ua1HSp3TQ/vrXAKt6mlBiAYEYbCm6qA/
Kc9051yLRXebH/i59lrSszaV7CcyEIDprHkccQSfp9p8lwPheVY7898ZW30vXEKn
FMft0B/70adq9LkaSUtySSpdVWZl3ja3XgGm95ZB+fqYflceCoSzI+Cpe/5tYrew
q2QgTf67g1e+T+0DbWb3u/1bxirjrfPrvSwR+4SSw7hK2lPiWs9TXw+9IS32szFo
qkHPQuu/ELNsPC+S6BrVTtgIKayevFiAgITDOs+ApplD9fJ3wB0cMyVZZ3Y6vKqd
bedGn7bWoGeye9MuWXXaYaF4/Hyh9DxNUJcEd2ywNmow9Px4Rj0dp+bIC8P7W4kL
rvQ9jiTU6/TyL61z2MBQf/A1qhn+dAoqy9hXBxDuzOIRXr9YxmmXvv7NzWtz4KC6
4FSiN2HdOtmp9+oNbOPAQ4Ys0rcSZGaBB8z+LRhCQHUIuSgjNjEuA692Ywx8xzCW
kqguESDbUbIqbIeDhmx1zCYOP0C63SFt/bkM7rZlamTOfe9Qzs/bE7/VB6QD/9dF
kz9R21UVm/zdqHvEVA9vn+NrjhhOCiHpZFn4g9XmKgKx9IasHBxCVfyH1i14kaPm
wGyBLUTaIiheI4A7YgCdD/ZG/ZJPfc6umc4UY0LcBpYyDOTwyqjidwfhMt5dAjMZ
xbzdEvjQpUhpVj2LxQGqSykkHzZes+QgLVAT0jeFm/W5z1pL8QJrK6QJbQg5rQ79
jYNKhxkJnEasyy97jY3Cjo6tomCcCrYK4u2Ipfjreot91H2ct8PKbfHA6pUPTQno
KS/9XOjb0PfRZqpksly2XxIDVeKekS270/jvg4jsGF1enTtFwMGBPRSm1rhClduU
DNdzGWfFqdAnG6rmbBFSuJE8zaRmRCaO39IYPRpAHjySmYiAygNd/9gg4bex2lz1
wfi0aUEcUfrAsw6DIO83rma86xGkUVXp5h75Lj3ugipd9fRWeK4OZt01nMlTlYGt
peoLWs1yf2W8Br7Pab4Fvzo2iBRbx6iu+plkoSXyO5Oxc62MaeVjjEa18meubeO1
Y78fF85lYEzbawRDzTO2h40noIZFvIe8YJr2hppuK+aZI1Skhh1WeCQ4K4L8QxaS
agJmNFsrtodAnmnq5mkOzhuAs4WLSeHUCRbVTYvccxSzUzdezaWDQ9f032TWuq7/
ZcE58RI1Tdu9NCUwuv1PNmjeQmF7vaa+98PNf2yTa6obUc71JNsZiSldXns40/Vh
2jwSLIPfjPnNYXOH0RxEErCMzI/pbb1Ivvyg5ZAZshvqp7gsDB5v94x34MVJX8h/
jEXeOLKYGWSyJpbb4GxgeqgvLu7Z3YLDXwMJ3sKpcjwf0sxZSXOHEee3h+li79sv
03Oepb3XxoylJKnKzOQ22mJJ2H8abo1y5K1qRU4kbVAdGVtjfmpwk47MajoirzYr
xQLLUynwZ22ScN5AxtEEvlLBQ7LQ7auWCZXGBwNz6zHoh4FAp12Flcoh6CrZGBbf
d/KMyFw9bQG9YqpKzb475J0Jy8W3/W27Tq2KxtZV8NhgIJbEYm8thYHATFF7EeUR
OlQjh5TdX1Ew857betu5mk9CSBLrLGHmyZX9/GUOcEwyeh+4PPg5IK8f9XcTkenk
V8YsJPeEs0VnzYENCLk50uSNidgA7m5zAtdjgYd6SmV0QwzekqI6WP6lLDyO7PWH
NoPhnWW2F460Gn4hP04ltXJoQSEDkCJkO0GKB9RxW/0qkQ94NbkHb7OqTOWoKUjz
sgEhKAuE+BLBD4tuIIKcdC+nrLlzT3BbCQ1RC50Cuf500u0ZMJYVcFl2IWD8wnIE
LkxkH2O7Po/pu1aGozT3qBA5oQ+CwcUEQdd0il8ThJVEEtwB32de6dE7PQtLEPtc
Fn29oKL/g2U2X6yKqlebBMZ0JUm9VAw8ZO0s3t6199L/ZN/WUc5TKFsKmRNdFBVu
6+/T7AxRCZsuYsS0BD0O/KWMiaGIN25dMrukHmqy0Su+WT7D80rqxt1iJV6+4Rcl
tzkCMZefI7Rre6itXB2jg+ZnL9Vjn9tpH/QTE01BUojbOLSUcVwSqF+mP8XpMhZU
hdgrhR9I9CRgAVfHuL2zVbRoGJ/XxPqCfaq/91xqQ8DynPyLmg9Qq9iXiw8ytxyX
7dgCHylnxqzrLUxABFo9OwsUHsRyecHxBtFyoZYEyJZHDm/3zd4f0OzTg2BAG8dF
7WEBdqDqnrQlQxT8DQJaV+W4GyBUljts6aHOnWblq9fZNZDswHApsf2mklmLhD5I
fWVutCN7wZ6ESOHgf7rkOHYQJe9d2D5XDoBlsxfgMZ1ZbjZXkBX54vY7uf3oubpC
fou/NywhrGO4e1plpwCuuLWQzh1zZk3SHpEtyrxapLXQL4PfjlmmUFbNMFpSrvfa
CKihV9eKZ0pj9fL5zW0AwW0nQCeXjOlT0IsrV92Ohm8plaglIkUQSLXwz3+Mqj3j
z2Y4q7G6Sjz8CVosp8SpWSiGd7uJXQqAMnPFjztqecphf/CCFEZSrczcT6VroCiB
hLbgS3IdEoq1GnGYcsPvZQmOlnBO+U7rcpZ+mplhnS2+uika4ZzAtMnniXQuIINV
4fYnTIbZstHo10km5jkJkOVekTLGJOTmomFndFp2xCH+QMiUqf4n7+yqcCJENCiJ
845rqVeN3GeFgY+h/r59TiMWb9EkOACPACnR8FxyYISXu+jJL41iWpWc1L2tVagK
sirSXhoIaO5SlZo9gKPJsh3ne/GuR4bsynnTl2i52Ukwy82YQKDbpvvFcR8PBd0l
l6vzlI8VHqczBGRhKAUJsrmq+VnlDAp2BeK5oXg06WYkJHOVUzWEgiVXOOQFytTO
XPXhs3P62SDtj51MQ4gjSBpQzjhRUWyTqXen7QIx014XeDbvIJLTQmVyBo6cYFaM
wxEVwb04Orm8uK7qRx02kEJpv347P3zvbnmx77u971b4pCgYJor2oXToAkpZzpxG
E2Xn7z58mHMmZSLLPWWvf1THQ4mXpoGdK9cjb5p+7A5dYRn0b5dczKQk1RvHRt37
E03jXjijTuqIaeuWTgWEXFjNpnj1PAeMc76r/w4VF7L/x0o/YgoIzuNKU4/eTtUc
LpV0IPh1D5Jagu2PdrQD2gkFLHPOSanfOTqRMxBSQ1zQog0E/1SrZHmWjBruHXK4
OdB0V4Zc+K8C1FFmGeXSlC3CRsY6Cm2bQ7MSREdOKfLDJuA72hZGKjZRGPpIaMba
cwmoDdiT2PAb3DkHbCqzgGz/YKomQFlYbHMhXrQxBdWRKZ1uxj3qOQT32faI9/Qy
Hh5oWDDJKVzD5dD6PrsxeqFtdsY+N1hsdKPvfgZ1Nk6DsI/wsmYVZ+OPQJcPcQyC
q9Bw9MqBH8WUN12+CAfSCN8GPRMmUkQdxBKCzT8SzXsfQKVmgStH9dY7+TrE203G
vmBfBkaoRi6LNUvrAjDOhoOtGK2i3ouRTZ0dqq855usYnBRNXBWAdr8O4KX8vzmg
11rNGYBBwXB2+XFzeez7wUYYqOl2KHN/kwTvBzNH4YcC1YLZc4Vi8dVtR80f+YeY
0m4XHonNxswFgdnf4LDKSsqwGW0wp21TT0G6k5vhSfpOSC10JIkQ4cLMMFrukOJg
2qSTjh4H03CwSn7zDbTBVTVLwZ8QuGNrVbZw6MZDORg7E+0lEcYvZjEtMPlaDiAE
7RKpq0ZlKReC96+LPCkQqHoUC+8vtIev/Kvamg1nrtB2s2KiwYou2MEKvGCHfbT+
zT02hjlHxY/rxi0AWCARPlYkm7r68XRdn13bubcE0U7U59KBkU7WfCqu8A8L/V8y
JOwveuwnLA/QjzWK4wHoWhs//Cx2dQ3gI2t+zxvjwKrYTqyQ2cnO7FleOcZ0XrW/
U8uU4wduoBzO6lq0mAdZP23bfU44jMnX/4f5VkyVDJYTbw58q7WKGmQqF8qOEvpb
e89h4XoILKiKTNAj4nbVW0/H34uQV9qqHv53tO5/xiT6xUFZQt0Fo4mM6BdvqjZG
LL2C87bawA4NMnILhjGdgXbGR6BlLRQ+Lhe6mc/ZGWJDoSLmdH/5xoAicaE2bGaF
dBNcVrnb+Sw+Vs+Uo8JC4Eus6GrMEu7NE4L9/1f+cIjlW6hWMbM0tlG41rHnTNBd
93cK9MxmDY1MtynjRox0OHaybzqnWMuze3EJPnRN5HjqZZpxORWaIwQR1tyBRvci
u4RSftbiyFFhJfMliQFYNMOmqLsG61YGMDLdbB97A9InxW8Z0UUs0TbZbOOS9RAP
XJGiSUEoEzzu12xQqY1+PkxItJRVYIyPj07uMib57zrBlISRkx5B7QyIDUW389z+
mvr/CU9P9/3GRDki1Tf+u5JNDxe5OP+koFzjltzHpUTIOOB2FVV8qBNeY4CRzilY
bCJ1jkBiHO0nKh8OoeLTGkLZNWP+okPvtW2PD6DnZjdz3ECrbrBYvl8kI1t6st+I
FGqyxP/3o+Kpd2xtdc1jpkEM5OD6UqpTdsCng6PmBoF48Jp7gfd4mtcLCnGmAISk
MNqe1w4/4AH5ujTS0SVXFLfjmLdoN3zjPUxJNmIPiLDPYq/Sx5JPsZvcU6HXNeKR
KOScPPlg6x47+U+UH3PyGO+KXPRx8Kfwja1b6hu1hXEPO2f6otXB7kJsgXmH7oxw
J0tk5BMq5eO0doKyk1q0U0DHL4TF+DH9Wmz9I7eIijVdGdwLLxFJK7axhs+YI1sp
9YhjqCjTH/3TV2D+BMVpz03HDF6+7J1Ruie6qwBO3HsRBC4x/H9aZ0ky5ulQa8ur
3TGcyJL+VEfOswMUXhKqGfFMddnOvbzjWn5qx1diBTWnFjDW6OEDYJIvY3uytR8Y
hQFr2NbpyRiCP302fBVDGWh7XrXgcd1ZiPVaYR/xBM+5cFD+NizKsskVlQz4mLd0
PsBvXlR+gAYZnRLf3DQhOlYkrSIvyC8Es92M6gKSlfpJsYfjzyMgANZAZnNjG5f9
luXfYZJS4Q5we00sVkSJNnM5vVQqEC0GFkNSwoTOFDUj6Ra22WQIQ0QOyOQIZmGs
Iqt5O0XH9TWX5qVuvN7F0RxFfSTip+19lNKpDSuH2JmIUe4a62ZxbNAX48tl4kW7
dLp38JNAqXSBIjXVGonh2+PPuKGHO/NC/oP3IwKbmacxNVuHzHRrv00yVPbBoM3N
rQjJBYSNR5OoCkdma/BzTzM4PN0A75lZUivI2BvfByGm1RcbJvgs95704d/V0BBb
as48Qv+LdeiMaRt74Z4SQ1a+juNN3BjTuzl25YbLBaMUVHaXqvZ8eEdg+LdQI2Or
2bfyp5mbmZ+BkGp8hmQYXZlhoPuQ+FJF2WlBFVaBT5LRtw+K8SmdnrLYnmN6lOu+
ioW+ew5U+k5YA06O14gPW4GEhdAq+wrOuiFq5VMo5RVAmu9nw/kfTsztqPM/6tjC
5BN10N0js4to8M0F5bCafB+gN9iKBm/NuTZ7Wxz3DD517jnOjoq6wT500ob9MeUn
IJmml3QhKUiFNGjw0/tyrCQNuUjcc6b5kT0XJe1Tr8bvbp7jdrzlYAKXXn7Rgfe0
xSd/ChqS9Na19jHpQcuZOmQU9ZxG4VtWAKQaPc691yWSX6nkxwIVUM5F5s3euwwW
5WHQIxV1BKL1OMcI2YT57dq4nTKQWXhmr8wZKCCpj5b5Q4P1sNz8MTsuOeaWJOrb
Tiz0mgbDAk/L7XlebR6hlN2qqdbHxkhdQUS8cJFLQw+qVNv49VeAftW5k4DbBShJ
LVMx9XUXJu8hl8U6622ffY1w87EuSznvAtYZTN0DHW3JaPek6E2/2KGJhtk8C4+s
Hge7KiFm03OiKXB1QAPPIeETkNcEAg53S0kNwWFXumtSb3Hf947ZkfjjX3tglGGt
l3Q60l1wUE+gHziHX4T96I3smdisacLmgfVgY7AzxzZUcwZ/kAaiY4vXo1y5GW3d
LDZ02Z0Xo0lmUk73h/lim/o26mCjx+LCqO9gSwAKzoeg/mntnsEA8OM8QfyY4Ry2
yydHGzNpjlHviO16D3bWXclhSutteq4+4Bu/7ShwqR9pt8K6SijR7y4LOVzzZ74K
xW4dLy4ISRa1PlhuQSsb11gV0JELP5S9lY/Zf5iJpnUQB133v5jKmDRHt4Iw1NMC
pfViT4f5Tw85R4TZFXlRmw8yZaAcE6ecUf0+kMn/4LVrERZHiKSZQqnF+HIIXHmM
y7r6vo3IBXrpEmS24P8HjDiSHM6TBJXn2osmS+VnMpQIQsNT3MjNHUQAP9D2Banp
1QXF67DbUKy2E3FKyocJAHSwYdfJ26lqAJMkiHtrhmkkGR4OU1OpvzL3DBINm1KV
w20rDeYrZ4xu78biG0RjRbmLlYhpaG+9R1rZB2DqKbUWoXkSysvnVCbqYm25Nnb0
O6KGCIvtgYnMqlxfRt0UpjjgBWSCp/cRyxlFyw/nVvTAvo8AqAdYlmoAs0IIIW5T
ZN1clIRGPPDIPRTqwzppCvS+Qh+bJ+l8shV27rkjvm3D4kxLcU4OT/KzbO5QEQ0E
BcneEMI55VtHM2YXV3DtJwUKIJnBVQa4OAH+EOOVCj520+YVWkFWMONMuYHvPsFs
i3q9dA22j9ZfWnNWBpU139eRw+nAWb06cY3L3i/Pg2gS95YnVkgFpSCjW4njVAXi
KBL6L4k4ozYvIKpueNJPRwpCR4Iey/DByqcP5Dr1oKU+z5QzAHdc8uKSCMxRP3O0
khFWdC14LgnLX+qA1QszMQt0bgDHZDcv4Mc8rzGurA6O6nVcEyt8N4WXzZDIMBQr
Rt4m6TfxdnvmtOAXZKBLzkJC+06qadYafCLwiCEK4AAiOsupCOLSaTDiDQnmX55B
qB9cMHa6MfDrlLP8tFUpaNzuFoKVSNx3M4TPDIHoXIDWlhltusXm1h/AhW3p8mBp
tgxnD5sH35MlKRF1Y7MWbN/jHi8wJxalo8SCh6ZhG2kgmqyeh8wtRUaEI/iauu/T
WVKdmptPBoOm8kdgdJb33Yt+CA9QzMqRrcPFUjOWd7Bu5RDuudpWt6zUfW8cxI+g
uJKWyCvvlDK099qMsOwlNySspllydnuHBxnTKLCIlhCGC8ap1xs+jGbsKeLaiUV5
g6wQxIEu9SXJDZnJBX0xsnzZw5uow2QFDEreTTIFXB1EsXHmBc0i43GpBgxonSOv
64eSTh5jcov36wpnR10/ezaF4t7OtuFrpOMdRPcKnoDPuFaNHSfZwlq/xVtgZbUV
hvhRgNLDDAhNzgYcKj5xmN/wSD2dQfASJRFwhH9KXuM23Uu7JCWfIUzPTF5C0AyR
gDfepc+p5cwqLXTNZgUugANXtsuMHYKD0vR3eqEv4k/dgOvBN5xcceFyQ/45QPWw
Olcu21QIC1CFzcn8wOp89VQQwRnp3CLg/GTOXcFF/jhLRfu4ksM6YlYfgVHfsV5f
HmI/0I/zEzxNA0E9C+P2e1OvfW1prhAxq3vhB10Waz9JKCg9odr1OOzaSDSl/JmU
WeNl0L4iUyrloeGhj3aha/PLzrpvFfJVfT6/1581KPpry078+KSHbqxhN3h8q2bO
S0F0S2jHgTGmDFWRxQusYhJMR4N8wyOrUFisiy9fLs5kPOe3xCtQYBSWpwzj1C6S
yvaes3zEvuIg3IfJiydfBDQjrD8uUv8GsPZoLQ/+S0YGrtTkMVLjDaBRoBor6PS1
m9pDC00GJsPd9J2EADAj4MlvrygaBJDhxObnkVLjfyJcZZU3kztRt5p2iABlzK8F
+OQNuWAY5gr5uRkhfu0J89sc27dZ0arsGWdTf9wO/coy99ggMnxCqJ4Oa/m4/7pN
oKhCvX8OeCHmKuNV0ABiNQZfXjH6/aAX3fF5h+i8Qthg1bUC47YQ6FBicaj04Aq2
H5u96p3oPnoFOYtPj70BN6Zdpz+aNI9+Po2LG/l+jAo95aUWagBuPqwwTFPyJKfT
9YOl3IyarhIjgGvAGwivh5xxpAHe5h6I9CxV1vdTcEiLSP+ZGarmHG0bGyZlsTtU
D3LqcbScs1FLncO25lAUy1w7ENZ4bHIVhv1Gax6o9BTsXF3wI22x9PBUVZNX7XB9
vvp+LW+DGMqDJ9ckyH8ChJKOhcN1URMiJCfqLuHK+RynaWdAY+pON1ME538b1jLd
kdqlzv0SeYDLuqoF1+J7lIJayvem88Y5FMG2BjftW/94Hz5uW+9jbK85AFEOWV8S
qDVKnFQXs0BFRHnUjj2jBJqnwVjWd0mlDJGlLk6a00iKCA0VB9WXlHTZZMI1hs8M
cLl5nKYpvsJuFqA/I6aXFyQP41/HlEV8pJaA370TsW5jpnRBRe6liprbSu2sG1Ax
sMTJzbtGuVvhUFIHr8EI7sbjX41wn9KdJXIrPZRcdJ4OpBoZ0us5vAAvApN+LJpL
8ge3SjFaD+aOZjQMF5LmkvNj5g8T+uoF5fAw5sQkyfGF2xlYQgU9T8TmllRyhkrk
L85qHitAV2NIYnpWbytzCDUwCQrevvFTv+GJzGAGnTMbXyczjqghDGhJciYiirf7
1boRrnriCodTE4T93mYGu1cszPHekmaZthv22FmwcYfgnHMTlXjd59HxtQMhPZL+
eKitt/44MVkxxbBqc0Jd0wR2hepH/M7oA7l99ll4pYdc6XfJryYuSwaXVzizESyK
dHWAcc4nybwSTxuf4OMh38V9EEANITJaRjHufQGoYSGl3GRsQPQIjImj97H2U9F0
+BR1cXh0dVdLZjgJiESMFiWUSI24+yRoUeljPBcA1JKhdzQ4rSM28L2ehEjYwXIa
8TNrOjLIzNNZW/Ob0Zyx5KPzdHkShxA7Y9lnFWA5CnaRBczSAIMgmu+xCWLNN+6J
+mnLjbhcaMy2w4AWTAyeZyKOpN7UuqhU5wlzZ3gMM5yh7datSh4U+o+YM/qbebxD
eWD/lYh4Y4nzK+akpQTmmAWMr4/8ewJ5ixdYirEHUhjFJB+oHugjRdwdDU3Ht25t
9WA+6O6GQ1Tn3gJgYtSlflD7Yo+y2L5elpiMXw5kO7dT2PdyIBmw8pbXc5U6MLts
sqxG8iAk3XgwQw5n+HGOMm0eYJ5R3i9fB3c9A0OXLB1SRGoY0xH3mOmwJDkAveTw
UJLxUbdGSGUOPadfT13MCrQ7g0dqamo3TM+Sm6XAcOicq5Ax9ZIsKOU78L1E/DU1
+o2qlbim+8gpel//xapgIwVOUEEYs+RtN1DWwYt4MrDG3fryjnmaw6TBOUSzUE8h
tOQxOaq5tvg16kRVh90zE2d/TXV8F3ybHUrsw1OgixSvzKmp4lT48r3Gs7uqU24T
sK5SAbkEGLgRZwkmf6LEqUs58o+mYUcZ9LErPIN+gUr8GRY6H4Nhz8PnuuT6CUBP
CHnymuZlSbO9GCdDyHNbkw5rawY8D5WFD4VdWxAqMheZPT1L0y4DJMcHlboSCf6R
07fvE0T6uTB89DkD6zNnrcIs05DKl/d2hHbGbCPEwd+PwAKr8hdbsq6G0LzXvC23
E8PDmG1e6pzKA4t+8T7B+hU/RFEamE1tmqu2qzBFvC1DP27XDqDj4iRvFDSOVgB1
xAeVT/eet5Ewx8RpDLSkzuS0CNMm44OCT9TJrW64UAeF44z92C/BVhdBYk3V+Hpg
QD2DrCCwGcIZXLN4NcjGTnN+sJGeGt5J1J0cEOCTNcBYDueVt7u+hBQBk2/cDdaF
LdKKc7kMswjs8MZHbwuWaf7yiBKQ3neWVZo8qj9lg+a+IlJmL+ahlnG73A71iIBg
gbW1lyY0RfKXeEYRicXMSvWNNGApByf1ae1adCBwuxoFaMh7chaCJTfpHoEA5h1U
Kk9YSTrtVGm8UCuxGjbsrPJZv/G2Cn/HSbnfRlBX+/UJHeEXu0M8mXLHywkrptWK
P+XQsQBXnExdO5YE5dsC07HRm1rLIrAkznm7ywjq4QBe3ddhjqXxqF0F/XA/IXf5
gkn+RCPbLKU2nG1QKJaIrTb7x6VH/pqT1vwiCYnHfEbMOftHmkweEtchQVw1XZEf
3Dt8+NTErMGJMSPIHjyL0XFaSBHvMAHQOyNZkjKGt34mS7AeHnAIWyJKg1qNqfV5
1r/BA3mnhHDVLQWGfAMhbuK3JooPvLZKMaCER/LlBNBxeQb6LXRCNe6p6B2vRJXv
+O4UBGR/cemJrfu9txNO6PjEkKAaTN0nlMjHNZ8hVD6ryYYXpryZvPrUDFNYO6FW
rVvg/ghJe8/eWM4RkYL9ZTACa0GvhxJVWmqjZTkd5LOY8JPIg+NNbM0iJgZomoe6
7WNBbzvYxnpCmVTLSFfsexmVf5gy2MVS/cUgnJZLpNKChdInV/8/cUJNwtQ0WTth
wlFX9cOujZKJ3rFVEjXgysTW0LxL0Fp+fqWXlZtg3TszEVJguZyMWKtDETRlF5H7
qQNNSRzkvduS2arm1jvjRBSaDS0Y+uQYzJsXKcugRCdw+FjWaPUK7Cg0al/a8Au2
YUym2+jRxtDR2SwU+xT+DFtWtcefpoifBHlv2cPERvBrYsoL69w8l5SzHAteWIe0
JvKqq9JtRG57v5GXrg/Cga/wbt9X45M2+cpaSBeg690U4evF4Bpue+CWk6zwDcf+
YdftZu3uqFeyv6NNHOAs0pnhHUtGl7Y57IuXfUnIaKv/9OoGNmwEp3KWHZYrWlLD
cznr74eKIcGohia3tl8erAWpMX9FbuQKZbAg5/gmvdXekKzCudxVj3RbVa9nnNmK
i7SfwWOhqFOUjp6tb+/Je/Pyc9ntTLoQ7MGpeBXG2xuO++DFj8dbPBxZeUL8G8gR
Bc9mOQDkbAThwQNbiBJTjkKk3mMUWxueAixYoy9a7zPLVajaGmH5kJVZVnaGQ9SA
tWlYNs8QzLaMJOJFIaej4M4sFUQHPItsAuhdLZrYrNTF4sSn3SCkH5A18eAjb4qE
gdR4ah7DEFQfybKVT0ft0B5/ntnAAUcuz7IerVfdcD/Q6vjB4YmiMKll93r2kWcG
6zbT4FQ0AMZkB1qcHLrxOqA/tg0VpEFQO0cMJ1daw/vOCMx3Ko5Pe2vLKjYwIQmo
EJpdASsBeYgNHoMjxEbxUMKyqqc+d0fttoY5T5BDxzCHRdyNUZeSebcZZkFuM7J2
fb9N0XYCxuo1EhpigQ+F5qFnUfexjQL4iNGpwuiYkwHJMTvCtOnojPWumWZ5HCUb
jsz9STNnXiii0lL0xUBwC8xXfIoLK+83kWCfzFpT6t7Zk69FHo/woQlTz6PdunxE
7nnb6Shm0TjsHijOqhrcfZwk9U1DBN5rRG9L3wXjPZMvn5+D6XM6STvEIBdZyM4w
ZnBbcBjdkzK0FWyrwQVgJ0mwt8IsATQzLWwVQ0CzONDh+oyT2yfmztf1sX0A7hn/
8ybim6LT7nvu88Hnjtgv+JQJFnYFei+DsdfJVxPcV2QWLmlzR1++2YggaFHyZoNQ
XpMOhB/F2oFkDc9c6OvzTnn+Lyb71h/x1UNeS0IeMuHtiK9+0445zcivkCBWBr2y
nWzg8K3sbmwz7LcWc38mTXbTwqchj1YpC9ezeWFRx6fQwHXec1x5MLsx2Zp3qke3
v6BTdV1O/EStGC//cTSnDTHwx37uQHRLo1zN3kvlyVQNWzY9M8SmUmLEHohJvMky
VAH4GWJSojdN2M5TWy16k5AMN6QoOuARs0tOgkvdUMWOsOiO1XCrMavduJ2ofdL3
WKDauIN5dCJf8DOW/ZI4kqxwd2YvTPZ/40N0j5lHkXYLMxCuCLnEDw1PQqNrtqP4
HhTeY3tJq8lk8GfCuPEv1ReshAgGUylJOyG80VShEtr716nSwJZCdoFTrBDTOKh5
4iX1d9AAiepVNejWkUkcbW2tUOtALggfeCpdrLxsOJiu26DEcs9z/wrlyoiWqAmC
oOu6AeesjdUSCAIQum4oKe9N+JOBDfY73ou5KFASYnIHFn4FQMrYQXyiq/tMNhie
o7mS6p+TQrPsuCtyLTDFb5IQAmFmLhAsXImv0bVFOAzq7kLq8bMoHEhnLV7B2uRd
8eXlLKrii3DHa0roim8cFBTCwB71j0zBtKtfPYDQ4C8wus1AT141aWuM72YTGCg7
eYSMdN0BTLlayvAhFwR6awkVGtvsowPbvxjMmr0nSNKQ2xZOAWn7KmWMcIARFE+a
5ZPF66kVIPJplydL/IashRqNBzV5uQyulJrSfsjZaiuNyeSY2jPv22kN0ihkFFAj
rXDK2GcQ3LXwaJ5Q7O+0JM/AC80snTzMmElpFOqmYQzzesqt3tAC/9ANQQZ2NSXw
KA9CRTzhuy7ojJcF3eGf8MTXtolg3snJUpVZV0foAQXyfKxe/z10NLf6gJ6UZEEa
7gGbaoE1UnOn3zPMQlPh7h2J/rNwdDM1meqi4neRzV84KcVoE8/4EvE0TfrzA5cE
EvO/b/OTNJOmdTp2bokFinttOGoxvAkiNRFZxW8W0tBcxbOUiyOze+uX0hnxrskV
ZPP92jYGfCjIiHR0ccDU/3A6Y/rdy9Bngjz0G2XJQ7NOgL5tnpp3G+RwSUseVZV8
2Y25bzYg726G6GzIhGg9d74Bd4Ogjv93TmBVQ57HIazhKivuYer/3P+bHk0YAfKH
XF4W3oKOyC0WXYN3d0zvEmsoBRYg3OAxV40q44a4bZ+j2zRf4D7wqoDym7B4NNjO
JoLicJXsMWAK0f98wV1Vuff9dbW8C9zR1cJrgTUN+lEpECvZOmnPMaF2kcP9gB0+
C/x7aU5McxcWRt3pPl2WX74WBvUkdONMaah8cun0aeRzgZApFrdfwbckaofo6yxP
xtdWPbe3mUgAF5mesDB2QNrl4X6QUuffxTFtJ4sCjjsm77kV6d0LXM0PzjVCbW5X
h16mPOtRe4Gi6QmvPXMi7xWBShGk7gq1z999/wY7Brpymr7136+sGhR+0CyX+9xi
M0bN7etH68b3Ad2JO8mfLoZNwppxMKKphv0MJbsX1B4mIU4Oxqfc/AKVJsDrBm/d
InBJ+fQtstxiPWzFNBD/1oYDRx5f0K+AzSAeQWxvbQJoEVIvYBicSgN69iotbxZu
fD1Tmgu8VYPmEZWcIw0nGgXoBc/4AWLoOL/dlhqXeigUpNXwqPeTzIjMbL/wOmmU
1bju6PFxcWI6Rv//0c5jbcqJdX18e8w59RzaXTBVAwCf1QyhZ+uoeISQ0sBfoGa1
JOU4Exq9nX9sR4oxsHkOXBPNl4m8GgMRp7nppik6su3nGJ2TgcUUy1XIWZXgfpc9
EjDP0fUw87uCru6mLFL1LqfwKqgQgr11HACe5p8/+sFXSrxRgHnaXESXjGYSfSnc
TCNY/VUr4eJ7Xs3/REiNEXIGXU29XuIGJycniQ5EOtJ0GWiFWTdWqukM2WnZfRrL
mnDMWWAO8RL8YOx67ELc6g53CZwaMDiIGNtiI2cVmpslEt4xXvbwTpQFQy4sNw3h
VbabuhVTNHqgyQObwokDiJjh+A4yDvXtR3SpzQZn7uvtEWxYCi+/aK66vhhUuQKv
LhoBj96mukpd9RlpyYshOu4oiiKYmKeHb2zAL8w/EnMmIZAHqyJDO0cmB2ke+FOG
668B1YGqiz/tAIj7irdo+BQlANJG8X9b4qkmeblNFd5XeAOkcZ1NINe1SedjU7jz
SgrGyp8Ivb+Zu8oJ4ITrwILey07fzKRf4Q3bEIXz4B7ueThXfgPHe90c+32uMave
EZ2n1ryKwC5QVnuJSMP0/PF+SHNkJnGuTO/F098k2yHEtnVGE99lB+PpXUbJf8yd
55PjVrayKDHcl5kSZn/JJamXX+se5IBoQV0GXv38l4hJWTa3LEJTCg/LCRnmqNN3
XtnESFyDxAyNgG+ChgL4lrKWBRzvN85m+esY/6ZCKfjThC0CE7siROrRl2sOUOWv
BKvs3NFgkYeYOniSskKq4EOzZMBLFZtOrXEsNmXNcqEKshZpigc9xYK9EXYbhDqa
XQdJIroUbtjUevDz9PhUcTR8/fuffx+W+w3Aeii6BmkZ7JWTcdWuxKfIFFBapOYq
74i4VDaA6g2fJ7alcxYDVRKNQ7z1Yf+cABuTgBtcmsxOnpVdQGSdrB7G9fyh+xVz
bCfwMGFOynyLiJ2l4KrKlW0SQq3KKaNHZvdpy1Qmv9y2z7MLqpG13x37HE63NYmy
IpG8SrVN+Vv2YpqIBRjCZnX0YVkJLP/EZSCNNwMwBJ4TGgTNOTtttmx4vo1Bd4Fm
bl5fB0svYNSWNXHbDXxW8QNjPZ8sQhKoOwajGAoM5qtXwM7uWfOx/CZV62zfeOKK
S3eVgz2wSZIW6+9cwFGl/FsljVbKEoJlru4pGBBW1SqQ4ji6pMGQ/ukDbxAiBWQK
NQ6H/aK0D2UMVq6zD3CcftBWgXAQagWP6wl0sGG8+HqMGKqM9dUw/SbUM3SCGSLU
jdEUnKA76uyDMh9TCt2AMnOWuNf9d/UFpagUq9DxUHR5PfXv2R6Cg/3MULhNoaNQ
4+ZDwAbDNpPRJj8pOrDo9ey3uoFykXMAiQah28UWw5Zoos6r3uF3WQ1awlE3nN+k
WWuh4I5kug+/yqmq3VTFBGucJyzESoefCYe8pVWHycYVPX0KglKV1Y5D6uwaQXfF
ejVAeyUqvdqBSz2y9E1mS8zqJ4q2ic9IWNSdja4vGJ9RjIpVt8i7yH9BhoCPvs8I
+3dd9jrVV5XIYOlWDTGDcDbYhj/LIRRRvuXV4uLvoZvKHbREEgWoEWv98TtL2nP9
Byv3cX4i6WiKnBWKhK8WbpdZ+nkojoY+YLrdlDCuiimJkqqW28+33npt0edtwvvA
N8V3HkNlikTwGG+BNBC4r4SIek+vv1ZuVY0troAIw0Roq15oLMSN3t0CT/EnB9Bb
/QAnEwCS+BuKSyOj4YN4wThWUc1tCaWYgO8jjlJLBQzc6fqxPohr24iT0hA5svPu
Tq3PT70MKW5RQ79UjWhc38YbvMYCwyfrBfDWmLFMB/AjQUB6X2XSC36TjKExCwLU
NpqZ8PLP79irxrYc8V6ZtSrVXR0DV8+BFdYAB+1pinZjY3BbTk46wDZA3IGAIZeR
yPYgNZztBPP1v3kCLC3tKNwffe+/kQl+uHOMtGXccq3j19S3pGjzMgNsL1q2NQDv
nXWlQeTjzCj6mPRSWD11ZnaqUUrWotQk/vwb4Oq+GJ0+IR8WSroZWbiQLqQEpyVV
pW6avNsIWX5HyHvtnWhWT7DAX/QrW9rI/5ve1INhJtx7NFwoj6b3Ca7+3IrnE8ex
0lA7XPkSAW9kBiMzh8fbbY7M1x2iYPUdh42GfYzpAuB2gd+SIaWeFTlRShXjCe6h
169RUuXDvfvDZ7pQtgQpCNZGDWyJwDhKN7vORwAYc6/EqchTNW5sRGDnb9Qbko61
ucujUNKfrPfj7MQhX6XhMfWYov9ZTGnehhN7jFysaI/BfNghcE8wV/jDkVjp3pCw
u0t5McDYwx7U6G95UMX2igmcXSSIu18iT1uMhVzHYA0YRRsGOONoNm3b+gyY9vBv
Ipt003+w0PYy9jy0y/1PD3ubuon2qdJHdsfH7gM3DHCNwEDjAIvJATwM8I/q0gqG
58J0shR5MGGjwuPiW9pWydMv1UDJ3Lf79taDAlg1lEB8KY9zh/BiRMSUwZ3zFoqH
rmCkWXOpXvZBW1GO9gnK+UaYuk0Oc1gJM4ft5m5MG0bjFt5EJykdFu/m4ae/bqHP
1CtACjjYDLmIL8WphtG39Cb68b1Pvqui4FzblrBf6fVPAZEB301dSTDYepWCGdAF
VFKCf0fhKBShW5x/DxAdAvIIPxzYtluycLyf523K1JD6DApVj8SW/WztPg2CbdYK
B2mrv1ib2+5aIJT3bSOvu97dIeVVcYv3CLjCs1JVcNqIuqf2Dq0jeyWHIKOsrPwL
Ahngg2wMFV46CiJMJnMLuSv+pu2NaJO2MdNUu0ThAPfKFpE/alv94gSr4fKrl1r9
fadiPI8S1/9sCt1Gj4nTVvTgNiUx74xkaNZkdHg5g78lKm6YIcv4x/VME4OV4b8J
FwxLPDwePxriS0RCQ2JJhN6Y4BukftnSJ89hkN2TPctFFozcJyCU5z3r0AJGLboQ
XJn3S5Slsu+hSi1R/92VvDxow9PxNlm6Z3Zl9k0QPCgJqUhIdNuVS/tJNaifpZ/4
bt3biBzQhJSfD6kcgsodjxIVhSGm/mqiVhz1vSc1uUSFZXA+QsW9AAk9OlSWdeUQ
tLqr20MF1jfejgvf1y6RHBJUbWPXJXLxzHndivlW9og0K8lmA43k6aCx4Lu/Fked
qOZt0pr7fVQImeUGbr1dIfkAhXFNP5Tf8mdDnQ+mwgGFPYwddaaAYi4baiMuZvoQ
/x4rR9kZPCl7KZhMjHIMqB4CSmN1qc/gT+MhpBOsPHib3DVcpHojfHfPZVeEr5lg
/l8URBVacjSGFPRt8mycqEmGsi+kAT1acimJVeoVfvUFADw68jEMZqOkuJbOAQE4
OSi6SzmjBwUzwGzk75jOyLUXb3xRT1CBI3X+LbCbupY/bMHkAJlght1jCTTkBXeH
FW+nf42+qQW2LAEjTuqiNMeveaXwGokEnon4w4UgEx5RlToAbWRJa5Y9mcQtSjXG
0KTlRbyebSyk6aoeu3sGnimn05o7xnGQsSBXQfotZrq6NV+lbfb7Y3VOi1YXIa9J
NTaTkkmgw8gdiVqHrvesKT9RlP9gGHMk7C0kTyffJAx/nYsolnuDVkXZGXyUFJQr
Gx4j7SGFmXfVIiMftF1kqxiIT/nFf/mREQbTcR1fda2sCNLz2oONR6Iq5VC+JYWx
jEv+kU29mzKlaMfcQOeLeob0GRCD21Mr8oipuqgDhnn1HCB5XkoGbAeOsRNo+1jP
09F6miZQPBi7ACpgiEtQQALKnPyLTZoI/ACPPDV9fExDCy87kKBIA7QMPFuK39zI
yQ/9T5ZqFi83mXbGyIVSUNzqI7UalUBL8LRF0QIIDqydqxsxA6vKAGGSgTVy4OdN
t1XMNqISvfp7RmOHGJWQLdVzMZmK5syHVSgpDVAq+jEFRNJNkz0CPdJCArbZOhtl
Zsv3U0LwXoLs/xujoEDGcNy62CMpYfvS+pi4wGH+bWxgmKF9WC7o1yG5g6g5J5fS
MuLA4qfpNKURndfKk63J63Vpv9EMlIwOQ3xLZw+Yba2B8UbAaVBEJI0SFnXEtW6S
N5bGEQNdJwISJfn1kA9oUzt+pM0Ze+qktUJHSHHEusc9MkvieUEB7OQKnLbxwmhr
JldPAYMM4fefNQFHq9eJUuUnkIhAR9HLTzLnzSe/cTLUdXhMtga+s2fnWaUpqmuA
Z5vJv+nChDD9gtNj/E1TwgnibZHzgd0GSUmix+fz99Ebn7DSHe9E9v1X8z5a9sKE
qBmEfAz99rPnU8vBc+ZLkRbdH03ByrnyLc2/nvOq1/6KFqKNz6DgA4aUA7umCc9Z
zBCUru9sYIh6QykhT056Z//1/1tXwtyV4hvVlJPxuVZvr9fwYjIv8eszENcOfrnx
I2e9k90e3+j4i+8Uus1kfd47kRgxIygBFblYO2vtxZ/NIZPmz+n/ktN54qyEiX4p
YJDf22hfK2+BO98wK4Je1icQ4M78o6KXLPk1KHrv3VGMhUuzjByutEIBhqFFswmE
Jh0cphVv9Mtp269AGQUkbYj+aJBPhfeQDVDTr8XWaeN6prFvWUw4KEU/Gz2L7rwx
6AinBHkjntWCo9Ge08RNlA6ct18olvCZ53qVbOtg+Ao0v3wS43XAe/c6FjKBXw9R
UGLCKUgZq0wOmeuB85PrC/bFonBZ1hCxIMc6Y3aSR8irIhg7o6iRTS5aJ4jtsFHa
7oyJP4OBHOQfzpHtY3eLlqDSR+X0+rlGqjWqBwa6A5eVTL7ZYPRwsBV29t3c0ERX
EOI294b3YfXxq7NPqv3Mo72WghpiWWeypn379nwu0bW5BBQC9HI6azfF6y5hF0z4
z1UqllaJ3EsIkLC6CI3gM+yBB9UhskqpqYfdY1q2cuDmsjS552wIyVBvhJgqXsq2
rBzebHTmsvm/d34XXuUxfXz/kEP3qO+SeG2vf3F6CDb3o3uzfC9Ro07t9BAFgUiB
ALhwQzkrc4X/iS3FTKh99WASVNODS+KVyhlTlx6gn6Au/wIrlRmwcm/CjF9Zcfwn
90JirZlUgOPquTQHRF/s4dXRVeD3IOoMxWy3aCl4fUVCtJ3uCygnE9BUk3zqkTr3
TEZx+wqJ5Zg95OZXT29knZdlj4rwyo6IomXslgp+qJLqJzC0rdTJlp/Ktf0YbYDU
HZIbxVE87ZJBcVnEt97dM1NQ2lf3LnJsDN5PLTJXQCiAakxZeIuQOSRkD3UuIVmh
pKKyICnxQUQOc/gkTbfQHGMlaP+P3HhInxHGngPmMqEyCRCwRTzEsv8/jk322LFJ
RWUsXYmEAtjsZDVyYnilFoLmk2jTuwjgOftf1iAFJB2ejtrCSxA6pwd8eY/F/TDh
3H2jaaowQq9utFfwQ4iFBeAi/ws+9Hms7r0VQmj0bd+PSiRYKoru9xX26TgWrAYR
HzrZhNYEV4tWnvYrXd70PgSmqNkiTz0lMIvEiabq8YBmC2g5rM4h2V/ALYudyuRx
aOAFOkAuSt7n5Frr3251PhjPzJlBrYyyqhhXVSwi5i5Pk5kWrTeEyEwrNPMH2Hgw
zZU6zbkhHf7pOqUZ1MDJF3KN16YKOGeHk3kpScXxgqVKtzh3qSddzqU9iLLLOUVE
CcZ+8tNN0Gx/F0pQCWDl4cUY+uumk5ClP3hpbsSS5nKocCgLMXA/ciLYp50zNljY
QobGIk55Up2g69liQWbBK3upr/2XK1OliuzeVAP9XNLKP87wG15iKyd7yqjEv2zo
IApta0kna77UCL6w9GfghMAP+NmTucfGeqlnOzri4Nz5Bab32oG80LEptILkoY/c
lZZYpNo53YE4Rv5NXbIuYJRT6TNt18XdemfpMq+Lf3fwdDrkozt7/lkMLFcY73Oe
YWKCAynzLCmXObwClu5rZoNzeeD9S+lOA+6yYNlvyHaRCM1PF0OMxbRIbVP6OVgu
jN2IVfyKmzExIREcBU9G/1qLevw+7fmZhr9m2j/8/+BtmhtpEJSxoEC+h4DFTndz
He5skn8l0tBEopj2rTd/RxIgd5XfISWaKBIK4VZJ/BYDhZi/SgyMDkspXaPDVi8A
VYac6gDTZpFJo9Uc5tlyMA55ZbZVNROfwZhv3uxzIr+bWTOVBZz5YYeHaa6h6ada
QSDVouSbPf10CYNlXY4CS9bom6HfuhveNPnvGCzixpD3nLlvtnCIRbJtg66P2fpm
OZcze/765vWOQwEqXCu3O7strw3NOwgnY+TgVvVVaVHrf3fNWPpu/v+g7FGRghmu
rmFKrXCQ4pkzKP7jesJv0lKTYjpt0GYFfpVITdzVn/y1FRZ/DI1da1u2jjAMryPt
Cr9Z9tFcrI4ZETIuwS1o4UZ+SwVRJvEYFubtPGhtHyWhN+OKCfxHK52hhvVHdhgc
/Qae9JDto9P7xtSzmeORi9yxd+3X4anS2Bu5r17L1uayGICVlMnOv1cnGkHweaoi
wHKFql3oaJdMZH1q6lKpghjo2oWEzdZ6sQes03a+nfdDz3ngGH2ZJSb0bM5sOa7O
9T53xYhJe86l2sTnQfQZXtBD48v6zZHDFjBo7EXd5oqbUYTaswxFxV2lWuNz4Ot5
OaD+G8F4SLFaYHDmieItvZLoQKSFOW0INmiL8B9WZhQYTgctpnfyG6rROZOOxCsG
paJXxEAmGZ4VC+EThWogAaiwHaROM/gujjdjHLkgIt7u4xua8rhHHSma7nqaAa/9
8VsJp8xlALr+NQa7UB3olHWTf7OWan1BW5RYPnxdTxvXqRehAoAuxUhPHmN6D2Bh
X/cL9vnCmM9iPuubu1eQi8nVW2R/VI0hrhQDqLlas8otT1sLFxchRrKWxUEeo087
2Sx8872DlyYB5JPEfpWzkDHwPnpWmAzDwp8Ok40r6cudP2tbMk6pstcwyr9qXjiB
ZrH1eIJBnLMxcfIzTkISOM+yN+AyN3lD64z7UTpkjMxav0kSECqlQkkqeI2SzaPs
TKekAU6PisLKrgF+fqczPSIV364MFzdA18EklE+T4JTnD2ZER5j/6JyeS0O6dWhS
48uQaXHQJu4QZy4z/iq5EXUUccExZTFHPKtKDeTbQX1xdm1FrGIvqOUH5NJ1rwXw
qUxLWfrNvKZJgGizIybQ+uEWorYamXoK2zLRRVIqc6dNXP+PwWvMsdLtoqAFMfhS
uOcY3Be0Npa2qYKdcGLacQj4V8lOXGMu4CT3yH05Yy19xy+LvT0VkdRLGwnKzphJ
Zn/hI1fvaVQ2jfUA8nbEE6xxzkmXdczQQuTteDmID0bFpG+vcjmiJLd+8hMd5ywA
GBBJhyWnDhfIuCa+Jk5w7k2xQivWe7XswkOk4v4q5EiQhYoODxWV6DMqrik+24W/
uvY9yILfNiiwK7KnbtvmqbpKq47ijM4xYGCPEJGdmlCCcKDnz47icCAHfcHK8Wcy
3iJxqCmcTjppai3pwrXnQHp0Y4A8ftiUu1ab64cOIGIZyVZp/pdEpcZg6BskysDg
dVuS7+ULqkkTBAumyOyYYdnwTOcGdzUsrgl28uVsHCprMG3PpY+Hp/QJ5Sf+I9bz
fJeaqwhXZCz49UJpfMkRSlJyOPCk7OZ3KKeHMmVUUpEk/EyqLvPkstqV9dmk+AAK
/Rvn6vwLgLHxbeEv2KzEMo5COrCn0u9oVlPFsLJ/kN/FghRiYrMP+C1DuaoUGtux
LqZk79JkrrdPcn7Yurq0HDA81Uk6EDqVqiYgde5DBSqrwrJist1D905K1SFfSFpc
7/+GRkZuftEgOgeKnt2I1owPgt6DnQFrjFcEiOZRfwL40TADWm8N4ZB5GioRhtfS
OGvoCsP1GUWvqr0NDSfHYLUrYYSZRRP8bHkCNV5XN/41zbfvUWiUBrvUtu6px1fo
qKgr5QtOOMn/p9gs4V3pfvo10N2N2cyglwrbSn7tPCWoZNNRt9HMLEVGapOGz6Ag
GZb4Vlhiav7JfX1LplukJV/Vj5iA81jaXmfkiUv7ohwB01oeWEWIrKVJUJSTWRT0
0RZgcB/Hg1fFtkz0Yv597dIj4YKr8Mm7Su8gXDtaS7mDlsQlFX7wXrZ7n0HNW54Q
uCZ+SqSuYNLBhs12Po/MTD/bgZIbke/bNGZTifiXpXkTyUMaHnbtmcqSXoSD9Urz
1+xKvKB59qDXfjU0+DSylaZHIfNFcW1s8agueIztcs92XERwoilHuRjdqyFmxcHC
EfSOyK/BXkzLVDd0MY9RyPANYyr/SkokTR3FTmLIEgtw5xo0ehfq7P9AQoAww3HK
dILRPPGcwBtjVHT25gQM2E8w9Ox9MIXjVe5lk9rH5GddSDGBxObZ52bHfjf3cSp1
gsCthjjAAM+nexx8o+GfMt/rWYQ0I6AEtoKP7pCEZVXLCO8NsacthqILkNat+WMr
b7LJX0ZWE16tlCZgmnEuR9+eLpqwNI/vDck7fLGpxMeE8XHFH7ukY7uSdxkIPh66
if2dYVm5/3lLlrBgZemgZxUr8tutau6RPOc1GxhYV/w14WdqtajxVS9MguK+MwxV
4nKxRC+0/pigo3u28Pzd9G6lzqX3TGLdEHY1Ta2VW/f4SyR2R5gR77fFEVgRcMQa
2eCeRKKxXuaRZu0frtNHyz3jd7vQ5M8bgwxt75l8OvfcioDnAqJAAoiIrhe1x7BA
hQe2mgv4rul2WeTUvUZhx5KWdMLzeAXKwkvBdSI9zVymnhxr5qGYwinPN6lmCKol
8kraZY2PqfHuX/MYYd1jMoa5Bkp7B9I/hq/beGTaCbSLtLsQT8rmxa58j6D8tto7
wQKVcJMkm0BcOwKo0aLoSlfT1gf263lD1PcRj/9/p51kDFNW8SFqYnouHW3WccSM
qJRufQBfoaCbRkuh+ZcXZdRbeBp5Hnpb4XsWqF2T9KlDirlwZuwfysjzTIk9mq6I
Qev+WtzeBIFCq9bn9RUP2tSHYF/VD22XdXUF1yVnzcbRtnenmB0qkL+y2+oP1uY8
zO26U+N38MvORlTCXv+pTctWCzMq6YRNXfhb0b+VveJfSDkd6nZGbBvl88eOiEvG
hxSJKwJEm1AC+iSxDp//Uqbx/8TW9A98oGyDP0lk+ztShAl4/lOOC6eFj4Gg+PAP
wJG2ZaaxF3yVZWCvH+qU5cWCNmKhd0MXvx1eLaGhe0GmLt9+3V3vrCDzCQdUDmRH
H9BamRZB3wStOHXRHya95HJp233/4s0l4k+hUfSXzeHdE9O0JhD/ATZcwdfeKV1q
LLhjQ/XHdV9LaAiSTYQd1oJu/0gsKRfxHUzuA1v0LKcIvBw45X23vKQJtvp1L6Te
Y3Z4I/d3XaSXsA7l3Fub5Rru0FAxbAQ3bVcGYGoQQIWR1DfWqcd8eBauY55884tV
21wzkaFYMOhrIkqAoi0JDU29EHPADOPKOM/WAP0l4L9jbXYAotG2sC+wmALFc3UW
dA/8F5QAFWIzkTjOUwaVVBoq7bMW8IMU3LrIYci8dUokaSDr9692nvpcnJ2/NZG2
fj3AW70RhAeKc4fMTt3TmP7a+UjWGD04JY40492JllaPML4tJznrssEjreoHpgfc
9kajlQZp6rgt/KzC8vUbIWq1umGJ3ivN7PuFkiA/xVgcPtzHEr7Q4hhWS6BkStro
I5rFY1MqyyBMIqNCMAT5TmYricbGMEWymWhP5umilIgmYA1csgoa072ndKihVHHz
tQ3KGPIJWc/Uq9iSJ2sQHD/ai0ciOJgPIzZIv1Rgx+UgDNqQo1tseSFpz1pQC5IT
cjmkBEtX/kcwOxYWUqOmEns1wD/rmY5puNEKUVlN5tsmh51X05QEgKk1rWyhIU6g
vbCBLvr2QZ80OQf2FftIkvR9C5axrFhYmX2KZdfE2Fou7kfZCnk0geb2BchfMzU0
0ntnA4d3phIlP3194HRAA3sD77qDblNxGmutdMxtwbp40HhXcM7KA1/wc2X9XzST
9co7Z4pudT0ihEvsHkr7ZAVdXHYHn4q5HEV9c8eyaS7OKoXeq+Keje5TReH2htAw
I2sKByooCl1AiczQ7hFMzS0DImNysyjqjIiXmBDGIvfI8EBOMN/0RVVldEX3kXSq
VkP60yevIevWabLPi6sYletipdT23Dns3BVkVY+qC/9Ckb4UGVPfTwdacYHnqgQW
m7sJHMg+gr5LGYfgcNYL0hL5FZkjdodVRqLL2NbG9yERscjsQ9WFctnjmYrJ9FnA
fuGZOufUQP96S70fZ80LE/ncGq8iGPwepUJeCGwSsRYQ1VXRlCnC/11quHd1EESI
T3caB4XgIQncxD/FTNclX39wn3lSpWlA0NiLby4laT1Ql8LMTOXQvhOMgO0IxZpl
ulZ3HZ0Nf9pkYQ2we/wYzeeBJQsXSDzLd8OdljLU7vBOV9UBqkBo1jwHmpWxcPtO
2v+3ySISD8l9jPwctmgXEdAdnzOlot1RrTLkqJYngJUrwX++NVtwLst+9LYPaKfM
sqUtnLd+pNXwECW0Rkg6+yNNdHN0Wr1srOD2AM35S2RkulLAv7Y0bFPHfa/V+a5x
OXxQv/+IzqE4G90otTaocRpIms1roPa5r6Pc2UlKpHTJqOTIK1byw0v1+i9yhAbe
qsD8n2zxxk2h346TZC0tfSRlgkbnsQzKMoE2tzhuRmVDqZ/ZncGsTtNDI/J+KepN
I+Eirp9/7FVtNm0QW7Gc/bOsbsaeR0AjKxcJAvZkdnXkwqP0hGSwGHc4DpImR6T1
Re27lca6ps/pbRd/Yn7vns7ZF00PHOLB8XF2sNfJTTr5KxPwcygRq1vjemEfcLT0
D1a2/8bj1meEXaVeP8kf63deKjvBL5kicPyK3Sa9o8wTI8NkjVNAkTCjAOBG59gi
qE2JW3lXC/fSLbaRe9vNRvK5RonpQMqTyZzh3j98OE/q6oT/Fn7RTZWSbiAeBn08
PXzn0O7i3Vp9nGpnBmNNUBei2EX7gjgmPvYyUtkynWjKfFZVIfOc0tVVMHxWl/cT
EDbPB7W/aqDhT3SuuD/OrWXirHwzYMOIqNEz+ySHVjf0QjI0+9QV7XnUFyXwysRn
Z1IZSMliVyzXCSr6e8PQRi8Pi8SMK7oS+jbqcCuEQh9WkbJCTkMz8Eyq729d/nRZ
ZUhbnMcwBT+uhsyqGeNKPzrmUPcy1Piz2WB/4sPCmflUcqAamldEubeVsw4axgSi
xgAMoU5CXtYFEz/MekQ+ZHllAukt6KNfZeSBLergfHCq0LnqwfZodkXTuaxF3JzO
7mHFGLKJrLHZH8Vsssexpaw+rRNzpS6TkpVYlq95tFU8XovqyJeCyHIhqnog2O1L
xKlIoEwh7hMsz8Rjc4iGwDGadSyIgc5B50yFmftW0DwPccD3szyVEErMyGcn9uLg
Hjh4JYSRxMLxf1dP5rlu/L6IUhapfKzHZ+yE7bRa3HyXF2SJmZ5OYrKBmARcGTn5
XpyhorUh0tx4Z9x+FZ6MxvImup5xXoWvAXZoS7S0i79/9FoX95RSKZz08B7mysnc
+WOg6U/w5O3Jy3CaihzCbrbsPDVYa6TBAzJL7F3sGLvfc15bgIW0ogzY/K1+MF8S
hqr3CK60kIGfpKAX/Mmmt8nXF23VsNB0kSFvqGHGrGajhVAGpzRE7rrFs+zUAmLk
FwOouvcCkyzzZpQofx03aXDwm8RHxDC2i8vf7laBQsINMN43IWd3tLAZumTRaF7C
xynOPTHgZl1DF0kl9ZFIMsW2A1EV2lWq41whF6kYKYBbftewia/G0kVgrRk9hHSF
ww+E5lWxXOIcaretkllM0VDgFk3YasiqeInL3TO6SzNf+WNUHLYHJY0GPCjXSzCh
C+F9tBbLYnED2dus2LkT5eiJr2w+HtRa92dG1f+HGYLc467CdYrXzss39uyMs5mS
HE3GLNbKZrsl6Mm0r3O+PnAkIjCiyTPQ0n3mMWRwO2yi/ha5DzaIbU84Of49NMY6
v6I16Y8Xq0kpymXxEfCOOIyWK8VSwdjsRxPOp1rwM+HOrT0kQeN1ArdUWVjTwXZq
44u504+VxgALYACOra48OVY0uSSYoeRgh3C2z78GQJXL72QvhWyRFJcigq1b5q4J
AIbN4TIuVvcYKLwRzG+tHrwE2VU8T/ioG5pbH2sU+xDSOQv7XvWGxEJ7dzEl7+Ag
mv0WDg6sgl9P8keVL4VljHzD8GhuuR9JyvBuZs0jRlzwmx91qLUvNYNxelxHwrJf
2uJVi5g5z0Lea62F4WXKT0btI251Cqj09juOvbrAJiu1aau249sHRyVNOE5rw5O2
zJ+c445vSIiXJLAgD2cgmMQ8Y8uleLa1p4mfANHbE8/W7A8gfuJRYKn1wS+CKyMy
vatTpfbUS79uGgdQf/de1LtIWQGXdHvZsWcfcDnnuz0R4wU5psMbE+QZpKOELro4
T2eFFXbbv89FAXS/xTAIRSGdCJTFqC9WXJH+seedHVrPAlkFZ+qt1hEqKJ8zPu40
c7A5IHSa2aCMKD3KjxoaIEaw//XWKjkcDyse55RUCg4r0wMSPZOQZuprZVCyMHdu
xhKTulLSKSXEs51NPGKFi8Z55a+b8jDdfcZlfSYMc7aMwEG7OGbPG01DOytBLuVY
SkUWaiPp9/EI45w3ibvaP+SpHcSt0jDijRRO4GwIE46tcBxzyNGyAhczjEkaNfWB
/gBjF+cRsDbzNOopbNGb7fj0BUqaMx5oDZNDCwex1ipCHT5DOJ3hrS6mpYaA/wSU
eug5G3lFAVxsmBpTdTuJjBWMf3/2hF1XNv0gC2QMMgePelfkhS+EKAj7RYbFBFo8
dOORj9B7BRt2s0royBxG5W5f/U7hISVwxv6/tGOyJGsVCagTyGpVwkiXcVsWrCdT
fivnQoHrDbswdtn1W7GaxDg47z1dSVIZud0Y32usnVWQUZYIwn72dhkD6X7IUWS+
BRfTBT2VbLPZcQyZhMDZP+zOCYVXoOX72QGPlIiTfqc9nzFLcwM80QwYl80g3vvz
JDj/jE9huZAcg4vr15rjNk9AhwGRQicwXqPl0cVqjUW/cq6f6oQ1TzlzwgL9FuLs
2l18okH7AHv0Yj45WyC+YrcwCZz31+E8EXp3isVxpLoQTMZnP89P9M7cd9Msc9xM
uUwYsuXBJpgXDIRoetno6FIjBqzq3tquwqmRZJcNIiTe5RObRg5ta+lAoiI1qeKR
1unWmKa5rBKXTyf5XB2MtWvdmPAoHj3ErB6N2d8UKmxvDUngJvUj8bf7EMsYtAr5
DWHuDg/4++CdZU6EW/DP547obG98aGky5NyDH+sqqRR4YJK5/pSJAhEqldk8d3ri
aFx1CKG4679goM3j9DpjSCcXoMKWDQcptOR2fYUnRAMTKyTsFVRBQcVzbmmJhrZA
rtZo6r9cGdqrRHlTZoaSTN6qd+OD9YMAusCTzu5cO70bNVqrVpg/h3mQQKdnfGde
DVBveZWiqmtcFAT7t12nWR0Qwd0qLdA13KQdD0lgdgX6WcSJ3gk1/4lULV9CxpqJ
0USYZMkkcDOXmmDma3FgKoNZL9kso5+2clIIJvrfRN/rVE6bA6uya8YK9UKwlsl6
0cSELDqbP29k7/VvgQi8t2XF1PIf5FjU1B866Rcd+8eO6SkQO1ei1waZC+1IX19b
VcncGw5er/xYXvwOqdFIPTbTNvx9ddHkMCixuJw2TBSzDR26Q6JH1k6Y6kWXWlWr
vKvxzPQ5QpwEdu1O7LSIYLICNIP00f4R97tKzDqmL9SUugCYk0xK1OLuJsu13DAU
S+XLYVQtqt0jO8OWSOtMv6qQc+f+Q0hOt6liU3YnaBVo/I/1tb+mVa74tJd9oUrL
cWU/B9Hxg+9A4dkdIv50TcBadAG59iYbHF3b8wkD74ex5mj9CVPA9O7CaFcz0Rj4
oBK539AP5vz3f92dRQANuSX6npWwhdz5xMBFFbMIXtXG6/BLTZJTV0QPJmRW+A7C
OP7cdsWus8kJRJZS8GWARWfm/zE6WEgVR/m+JPV8QYbIrm3blgr9S4nrt4kPXUrn
LjRdjJIacUJn9sG5Xs/vdWVvwwah5ggHxuGDPfjcgoJZMkLUK2bS5Ltzfm8rWgPl
+5jUY7XDyk/65aqdbT/2S/Mwmyc7oobooxOcSlxip81F+AskB7kYXnTe1adX7gY7
Ot7nHx0Y+Wmiy8Eopo6QCklfSTR7VOnk5oSDDpvfUrVjZ7LVn0ExYG+u4Xp0SWe5
AyLEH5MZZ/Ebdyj22aK6BmJKvE+qCwwZ2k4ypeoV/R7UDdIDl8Oxu7HjE6OxBNaq
ZeRbL1p5GjtEWefftrXGmnaHIFd6l0ibeR0ltxilWpvnIOQBwHMhNGFCCy3c/GWV
+dbLP486R3R0y8vR2YFelXDpk+Jfg12AXGV+yRB2H9yaJCaBf9NKqWWb7CN6m0W3
vWns38T5dxuhKxa0JbPZgXEyprTBAqbVG8FqRcxlmt5RLmKliA5rJEpF53LDLalQ
XKDQN3liy+qk95k/EVxc3ctvyR16EO5xIVRUdC7otJGpZGhzJUnbiGAIRzfcGQIK
S4D/7iKlaMTHDddaZ5dV79sSujm3t7BTXknmaOL84Qg6nbgB8rqiWdtE164S9w0j
4G+R2yQj3nTANwcTatGC3saxZ89TiDvqw/7PFxHdEAGFvNMa3cwsf9ZWAGxSW5XG
AZIkPX5txCbVIfzcj6N5KTLjS5cIlLjdmTcZIksYcoQU2YfkNsFJpDfoI3D2wWNF
+zF4Ahcmyso2Maxyq7PjJYdSCK6ttGprUZJQW/kdDKdFqkCuNBCLXeqpte8tT1YJ
oup9ne1WDSnQY/b+i6p9pGDGHKUgGY8fnOkycvoXl35KHsHT5cVLtJ6euOEYaNti
Dv3qK2lKkJfcFT9i+XQLAHuuIZHeuxJG1appTbddKYC3X/o6+MA0jve/0qKTkag+
17nO6+7IshXEiDI+R1VqRPZujlz9oq5LQJEZd1b8oHBXGflALE5TBsFGuU9EP1q9
4U5M48uQtEjtg+PH7EVyCQmK88aEhudFttJ/STOkKKmIuPUn61cFsA9X8ukfzDEg
W3U3QfL2tZZe4AKnRooxdSnXzcl4UiMxwvXWLhby/Q9+sbyTSHx3Y2U7CSOwzyoX
Dvzx61MmS82+nywOZXUobxfsDwlmVKdYW956avn88dpnUMkBXXNN6Nie9Q1UgssB
LHo0qB0vM7xNSrkXiWyTQiBHSh/SVurf4TzZjB8eeZhjYLwQNOXIMwRspMJmi0Y7
S8h4n3qXVQvKT2DTtJ2NjAQmLxAMgK4s13zG7iNfx8Kjywj/2J4fckFxx3m/QIt6
flkNJRHtyjMZXlyy7MzYSJR2n4sZ9ZyCK+607TLmntVbY2vPyLrLzC5b+6LgBP+x
Em4yXTBYlzh7vrwybFrTC1brqUT8uWrdMTOd6XC21eD3gGqm73MHUabULTyGRGKo
LWplQe7r7d/jfdIaJzuGaWlKLDMJMqsHGu1PlifPtTU2LBCJuxFMyOlLhdqAy7uP
X78VZlq2YXMlB4HTff3hMUVJU7sRr6J1bKzjKS8sqyzzTI1rPxR9MEjCjXxUT8KA
45YTHHn7DpwJH5TlIgqAQNLPaMQW8BqPsRjAajgjJrJiBScdSnshP4v/ESIjqGi3
ThRZAGu2rRiH4pg9uXEMEmF1h24og0Gio2FP7jW6tldu+vYCxZVs1XrDCOuSV3uw
Bvmuf3liP7Fsay9n/juUbJCrHilyYFV62jazNWId3R5+OZlRTiPgLZTaNa9UiYvQ
+Gtg3pbUwr4fvimArYRIw4jmLZHe8s8t1t2NNN5pPrcXdY8VoundvFwIqriZrHYA
79XraWESiU4Lxm1/EjbQYAn8e0zBr6AmzM1KtYic4j2zgmuuPpwQvKnBCn9J2TxR
/BCsjErUoU+EBQ++X7uMoFiCM/0lSf9OR42OFDP1Wh5YFTEmV0ScWRi5E946KvYD
wLaSWYsY2aaG+Y95GIMq+ye6ZrNmoqOa8CdLz5N5pE47B9eR+RyXatz3b6Uaj1jG
h2DCTEXRcvyTkvoUivMC7LUNi6gslhQ7PmXDUyYvwhFmff7G1EtYlf1QMoSUKCYj
pn9pOAJOztmhruFWQeaE24jcFW2BkJRmbw8Yu7rzH/3AjI4oymuU5KcYDg7AJdh+
WTUHQX+f+B+cUUX1XLz5pRPCqztesa0+GZEpJT6MmNLvnOL2TUgqe+S+4zoRJugP
d/uPVa6c5+qqkIRiQsIEDgQbp6WekXhETXkp1GC05ZuDirrbl7WWrjIePnLUNiRM
fMMfLhSGq1ukVIZ6NO861llULYNuqnsa1UYoTzjSiQigk2pt74Fso+mHAmjHlnWE
g5bhq7ZSJ4GAkCOH6vcCsVk4CAiS48xLjEtNjxUVkGG6FRdlJQ47K9fLQBCngP2q
ZVPWUbh/yX7SDFyVsx9d+0lIxMmcmOV3r662PQySpuv0kiHogxA/abNKi7L1h9m/
g0Kix0ZfWAkIPhQGwdDzIzTVpN/mBF0biHdcqfvnGcb0mZ+OSWTOD3V8BOGv1ydE
qQsUT49ASedasYMkh5uAPADh8iTvCgzOYJ4mWUrOos2zgceNA5KG1uY9HfD6MSuB
65nH7yQDQhHSyai8KvowVRjBHpZkBrhB+qWgC5RpU2dhRQE4KS6w0R8t3aO8eogL
MyjCRZ+LzgwqA/qz/Pm+jLeoBtyJEaTePGDAkgEyKN1YNVnRiqGl9+IDdrH/bfrg
y0kCO3avTLC4SeWiercTrRtPaG305GWob0MNLXnVlwevY6De5JeAbGlCc4h2txWU
w1Q8OxLQ1Ccn5ffEgR5ej4d3J2pRFhcNwlYGcWm03r2n1ull23tb/felA8zAubNe
yiSnOkeFsYtdLoJDzLkNSPlukYEF4PQvH90afXcNE0jZp16YbIbs4D6ou2nGz5hn
qOJcgIPvMns5LImUXQGZdekUxyBP16t8gubqx/+u6ORq/mwLxiuhZI+L4vexR51C
PRpOUnnkNVsnb73fPN198zKncKwqZHhMycaHi8hiOLMhBRQLnlP6fe4C/nau1N4X
wWyMqNZmJhn+rZJ9xWGyC/35R8Vnuuyfwov2BddDcziLYza/HRbE0iTfZCOzGisz
ht3IpEReoAJBZlm6/0sCMHpkvBPa9OpVrqkP2z6YuCMEJdYOnhZpLIVp+QSSlyZW
bIiHZ55EM6UNPYDJcyVIJ8l6rJpLynSsNRuHnGEV6AXwBa9itU+7qHeZffhBaNhq
TTOQY9YQ5D4k4DYn7WNGhRm06YQfQQuTRRzRwSfuOyQzk9YvkEHugE5wDgsdtpXO
HLglLEQj+wrs3xhKsoKZT4p0AjHME8cSSqMe/4Z1JM+7JH6c1RrGk/gw3+//33vx
j1/XvoXlfP3/Py+frZP+N8LpM/4Lq1aqll09x9qJVMrgCiQPNhiOClDm5ydyUPJS
c+08UjKqUDAs1D2NAUXPdfgl1uxQhbvNupjmd3A8+vxIk7cz0GwA7xwji5eGh50x
aPxkiFO9LXP4PDqiPWRA9eRh77wvT8QrEvxsQzirFCoM3FymclEOQ4QlsneUr0v8
YswHNAKzoZeOE06AQ/jaj3slQMJsFi0UPWitZjUuSwOrNPz2TqZ44pWltNbcxy0r
rX/bvWie1F+YkoV3qg+5lP7IDTRUha7HKL8m6z4ZEi2PqQtM4JDhXvF5KFjdB678
0jSAtiJmPwSl8bksF2kf5qUon25Ky3yYsil+J9iNQtcsOuqQWk0tVgLPbF45vAos
1PyDc34JvDqOKxYQV2jQfjBWdfV0+0NBvpnda8r9y1bhPBQ0LlN0BAVBzKzIS9u0
LzRqmlLyqvIMz1/GIPKjct2lGyrOkZaTx9Lfo4u95QgI2fzWqgsyTEJLI3Snhhf8
SPBgukTssql6liGC2ZqOMX1qx5vlZOfqe2hR/juDt79MdFVIIGIq4sSgD5hg/wEl
IbKJ9ucbqm/iCeE+f3LRcJW4twrHWfBe3UCv+zhrdw/GdhWeNKxzLqNX1N49aUII
++UCNkOg6sAU/bZ8GHEKvEtVwNrymSg+zAFJoYe0IqGW3UDARZv2UXbSB5TBDd9Y
1Uq8u5h9q4KWwkqxM9DcgJHh3pt+hJAVK/7Ys9WTBJiyiZGKLff0mMnCLAvMjKXm
zOAAISyxzpG28eMhLPyTcZkWlN6k75apwGPPRtmN97AgGhcRi1yzFkYzDfJamgtw
QBGE8J3WoV1V0wQRec3tgTNzuTNxKRUP0s1jY4kSZKgvlRmy54sKh/LYyohnC9Jt
ZmTCk9TOmwK0/ep63qbU2Eka7wmAtx9Xzv+UoAVYWawXuBbjzfOQysgjaEy0Limn
Ity1+esidwnJUkIZDBpPDLK9GW5KDar0UPRsZaGHoeN99mfYNcQv1U0E2jW98XNL
aGZmHeALIIqC60GNNdTX4ScsxCxbkXa/s1UGpVe6hxxb6CazsAoXj9g9EyIf2MG2
LyZM9fMWuJMlg+ZFrRSUEkTY3E0ariU4JRe95yE3i4etgKFyPvnpVpScxtRqJzMs
djAvIIyz8YqWxNv/Hq//pVu7ahSfwVMExThF/rcziblioZHLg6Z+iEs0r4AIS3nL
TrRRmAOU7CcUooe3Ban8giWhKe2cusa4N0oeJTqhLZQw8Xfz0tKxScE6LweJu4cJ
G3PnZ6jM2vVAjfk6OGFufA+z0TREvd5CwirAWMC/sDQWnfKiMaha8eHuCB3ow6+m
l6u00vKmokkExatOYEHRh6NrWXNsPNojiDW0PvjPs56/tLxhmPPRgWUaq3xRwG7K
ECI30ac9XVFumndE0CNWLa8CBtm8o/U/EU7zvjglg/0nGorc/vVrICAXrob1kafX
4f1mucJsZqdhtxlMWkaWFEXnGz7ig8yyX6TKhngNZHOQgJKqyOXhUJPwSHQltKTg
0K0lWFXauvCLXfyiNpPug3XrNY8pPCd/eDRqVNEmFiHmg+RREtkl/298gLI2idFX
c6ZuPZofZuUiHuRZ1T/ZjXc8mhb858uXurpqzUcfgf3hSeDgWHfbWHqrkT8Qx2uF
67drspBVqOWLzk+h6LAzHEVbQCWZIO/oNXetaQRsyKNxIHYiC4+m56YY/Q4Q7+tW
9ZpHDtzqvPyHEdc/upZeg3DA7Jjn0VOYMuma6to91qz+CVTCC22Q/QrjlP645by7
mhagsrD/RmiKGWwghfCpE0L6tKcdzA5/7RVOu3Y+bGhbWHA5EOoy8dfGcCcedX1d
JNoy1uEbK/FIpiXB0W07cUu7hyh+sJxfpJSohmfifCouLrmCBxO3MvAsPKKSbYEE
tI71KLEda1dxLaoXyrQoRZU8MB3+Ug2TH9CTFzNqE0aV2EhcbFZ2w/p4Etf8XHGn
2DeYqfiYxzPzK/TmjuzewqKzu/YMGBl8NzXkw/RieJchD4oVXc5c5lHBqPGN46mR
HLKvqYLvI3AWtTna66eBhYoeDHtxhImV9OMdQlVXS1SKfjAE6VCt4vigI1xlkonO
kR28grrQ5cYBFmw9ayMIwzWIwFZyG2NNcvc6TxvOu/xDJi2JsO3vj0VwT93wCiH9
NEu9Aku2wniWC10nP7SEOZG78aFc8udTQH4VQcdtjU5airdbonbeX8oHOlIjT1Gf
yZ6x8cuWv1t6zlNGhRQvUeA4P8ETXumQR2yhPb4mhh4i05yBoOCSiYP2Y5OLkU8H
gwcZD6K2+TYnBZyTvw9RVFfjLfPevLONWxfVo9vPjZ1ZI3scBmz5wvY9qWIs1qRu
HbTLLlVyAPBab6q5iX5X4zLZUHTUUvr2JfnYgk6UwrzMIKV+9SSfFUkl76mPfxpZ
opHb/8M0enuX77pTfowVaJumr/m0s0U1NjTBDMD/iwMQIRWZyTiXUA4AOsPtsNtj
4ckP4YB0EjL8pugr6SsGrQrhV4sucEPG9TwxRlCENXNRrtGU6g9/63POK806BehN
Ua8oEIQRdnlldyKe6dg04zqEtC+iRatuWnmk5uy15K6Vz44vm3ybmnxIE3wqmvRc
lEvKRlNiEUXTE/gn4l2/Il2okq/+gWszvwluAHCxj2ktN1MA39RQ4RxEw4phcgGb
xoJzECVYsyCnCjxv8T9v7IMXqYk76E0qsJ2zWZ8y4nu74/3ykihI8frX+rdycfUq
0LGADNiZ9jOCLLSPEHu/ZBTTFlm2kfh8+g3HQ91/gmfawq6pKUvmUlu9CDMyH2jS
bVEmJgQofKLN4Xh4JxW5TvlaSbkDpxbOwsSmtyvD3VTeeyk6hkXRZUqFrxCwpDkg
Wx7OHruXRXHQ7x1jhQxVtaXsshML8JpI1XZQiOOwZIjNDEpbvH93HmLvifajY0sP
0uIPMtTZn5/MyQf7zt+KojOOs10vgWIVSC7fOQ4uonegS9hHFFw4MACBW2XNGfBh
C7VlpksFr7KadOyiyUE2Jv0Sgo7kNbjeNc3cWH9otFax3BPvTUH9+WVmheHgy2Qq
+twq8T5lIi8oO5K8mhcVOsxoGtRA1Qx3d7hF994E24IPRMLHwINuQvN56Z7TPykt
bfSCkdgihbWMNONygJxItdHWJkpvkuMEe0U5VqUZ3TmdxIYRdjIlUuxmFwTkpRCV
OztF4qVH9pe1MZrfcgUBw4XXyhx7vJ3vK2E4uuIGGuvTYVn2wFVkVf5buv+RHLRS
WU5m9ok+KWlvisYzyAfTyEM/gr70SDaGdPVf0Oxd+wRWcfSdMyegR8Grw8KuXkVr
I+Y/3lZc4rLT7T4wQ/aI46bLOUnSCCi/c7dd2YI2lCO66GBQ1MmD9WgRAprMkLR0
gj2ZB5EH00n5CBw8gKcp/uIbSud7NWXv1Bzzh+vWaJdW7r5dHWYK8I3fRRHmyv2V
WM1i8r8wlVpdOTlFlDSanpI99NU18shhwQZBCTqXEZpf1CB0tzN9AConx4QBlvI3
aUrG5+NPSOO9JRZl50vdO23EXi3LJTOxVaNBgry66hNW9yaUWDfQJVrmzpELDNM3
KydrmjKGsEH/IHboHMDe6KkPKHWXFw+vly17sfR4Lcb5gR82vwz7rFuvFBF1o3rt
AY5gJoh2Y9YKdYhvRh08Y8vuKmsw/WQoFIm1vRjsgJRsHzxdQFkRuXym5Nja0Xc6
CmjaAOM5URhCgiIVwy+Cg0Hftf4Z4deJPWDG03kDVsKKk6utoo4mR9z/p5UmEPBe
5EUW7ZfiGQYXPSsj8aHq3wQFMpVRDjPSkFqHes8T3jaowp1IsZq85mCEUv81qHrD
bptMaOZIxFDQzx7IE2ilWV8gMyHLJuFTCPeu0zTSJPhVB1fQkBrscTzJV5GgHwon
DDMvw+Gj3aGEELBMnTDC5gxdu4pV65mgYkU9VzgLv4lAjLJen10THGwaCWmEwfAn
u9i2Xo5Jhu3Lyx29eJlV5iOV2/S4tcF6JV77Ncx6Ae6aD+hQt2YggTbqUWYOGUbi
b3L3J8OQeWWCf3/MwQh1Gyx7nI+hkHX8RNRcfGCHdCx1oqOdlhvB0hFvB1fqn3mR
2junBs4mV+/dFO962GvlvyOjthWyIqtY3+XtVcs1V5aueQiO5UDvLhxatQJFKKDp
pGyQi0Xb+i7f9uvq3vYpzwcsvKz734ts+sPxLkbsMwIftLFe5QFZQooWe9sBySgK
Y5tZDBIP8p58VxuwsIgHYiTC9WSsk6up2TxbboD7sWNf8dwTh/zlmNwz0FOaG9QL
u/8rg1izdMF/ATue4YMjfErTn14Y9a4VXC88i3tZDOHLq9r4w5VUh99R5dEuBMwT
EpqCC+u37H9rvJ1NKGJJPTH1VGKXCfmwfRB8iu8OMvCA08VOHT4NObFB/4/T22Iz
M8q7XQn7OBGs58BlV36B089qvv0XmLZBKE/LKGpn6GI8QgsyfSafLydyx7C1Olt0
MWk6d71wr4hgZ41iLrhA631mFC4w+VE3cpzhO+coZgOtnkq7A+nH8/eaUOrmmdmN
0RLReM6FbyRPZF2M9UYqiubVYU/W8IAylVHwoT4h68udcxHc+HEbhTdj+REyh7jc
oWxqkdrfO20HQkLK+ZpTCq9TRe8XDJ/wYC8rAN4cNYSh8EP13TxJnoF9qtzgcHVZ
VF0rbY6nYuAJqk732GZZvrmDn2FmAF7I6Fgu71iC72vmvrxaXO1BmbxACoUlRn5M
2eh7hoLGbBl0vFX7WSYWbKAnUzRU7Mudthg3kUSoi9qa12DxrUSkd6Myvy3NV25S
X2MsH5Jxe84OE7jpPn3134KVIsHfP8bGYzUa2zRBrzcTgjJgWNE+dWVp/vYMryC8
vUT0P8zqSoMqgYyMonoq7Rxb0IdDLPH1y83eGaP6KBWfDpyESdeTBTiG+jT8EA21
YrJgE1VFkaBNgGJ1055U2mP2mwwA9EX/I1pqfaeiJzUM57TWMxoOgjs3CibNh4Oo
tWAcJyOUPN5rbH5irFcKjzHiStQ8i2q22sl1hJJbFRfp4bCe2jBUcGoO0GLaZ+sP
JLCsdNhVfp4khknpQxVsN92utAebq5OaU4rQf5iUPFwugam5RmD3v+VQD6W4mGYh
S4xYziBBZW3WXOrCMtSt2X3L0Ld1FKd4o210skHe5YScH0rwoapFj+Y/gVsl/srP
GhMmZQLTX9IwabQn75JTYqETldm+d0K078YZQc/ynjjTXhtJ6G50l1YqekRCk6aR
Yv1UVrSUjE4kJoQgPNjeDDin8Jm06youChq2R6ErWmeArQmMigou9BpLJL8RG+Ix
Ky7qydC0JThbFHS+V3ydlW/eurbfYDBWJceYCndB4aiP+ySMcMTX1hPQsZcIAaTQ
D0w5KFXv8cJx86mkG2Haa+MKj5Z16L0V7WpL+EkLhksD2/n1J1T+d+yo3OizySIX
4UHK5bfI1xjmdLcRZGk9ZDtVWlPcflsQDYejiJqzNmy0AvE+/PCi4l0ZY8xOZldq
K9vSqnhED6EToa+TIXHns945cglAZ0ov5asFcsxSB9kea6BWrKR3ifA7yoS1tIIq
U8Gh6cWGE3/O5yPsHErqJ4Hx6cTuZL7tCMMvYtxFP661hbTbntjcN9n42xP2HNvj
JXQkFgm/Wx6vptCav32ieJJpDx+0Z3gl23q3r2ki6P96lz9V+d0E/zAtfWITewzZ
aRm+dUyeVQT6W5YWxJBxNpxo/I7P3etAetbDLg95C71XbHeG2yjI8WRfVW8Wa9z6
gjKTOSLPRUirF/j4q6om6SudP3Wq7hNerL2Ocei8g82YaTksEAcyQ90jpOFeCzUy
l6zUDWDXc7i+QITtzsh/5JamIviXpQ07vKI26N/op+S2+zJQKGqfTE42yHzG6Pkw
PsG77ikANwrvOKrrnW4+qIZGC1vQw0memjy6IrpVIg5nuXGzwkYSQJoCE98C1+Oc
QEGbe77BJr3MDQ5x693Sh5oQxsvfdbevKUHCIMLfE9xNnrvnt3OQk1ioj30RRTMV
1NpZAG/XAahjHRhBV6FAGxRSUbNVE4Uo8m4+zIQpMIq2uTP/h/cJhlD+7At8sH2G
LfFFgoO6aKmG1WkDqRf2ChivW6c0J/bKUQBppKzd9veR1I6BvwzmqpH1Qm5iesK9
RouFN55k9VGdZhv7eekZAdI8HSNM6V/DWG+nlcIKzlYvfI7TmRZOz9NnL+MMiOoB
Cwlyi9+P+m6Cib1KIUheFafiPmjQ/EK7tGwbR/WYyDKxn3GCe2nXZqfcvjXFUQMF
l7OuHLaMhUA4bpWeMJgIMP26+T4yRO+bOiYpMMQqAxB//2GqBBqccZfHjL3MwA9A
MCcghFEe6Aq6EQc558BDzx98QeTKi16FZVUiAY+ynFSXr3ohxYWokom2lswYI5MV
iCP9TV2y5Vv+f4eyLQGP9SNxGVgRR5zxyJVGM6NjPFjyBULaYvoqgDzgi9ogZTll
bPR/xMTNXK4bj1oS3fgdLF8M1qbiBsXPprxsmhdNy1T+2ZEcePU9hbz8K6SCnWzt
FwhKmk85MZnOoRs8UKTPzSpkiQaCT8FN/289an5RNWWKxEyX2FIxlu5zo4ic8v/O
cPGmvBgaVJZEt6/sVuQqYXLkl4EmZkv1mV6SFnuafVuVsgSkMIOn1+QKmXgP9u3Q
5Fw3nVo/HfU4pGWS/nxZxsiaqNJgTzzhEsyzAYKipH02zsIUTLqO9Vuc0EECCWQu
FXdRJ3jzsOjXZhNRf6423NxWGynKZc3R9eFCYBrixv0fVmvMAqZqOHkniGeKY6pk
7nObR+o/X4FtjV/sg4n3ZSLiSQsuNFpE8XJZqcZtQ3RGLIcvtPALKmU3PUQuRBj7
4dCvF34obH/of3OcnuwcoO6LeL1aByi6H00/A8VZ7fzq/UaGJ3623CIYmvZWKXlZ
E5SLGDtNN82YPviIxLqx/bpD9I5BD6G+lIMYwuMUH2W9G9TyyogxIKS+P7KBkIER
EBY3UvkLl8xMgRCCaX3PYAtTcM6IegtZxRIhtBdDgdvqXRfv1yyu+DryqHlrdycb
STIIJsqGcgcEqrEmTXH6aB5nxM2FkYurfDpAxt+uFTQ7EYiMjrG7JTMx+ZBcI4Ui
c9xWGd4DjDOuffNVw2rM9kEdo8wIUuXQ3Z0U+pJK0A206tUkP67tKZZgoerPzALu
9RWt+blYSGSLO+DUSZ0wSwKATqgR42paCb6biWzNUz9IdpUP0YZu1N4igLs3rXdk
de4Or/F6aay9FXvCgxUHhuOWyo8yy09U+Ht18Sg6Vd/62+X+csf++sHVd6a+Gpys
5gdQXa0t5tKY6XDBRIFlyAnDHrxa98NO3OeOVflpM1AJ1mDIf4b13LyExQ+HeRI/
1pIWAevVdsqxJ3z47R4/CYK3rs6lcisGjxLJfaG3at6wyCs+cGl2ogiFRK1ck5V9
/FBbYARAVaAfGP4UDpv+/t1E6AuTFRraehudeRZCSIWLLpVk4mGZ/R7gEAY2eSzW
8LIarqzXHa/dargQjZRv/ilOVuqkEzomGzXajWppiAYlbg5fsLfscQiJhjHTmKxc
ZpxEXkEd6zqL3Hnl81I6zejAOTjwIqWoXM447V2tzPBm08pgix/ev5jprET+y6jZ
Ix4Pm6ajZS+jBDgSZXtAVaadRWrzZzhAl84A+VdNn9dgFn+qPztHHRIsDQlkIKE5
3rVupqRf3GTQqcsWo7dZH7b5XBo7ueupJX3GczgBQz46wnHepu22zX2hrJ3ytA+a
FF/yAQ3Hm8DF0R9rpCmNRZR9MJDJnzzJLAaRuiSMZ8pWOmd4/xM1I2kzWMIlYCLb
0i7IeAAVf4SrjL+LBAchoctGoHTzXvewp8peoDZuydAmVR2AAh81ZBFixAGCFS/0
XL50lTT9FbPcx5ML+QOlvH045CzvfiOYi560jxlulCAPx0Rl1a7EZucCmR1HNZQw
gqj1r1QqObGLaRy+0wq3dMVqloBV1nFXLb0mszGFTcCkKS61v9urOHr63ul2z61M
QUtLVTzWV6I2KA9p8Lo1cxpPZ1swBt3cMq1/hqCyrQ9+SGXodgODK/T8iLs2Rl4D
zT1TQxZ6x/lcb2zP/LISuix2ckYnJXwYfPjVrHmR5CpThMkhGkvM5yfkhPnrGy5y
DTOpouKaDYFPxfdevGobpCKqXgPrNwJr/gPVVpXwqf1T/BqCkSMfA0KwNuvvDxO7
mWOHpEClRNFFEeGHQUbY6gcPj6m+JVRTmraw/fUXYKGkzRaQyaRngZQPdMI77UpZ
JmC6g29Rtm04r8UZ2MYBRwtP6/BUNj9AuyQm0EiAkqFfNQZrnNSChwPkXoe5q1fW
Q5UIirboy8iMECBVc91b9pEUqp3TFBlUOwssBCGillaZnWxCOo00sDjl0PsdFkf0
yV3FwfKG7xmW920adh4/VOmcrxd/qP/ieLWUrcICm/xjDyTTfH5vNT84BZznRNIs
njaNMWkaR0zxZeqB2WfMQiZqjZPsdUO7nXFONIItYu305cTfDfhpQIel1ovdVfav
lDyO1soYWG92moLfHB41QUKkaAuP2HNfuEFzusAbOB86eiEGD+cZrTLk9Wffr0Ir
HukDw41E46MjXgr7aUvLBk/3fpOpY6ehCHRvyBXS/PplaG8AtF216jOrpX/L1V4x
lyPs0ASA+1X2mGUPFAkm5RrHk1h0O9V6y2Sc3R5bIbjceLg8G1A1fmc3tllPHmWC
Bt7tCDRH1lfROKFK7wljAIC71YL+OqdVmTyBuZ2dCNnuroCnkHmSR2MPfV23hUD+
DHngu+GQbty/DLNacjAX6rt7hBmTHlFypijAaA4j6H9yW3FIJhRf1PfUX7rT5buq
6KzFhLZvj4C1bk7qQtd/7DoDtjQQd89bhhdPdOGZwbESLRl0uf8HBWCaAIcfQaah
OHXO05V7rFbvBIiBltZqpGk+sQafDXmAIo5u7Phlh/rOUa2UElpIMvJI5YxCQeJF
GWAPNx3lzQJ9GYu9Jsk83anFWHtSzfuWOecavupjMz7OmE700KChRK89F6Th7h6z
rXLwEQ9GCT+oPYElPp+QNNSetdXvm1cxlDC/L9yjDhlF5+xaZV6MOk+QnL1mTxCQ
ZViuLF1HIL5LbWH/vGAOethiIWo1bdjmX9GV12LF8I+k+lm1sBeJ6E+WuNKC2VQr
JXHmIMZwjkTKpnc8adeWyH5Nz3B5WdsrYeOjT86HYD62VuOWxToJvu3y0ZcWUj6G
4t7+TW5DsltNk6MMwWWmvHhUCl9QJ3r6hne7UR4hzI8uHmjJVhwc6afIm8ae78UX
32GLNMc/EjsDheAnX3ciMlGvLPgaoHGbfODyg/mVF3CBAthB0xFcElV1Wy60FNQp
CbrLklop5jlmt5JPVhu3ItNBSZo9WKUHJkd6kLr6LjuFuIYNr1zemstIdawT2rkk
lEhZJ3SNubdl2/Et3WOR2IWQ+Tycm33BAUqieqJkcxMk6Z+Lc9C/nIi1YJVS5xFO
kc6Fyn/bcmklY/MAUcQ44WLAn+cO67MSWD0UqQWlicuzErYDFp4OfePHnQrUOH4H
yDNEcjtpRVd2e5X1d4HXEnS+hxgRc77iYTdQjjs/bDysL5uRHbOQUpQYnAIAsxbx
zk8PRfBMTr3hX3FfE4PQvDuRmvxpg9JvOpsk7x0tUyRk7+In7nr00HYsnLQzvkdH
HOglKf2EUGrfO0J3H9mmJJbYlrzs7FJODKRQwmfYwTSfJU2YnpNH6S11rGajDooN
Y0wdPzKW2hk1SGcWKykYKcvUA09q4gPuqtOnihrN/ClJW983KRIbYM5Xl/94b34E
fOkvlRIt3kRF4xqO7VthnQhGbHPB3aRnmYryJWdXGrkJOPrDX5dN+PSk7JQDnkE1
wj2efBWR51ixveWSq8ETu7h8Tf5GVnOIdMTlA5byY/ZZgvI3FYcQ8aHR8iWxRPmG
jJ9t2cEfAn0W1kJfR+P6TrM6IfhHrHdkv/mOyrCWNi+9U7JRi4HhYTRkMfTb0fYZ
OXfSoME88RKdsAZjDIJKLK+V20jB73QFGgpOQi6kBY35GcAO4lwntcxiJY3yjBL7
tY/o62urd2Iwa/hNMYciK9sZ1nb9bv3aquzE1iStAVDMZwIYVsFCiyqnlHU+Dak1
n/gqVzHxL0pOPSdNnqnpT4N9kKP0aC13sIBBYM7jMaNMlHe/EN22n9cDuoHv2PxM
rdMxDxepwtq1Qx6jY4GOIErggv1kEECys4/tZumMdrEo0A9pyBiUry8EpOFKxN2m
+RVJxTQvmOoWC0lTQecnxCn7aCwAzSgfN30jvflo3cU4+acQMrldX/++m7EW7iTk
2u9XEXqbs5cjJRjDsjx7NMz297zAWiHnplN04TA8tZnGvnR6Pod2ZPZ0U3FSEaRn
8w+LvWbA6zheoXU6UT5nhQnSBJCEFAA4gnh+kX/MrQWiAobqZgATXUcL01LGksqD
tgDCMi9XD6UOpEI+k1hhoKTQuVnOLoSwt+fuZbqX9b9aGwMlESF+8eqasg3QrM9v
1m0ZzuKj30ZsnExv1m57x0NxtUvL3ENjub7Wl/Di+uCfGKl1x0srWjMf/+UGUNxd
mKV6zU7h67Sm6LindaGtzoGWR49Eyk7X8AG0kuG+GdLqQdKpNTbk2OXTmE0B6URo
KwuVZUEtxRYT52R6WjS9AK5Yb1B8a6E4OhjRK6wTEJgkGOrc6XtYeAojw6Fh46dj
CD44c8VLRU3sECWwLutMS1np0X2SCYlVqkyTP9Ihm1fAsttM6unLzNKXjlxzXcF+
jc7Y5wyIFwwKKa4ZDH7e+bvopFrdJ+fdx2Wv4ljiq0NMCLGdgzM4kj1JEvrcwV7Z
wax3YOmJVmHcqYSfRi4HuVdXPGKBX2HexJ2viItGoxzgRKjLgdVF1ls4yc8vceIp
czyEPeJgFsJnC/6I4W2tql7psAwemnk7wIbVt/g6D+V5bROcQeS0hBfOBOoUO66t
DZI9iIIar8FX23KxHwIXzeJPsrIAMooWxlfkeLY/JOMgAxi/2guELbbe1GkFlDkZ
Cp8H0dAsxsxX3gGNs3Wy2vTsjUBfdJwWk55d60A64Z05u115be4oTm1bfQK+BKoD
/YoSgA3RhEsQC5jcy0IaDomPtSK+05K20vJB5gF73VSmQmgUqIuB75jc7aHddaCZ
ewsJwAvcrKmOeNPvci9VF/L9vvYJRHqY2fzgXv8VbQ8AI4BB7kZilBklag4RbQAK
Zm3sOPENOIs4KrOBy87BhSAQ/OKMkSoc8sOBQ4oWxoEPhSd4hv81aY+Qvpb6jsWK
SmZKY/22934sJQmsyOZr4shBgCQMI8Ma1ggktbPJd3mQh1QswivRgH64d9+mE1UJ
zgrAP2of6ek15toqRsuhB5HhrPom2FwIpry7gzUmB0U0RTLlBKJvxgc+m50fGZ6C
6DkzrhmDvu9kURkFRTsGkPj4h43XhilvJlo0sqqvP1wY3a+rWhaPhtINX2bcrJsH
pP0/8x5tf31ZN6UcznXj3ezw7pflHmfJwQffEJDUJ0mfC1Y++Iv/uwt1XZZ08YZy
MTObn8GvFCsatt0EvcfXH7PjaQ3zX7k1QTaOLdIWFxohdbBwmYQ5psX+HyaPgE5X
lSXlZHcV/EAV4AUgsohR3r/vtB8vPBiYfSS6XHyCJXvGFftenTWReuHfuBmvvCmG
9VD29lS97Lwn3m+ygdwWsBo4XMc/0oPBY6dYkDx/S1iyY4iWYZtnhmET10IzClWC
tbhgGVLmS1a1/rpMOkZ1lKxurRHdgTV2dekk8rMK1szJBPz3+xg2dvGJCt0buBCv
oZyRKiLjWyxdlAcFpbuRabmb7X0PUcAo4pyNoXqEXzrgC8R7TwTqc7nZgo05mCec
iuZsF8K9megDfcwkot6vWT4WXTIs8cbVxsK/GLaM8SChF+k+Yax23qkgrRYaYNZk
6C5CzuzUs5sopRtoqVgZ49lykfl7hcNT1aBgpM7NsUq5Xa0e+BZriTvD4XZCv0dJ
ULEN0h7pkXt1H4thOsD4mFlLgWfx0IkZsTInIHxiG9Py0kDRGvz7DdTSeB/+vCwr
NzWuz4FsN6QVR6NPNoZHI5SPMVOW659Syt4kEvSWFcY62CWHKGLlaAIaYkauBLzy
mqoBHsj9nI43gu8BWCT3oyEuFw+vj2H4IEQbt/BAGVGb/sfuQ8K/2CHIj9OrpvpC
dKZVjrcTZf3WNOmWm4XS2w/CdHrNT1fLf5Oq2HbWyc/nlfiO5BwwBFznGpJF7Abr
q8XGP1v3jibNIMiXUA6QuXrtKoxdBVoH1+8KdS1dLxoV8fxHDPJa15B5cMpNiL6D
7SlluKkjyt8a5CcG23ctejQJNKmEgvfj0GeJcw0LpW0gUISJ12FgzNv1twkqjxfX
Zdz/JTI06AODebaj1K1ygNNryihJdp0/oYkxe2gvbgYZtlaT5WVWHQMeESQ9ag5f
4FXYkuh/QKgQn9InubyAQ2cddiENYWmuaCwZyw+dVoK6jvlJIdAwZd2psJ4wqFlq
y9PdSNmzEpT5fBV8t0KjOI5uuNDLtV5rEjBM+59GcHJF90xi8OUHaIn5n+HUrFrR
zM9y9E6box2NcdxEowv2tCLbXANITMKgxmpjUwJTFHoFhTN9rTHlPg+XrUryKRJq
HJqQBJ1l5WNiVUwd1LSuvhMYWt+AW9OortsMQFQlogexCqDSpTb5QbcCKepWhk1O
ruzrC1voTWSV+XP0wGdi1RB/GJ1G5w9HTa7QDIZO9lVVx3e3EARmypCZU5M4nwuG
BBhPZ2QaOq/io5g7Ve8xyHRasEWIBpTnx4LSOCko1DEy/ezmGgMn8ci1tKfhdQyR
ARkzGkiXommg6d1GXN2RZqogKTxBweADbX2PIbP2z9a0qxwNJ4tffqnCgms5ZN3a
1DYNSOQBYyDCmUlAgdi2lxMzc1LDcPAx6I888C6BvoWcAkYuhFmSe7oMSSDAt2h+
dU0Nra7MPAjao/DzWsIVbYdgqEomHiHx7/42NcKIuCndk7gfgVbHs6YMUa1T8vtf
IqgK3SrqXTJpI5ygfmiPnJWc/D5f7nz8WeV4OkjnGnMhPBsbkHe/pmzojiOdjdpT
RA2Ouo/UC5Lq8QgOalOjvVjo9Eyc078ArOL7SEokOBB20PgN2VfaGykTY0mAEMli
ap0tNGxsbELef1rJw3LciDt0326g2G/v0FPw18v5eNedlyoZL4mXbF1nlJvqQA6Q
mQvdWvDsxHUnl5mpY3SpgOGZqWj7HxevH31rp58rdFpGwnTRgCOLt2AJy3zBJ7yS
B0iI/giXdfvoWMSbs9nGshzKoECHBCYBdVw41F2aH3oTaXTKNY9whAFNSe9fiFxr
JiZlQKJI8ab/Qr0sb3pQtXBU8v/nPxsVpkRkylP1Mim7xTi70+4JgbCgsOb2hd0F
Eu7KenHsM/+hozFhTVhvaCs7mCvdsSfBIDIjsYjInIOIrJHAxk2aTUlgkqIP0yYK
2CTaqFmYK0jaJxfN/q612SFBaX/Dvsi4xVQP9wGiBQ3WYtf7wVgg9A2uvJ3nn2VC
J4X+CSg6bAb+Whkwii3B82b+VZ0hjuS655xrUbC0tF7na1e97EuOQWuLyzf4tPyN
5pcwXZb6xO8Hw40cQ92oiOX8/ki+cxTxec+LD64Pza2FAm53fmv3T7fswKMnJM3h
Lkhz6Da6sEDlGWg3nzaNkPvkT8nlXIDpPKqsz9F3tCWekV5C3E98/24HIr0LIubR
PyBNdJijLmaxLv3ypzDSEWpmiTcgN/3K4xn3pOhEv9LNbRUT1uowMNYSyt06aNU3
7a4Uon057yoCa6Wl5LMkRQUNMZwN+BdQr8ES1czVIuE62H4JMucwHVSY3w/rsQZh
xYNXfHd+YAjLn1RgRy81dJubBRnSfSNbEob/tZwkkbpde8S7s1rAK7tmKHO2wRLz
FzxXp4zgGiIGEbwwKHGhfBbfyg6XBdYlVQuukbvfNIktYUPBNiehEy+M77PoPlO+
QVPxIlLxcVLQOm2EtwSRwrKLxAB65mY1F1q+1YTXrs1P+tvESacrQ7FtJRX8c//Z
3SwZAK3qmQzDVytNdGeH6AkgX6ZCaRMXXLFwNZNrHTR/hmDwfXr+/nM5EPlJdo1f
nLMCSn4mrTWbhCKZAPj3eKx1TLBG4hl383G5uDfwjfp89XGyrXm+gtVRi1DayWZz
wfFKOXdbkCK2Ta5dIpjjnw54OXPQTWM3JqPiSqIPeml9vpAUdiEEzIvCO85P7FYq
JvS8RKfvIKTW1FJP8lcysUjiVnGyD/FgV6i9FOzhuhZUmg+sB9bQZ6KI4ubQzu/r
e4rS0NQrxwK+cJn4hR4Rvbkkk/+Psa5KPccZKEhJCw+nzdhHgPHUki/6HSDyDJN4
yAcyM/9qcH3y42hc9hyy4jN7BPH0fBhWdxFDqdHq8tqPuEvbCX6az7qLmx6xkZXM
wm9VAjagKsOvgy1/OOo8sUaV4x+BM+WlYcviq5HFg05zi/nnOwKtzhLmGEZtJ2cx
2TOYvIEzxsBGBN+WVC9i0zqUzZ2ytDBbooqyJqyz+oV9MviEt/h5EVmVqDHqnEsP
sWPfFMJUtDUVozP6aUkZ2v2sjGOOMnNpdN6HdXMIboes7HTqNueAZ/58kr13DbkV
Kw6b60O5SqgIQ+Qz1/eg8wRuk1JkTPub9bRW7k281Fd3sg97iL3HsLzGuiVJLrWH
+zrSz+6Y0ldD7ZkkeEJDXbdrc6EQkvxneUBeOsI8pm7QYm+TFZjZ+HQtGXZlzL6h
zSSKmTqccdIQGAiBa1yd5CRB7QavJfcMvAwr5QdY/Kh/8cQejJyGL/+AVvGMMOa0
Se+LDtvygYqpwuw6VIUcZGtS8y4kiUxo5G7DeAW6ABr/+Z48UnqAywXLi9jpzc4u
gKB76wnt+sjOta1I38nRj+FZh0IQ6ZEleYzWPLbCTOVmVjXRkWRrOT5gRlqP1MyJ
5gvNFoQ6v3cmZTigWH+0IRMwrQzt1uAghomMGMQh0SAwlLxeSJK5UUgUoVxgtQ07
j6PLQL6qDGyioHywfClEvCdEVKqpFoQi89uJSkdMIvazFJHFvjDUJ3jg0RNuzcax
CyXYgv5r3sSOPBjRKJFYHT7Aqsvsz0reY7kPaqWSdrPtOlS7q0G1jOWZN1J9ANfx
qiemUATcSltzoQeQOXRwEkr9YjSsbf55+pa8Z+LDtqUfg/buN9uCX9BGG7cI1+nD
hh9yDkYz1Zs995xTZIdST7hwaS505m3fU8K3TDoIVxLfEjdyRZRp11N5y3PoQIHd
6Bn2p5oO4W4VaCFuSGMiwOSLaAGoBgNEg/BYNayRDnSPPYGod0RDv+Bh7vGfF1hd
dEByM/4YPweh6oEWEbX+BVtYbRY1cHgyhBySc4Atfw7bSBLsfWyKGoXuS0ionp5F
nNhGs+QK+cseZVCv6r6x5XXy6jhe0D3kdntnIwq9kXvPWdlbbRW3aar/C/iJ9pUr
HH5bQ999U4eOagZFD98xFtuovKQ7An7KloCM7VQbhDGBwKDUgCdEb0K9xM8L0lTw
+rmjPB9FzR0BYn4lAMEW9Folv+oX+T5luEnq8h9FGOiBu9L9RHoS+coR4CTNMqmA
COXjVgbi63ql45jND1VaL+m2Nb90K69K6LBoO2o9BPQY205L7rpi02ouz6aH0kBO
/GsrOd1laWdVH+R/8VxgRs5GE1emR17zEV1Mp0QQQH5wjBuckMfAqco5fwhGne3w
h9reOTU5U0h1Y98/Zfssfl1fKTwxzJivu4Oz5/tyHzvvtOJe8aH5kGpZeRU853R8
J0KfP2Kd1/wv0QLtPwQ+8ypTIT+wd+B6nUORpPjyk7zbipUdyzOb07Vn782le48/
nBhnjdxbSThkJs0ngK45tJuMiJLL37bNnYtQgsGh5WbPJ93EW1gWSUdZUVyMvpj1
Wz9V3jWyar85tj8QuZYQoCe32OyCnZbCDbZxK5HLwqzwvFxDnHKdxKGakuytfXdE
eyhD94sjl+wEQ52RIZ3YN3S57ZrfDQaGtHoMZtgVVG7sJP5o6VLa6kkNc+BPe2T7
vr9RHrPP3kk4p44eri3BK17C55eYlhYqs+/yGbwvdUqnrdhTgUhxSh1+FD88yqbq
k0lZbbANLOVZUbyAhNmemPOFgI22WYSfkwqJBCPephg9H76ZJFLcs9w8dTfGxow/
ae83bYFJuTqBPizkpHXu0cST0brWG/667k7UPdiJ8+1nllfMubBeZuakrScB31VL
NG8lVyQ0oRwjGt/3Sez3eD1k/SezDU9Ugd2Gd8i3bYIMSsTNPj9Tym/+yWKV2Iog
hMMNb08IgFPuX2XevYZKre2MMrOx4aoNB46fhEOoTSuHBpYAETrKc0sXNfltjDI1
KpwAo5Ad5FXV2QgtVOUrKHV7OUP/YDRJ5Z7TLluLeWuvnOAt4igA4uq0gABQq+8K
Sklc0/1ziuMDax8AZAa/vPvHpTQKJOFJbe4hZdi2xUcLkNnLnMBP21lapu6FNnQW
MeC4xhCu2Lj01LdfW1btEW+EunO2wXFJ9A7nygiiDSvfhXe+Fc3WQIJDFU+IfCNE
hQ5rpZnvq9p7Pm4qFnZK9gzE1kb9bTEEE1vZtV85FLkKwHB3pDYJ0RcFJ26LymCP
mtNTlkee9JB9lw82+xOL4AmDMDn2UGcRmmA1zNsi7RxqxllEIlwFKhCWdY/WT0aa
2PghtHDXWgmiD/ShvqTHWaaWRlt0wHPcHCv1nFSYBjKj1XQPMhZ25OpSY63Gu471
q4CgHtXbjbebbDwI9+qbHVLcqw+IGNgVTTE+CviQxEi5HhyoZm2kXbGcdpVzz5Wv
bG0wxW54mFy3Ieo8iQSl2UQvp/lKG/CMUVFGPK1cFhn7VTeW+nJjaC2Pp7e+coSh
yHMZZZs5DcknpJJSwBOiJEAY6E0/N4EKimmXLFO4xBKI3LiGfOReXDC2LHjLDUcD
j2zLdY7tdGR/RlrrG/4rRo3AvbPM/f19i+oXng76Evl7K+4npWww1vKAc27UkDbz
QoICr2YeeVo93en7KqFUnuKQs7R8xHuylNjT//bGS03vGxNcV9vmzidJHek1agbC
r9MJfTEeZfyQaJDWc9D7rE5XKYegIuoDanWrF1a+GVofOaM9CzQlbNbTJuGg/HyM
31gxZt9sDXcP3y1uomZse7eiQo+sQVemgWv9RzWFhyn1xgnSzaGiz5HnIU8N497z
jDHSFA23PmMjsxrfnkxyEakg3M5eJfsCDIwHEIpWiZvPwQKt2vrihRhr5+VcVxYP
tygjBZN0uUROw5c0MHJmTZLke33kpJ/XzBZRO9Z4zcSdNprEIy64Jo7dk9QAsp+m
AmfRqbRjBxbK6awMk6BM+QC5AuzV1j+t9MR04XwWcm5lMV5q8ykW9m5CGD4C1nCt
tx3YtDBeXQjyUObgK7PEI33CMgqgjL3lkJ3iAtz5KC10/k1FGwFN7EPEzacJpuGd
Q4LYdyldqrI9Ndhf/WFsLKZ+HClfp9X3ACPB+r7K8rGVM+JaWDJxXOm3hTgMJuHb
b1gp4a/itVtzzVsIQKjs3scpqJx7gmdQQQGPmx1agX7FIrL4Da/wU5PTfVSOkUmJ
SjnAqDLseBfHmXuXfG/MsG5uRPuQ9iB4YR1jOrMCxnWlWJI9FbVHnA6f6hYq79Gk
VBGbhHefsua8mnRef/W+p9BdZsvuJPf59TITwZO3aSOU7TIZQr6RYYGb3lwULcAh
zJ2CZIDDrzEAiG3PXco14thJg1+m1c0roTBz9P4Mh2ZzU+BBQ2o2x5XuFn1jMaTZ
fjoss0x58ite8hRKm1yncA+9pLatTTcnIP8avKcu3clRHkRiRVcml8Xrw+RHl0IJ
iDayepwIcZowNf5CvU+9PEUzSjsPLX9dEW9Y1NZmiUvIFndT73iQjkSfMtmzFXUp
q8gXwqdMQbeetCiTs5K/A5B6XKOaaT/rXz5CiYFJBj3fSxmXQkx+OA8xWbJql/Bv
g++oocGl98724MzE+2sahfe34ylqCgmqOmflJkXN3BpMigmRKpQ+fww/XHdvqd/J
Y920KiDnP9FeR9b3F1cdrPzjDBaPDfRVSZSz9SVWh3jpkKqoIiTGb7z3enuZnzZz
Gm35O5ColEtYxfav5AKinAtQzo+RPMK3AE9lb7uwpnRQPk1u/QZs5qWLeqVOa4Rg
Q+Kj3gQV5T+s93wcfZzhSLDXSTXqfhyDokOssahufZS90N+FyUOKGuL41lX17W9Z
o/52RD1fc7ajqIOWubYvzs18Ni8wAJ/XdbscXDN7zJWHvqjeB0mJV/clyEUJqook
4MNf98NgKPfCOrZnqNGeUS6ZBiUWyDlwIe2QWBmZcwsEjyF5fYRARp1harpf01UT
OBELkBVC/Xj32KGS+Qp/WiMLQ2RdLQUYFcOcnkZbrwZwRbgT3Ubr5E/jrnrB4XJ0
pzBaaMYlQL3aVAizRGeEowjVhUHrSOyqlPmxJBOpJxvoITW8LCxdd8HJTa+Q2N+v
8hzH8WhT5xrszHDQMXg+IoOKcd2DN2UQSs4af5Xi6A+8M0LIc+faKokFwn3LGSfi
7YdBYWJc7u96rPRDm42qWDZDfT9/Upl35JHCnV15rCRo/Xy/WL+CXkgrW0gEep/9
67f4ZyCabMPOEZn8X7fqNbq/eOODi0RBBbxFPjcyBS4cuJmZaTu1lOYw/VoPj+DV
ArgNnc2u8jjkTPPU/g1e77xvFFJRM/1ahJ3mdu/iIebIap6BrRN74OqruWZvfOgq
6rHeG6yq2+8J5ui/XA9mqx82LBtX7jzW18htei1DcnF7lEcAUoe2IVD1kutUQ8cr
JbZh8TqV3s9bI2q+IdDR2WfthYYDJqFFIbq6nRqPNJASE4fVZ3Eaj9JfOs9nYi5A
7pPjBy3N14lDNFFEOqAvcUXQrzkNSZtZIu43IFCyjYfSjnNtT2EAwgqVdwDZUegR
TKC3hdHvX5rteplCcog63eReTsR+LXSvVCAVV3kdgvGmfll1FSWP46voLKG4mCOp
HwjIkNSGnYF0Ejc7L51QzspHeinFVTFM4bDSvY0fcZBVO56ETRAP/5ZM7rDtOR6U
SOTbzIeTxgUAOXSjs4OtlDYTXNja/LMYJzXYKzjzAm0XyDtJv4jUUKFmK/QB48+Y
ywv8EvBk7uJZDwTwqas++hedzoBuJEKaXA182WC4oywXlVP/o23VLiQx3FTQ8Vka
ZTNnfa1U2CGJGG42RwdQc4Uirdl2RWBgFyXCfskBZDHs0MFDPWGuS9MdSrsW47pS
vLaYRHuqx2PggSc9b3nn9wlMTNWXq059E1f5FvH6oaWdLQU2xRpYlXWXLSMv5AyV
vUUuywm882Al0KhQGONfjxdasMYl770vlzMq4SpN+5M1rl5SX2+oA41cTS0IH6hs
WTXo0YSCcu4GhkAmIK94rgw5QE7A6aED9OtgWKKnC7LqFc9MQ+zpaqrk+Yb8B7KH
lsyLx+m5dswYDPtp4fnexPBXkwkz4u03Y27TJF5bhRfvuApT2g2sLderawKTEwV4
UfMPr280X8wA4n15vWPA1khAX1ygreqGNtLZp7Ee5cjv6FjM4r5/nIY8qsk16VbY
18Q3ROMrjAlCjFVXpQggaae8+5WUHEqPfhd3AgE9zqjLd7ytIpHLr9Y74DXCrYAx
I3pjDRlF7bPy+JkXOZRi5k4QC2WQSEEkf9mXFrUN1deEKYyuddL77vQ/NxmD9FrA
U+R3yN0WQpsXgWoHf6IdS50K5vcrp40fzlsFnPDwfM+PDVv6HQ9dVFBugy9oeFF/
4WvUcDa9302Ro7SkaS0d+iXAYazOh2RdSUuwKBYzoooNAf4hD84lwukEu1G87Nm5
yUIH0jB3UgdtcEw1K2oAZZsk7PBp5oGQdzCYe3WZ4yYYt0Y+Wyc0kg4u53p3SGPK
mw/3ASPmpmmj1mkpImq/x2FWa98Iw97ml40sdOyrl3YnEPhzKS3QpiWMNBoASP1q
MFQKWCdSn6rcJBjEjm1TWMzUm5OMQRgkPqi17tXzZ+kE3Ydq+oOhaRax/pLo1OmD
vjr8xfHfMPouBc0b3oeeYJH2ulsmpdIk3F5ViIcm/e8bSLi8YtnS4/XZe8M9xOBf
XDpxC8/KPynfnH5vdFApe8NvE1WlPNofAsqsyLxpQB8Y1wuSSXsZxYKpkdG0av49
eTnJ4aLQd3LV6PeSncKOjnGA9cHnzji0xkDo1Kko6vVyQWZGTLSpBS9mMHBLmMbK
OftAF35uD226HSeKzCKqyzNROrpc6uZg7E9aw0ER38eBv9O4V5vCCP+QQpEUUphL
7plL866bdBGMoJT2m3nw++SSnPyefovON6m/LrwOnKLpmfjSJlGh3dpyVV5yx5rq
NJccW8XiiTKbLDIaS4RTQQ1znRffjHJ91wkBt0D5p7VIBKQYGAmbe8HLLZnkyNNm
/6i/1I1pxeiJ2P8c7PvSm9JIzdEp14Q4PyYskjh8PQgnTvtibuiFbK7RAkKleop7
8zL6RiAqufvN66qiv3df4umefLiWbc/oT7iFVcWEwuzhfC8RovtZgbyr7QHkiqOj
BjTwNPS8gw1PTDzeW7Bm4qIZMtxa1DoKFXIaBwudfASXO7VR1m/E+zxi1g8oZIYs
GaXpnxXMBLXFu73VA5EQvQC0K3C2h82b7JfRsuw1hX6QBNtOy5fRPEHPC28nQHP1
10JtCcMGqmX0f05bM+z+YTpkSwRqBlxEgWGGku11ukXPnLCAMeB3fah9g2OhpwRF
gRaS2DfBn6/aPPbpS6XkWZR3XEeLx0oK7uEEivvnoKziujzUT7JykUyjSzS0mq1U
U79pJBjzTvUh50wcN+CzVxG/ixS29pF1X3Op2rxDHR38db9pWrBazIT3iFxkaKHy
4b7jLsCZD/Cdc6zp6f36aCBt/6vU+fsTCqJGWF0aNwnsAUdIe/aI56gGKvWfLfKw
jdEGjxmHoMRjs87QD9HXRB5lmgaVI/QLDXT8L5sWC/sVgKDHFK5xdMhL4Zsdynsc
n4TaYLMlS8ZqLOCQVm+2k+jNN1Pylt324xpNHmQdzchb0ZPt64ytOzFJao7qAOiH
WuXGssM5vqm2+D7gBaSQPjAFOHKBacxHlU6ooFIcPrZ8yaq87QiNY/BZCW71kjfS
3Jm9+qe1M+0OZpDirmV143FAV6gxP26LrNzpcJqBlCn0W7lkLPSudzNvVfr33jz+
qMb6a9pJQh9vpTISSVSVDwdizWAmBtXC5EYdznNCua0qZYm+lDzhnyUDqh4DdxvG
wx25CwYanOF5OXvbQH0WI2ZdWbO/bZvwtXeLUd1kBuegzcufiH7gkAZkyiLsbdVN
4vFn+yQWIF8pnjiL1rxL0avezhawNw+MrfDIK2q4Uk+Whhmm8jTyW25+4Pge5ifq
+cVe/c3uT9RU1XfDORuJJHBURpky/wu9QopNNFf6JdnQEKKuOuJBfq2vh5duY+f4
R8E7fiozouPMWG/66SSXAtR+w9jrppGNjQ41ByWDqh4nnCtOiJTIvzvjlZKB01BI
dXrM6KlmXHQ23WgIN+rF6a/tKputTXntgJb0XbcS97nVAr0FhzpkQFQ0rrPb4Qgy
gW+/HI+SF4x6bsHEXHKnXkBE4GN+N5F5hUABN+uTqcDkpZNqaeqymj5F5bMmh6vJ
KgY0q0mZ6WRpuZEpPiMWVSam+cOMcb+p9ATWKMyRSdhCY0inkarjNq+f24s68yuu
UwetvAzQoHfFHX+SUjbjNWU2kGzCOtNUAx2W5TUDEjTmqovVLtgylX+opkxHM5OE
aiYX3nusBu5QaRHxS1cf87GfPCPOaFHspkjXMHDnOVWOdXjf+Yuo+EZvsITZbcVE
eoqGMYf+O3Ac8mZ3Bwh1BlqPmS48kFPZHhT7PtDUYHLW0N7ChNg9XMk4oefJAbwl
oe1mDoMbEU644JieG25cHwdT2LP0kcyyTzs6a9K/BUPTMqoPeG+kaHd9n/BC3V0e
o/5qVe2pdmNstDdL8zrrRmnwqrgdgylQW0scO3laC4nXkjjqQwUjvf+mP4BuXt16
qUQElKD2QKK5JfK71cKD1i4hC1XdzWSA4VZwzNoJG+9jaUachDRSSBg8Nl1JHX3s
22sR4EQJPxpPUqzjAeXle1zD6JwvsZFyayVY6sDgkou7tEq12CWqoAWNkQtOA8Dt
2Go0MHSv86tkwdYRL6RutXm2z+HheuIt7DRm3FRstAfhiIbjxze2eps/0iPTezG9
WH2kPiHsnXHranMcbyR1DsmKCk9bRhcEABD8SFCXUNJ7dAsi4v7zaksCQwdBFVig
gB4nIbay98USixJfdqcOK8lERGq5pq8sbFftlRLrWSI4qYy4zsNwfSdMO+3aVJUG
F/Msa4/awAGqIW3i1SgR+2TrZNRM5kx5NefbFCickHhCl7LIF3fze1WfMnB72aYU
sY5+4lYesJqo3icSLi+XgTJQWjAcSnHXO82uDfSa2y16AIRdJksU25gdtxt01Viw
aDQ0tuE0Vqx5A3ZxvtIRgJPq1NLEH3aYoZvqiLPy2hK+pXon8RFFAscATzsgR4Ax
aMwStUERznPZW7rNE1Pj8vkBZjoYCoan+N3CD0CVodKvLL2KpEV5OzCp5n716N20
fBpeVICqJz2VsFQXPLJRFxMpoGUrP31R5fBDorN41D69U5OcCHwhJxzbAl3/zule
5XoX984+GBHYqjbfqr+JZGrfN7IwjQSVvSdqCjTcd9cNzhbTS+XNIAGxno9xgF5Z
C6ZYfCWQfR1h2IBwpgZmMTo/82dFuZ9FHKdpYMSr8DTehEUl0OgFc0g9ZaDeXWIn
kCcXFJwukJSd/9ACnXS7Nqo3Qpyn/1L3lwYO8TPkKniEfcIopUNHZW1fk7n8LiJw
1yiSzpFCA/Po3Eef2/qEtv/u3RVJpWKpUOJP/Nczr4TrsPsSxogwxQZbPoz9cx8o
9G45RyFeYqhPgw6OGc0v+ckIeU6RMfM2+WY8uftzTKizkDoBi4E8Pb5yGf5DKYMZ
8v6IKmR7/mXcYMmvEqs5frBNe1B9I1lOvLEw7Dt7f5m1u+gcc4U1HhZ+joKp5fBh
8WbJS0beBCktEBq+F2orx5caeShlhN5r6++hQcpduIn0ljfpQKW/uZ2hQOrIisNh
yXT26rw/d7kXMoFTvHb3XT8JZNAdOLn+eqevfhfoHRcnl8WlY9ZJPs8q7YEJ+wjP
/q3FTGH2z086LlF01CvdoHtbGbrQVVRRxfADABlnMEk2A6IaPEKYAn2ZM7KY4caw
EKwxGATA8giQQK0Q+/YyT3xJE31OJwC022j8k/fod+0XVYzPNVgK6AFfSA5do3L3
AokKQVfYAh/h5b95MT9sNxNAL+nj5410wArlIJO5eAaKuRJwQ3QvtsTI3j9/rdKU
CeYMFBZWpdklkIAcpI2juiWqcME20ASD4d2bOgXhC9ctqAXY2nS3kX+sA5Qjp3oS
Vdbr5+6ExAPhtBlh1z3USGqHHjSn2ZNgXSz143uX9dFhW/OYLDa/QsjHAHcBxMV5
ecxnAyQ9W6dvzOcWD6INrDmf4oqcirIa99ye1uA+zL5L5G0SttCUjTJUhhrVObIt
uNCAmXxkrVoartncshVuXC29U4fCA6sh59g4MahtQ+TmDyIs43jCgnYDdbJkdeBp
MduZAxixHQ8diKKmwDN8eoAzESziswq+dDeolAGHkvDC1232BdbUJKYGNi7vbS26
Ktdt79QqaCBXxWIK7rf69grvxbxCAfBExyEhDj0TW/Ydp+m6tZfnfF9wJ+NptayN
qvYnWeuaTimkbqWV3R2mS9r1VgIbfkgZkCsiCm/kUcr4BLd/rcGDEu1N5dBSMtRm
jQ7r09/Y0nz2i4erUrJtcfCCeaqoSQxfRiw+vtnT695+T3Lj7Unsb1MDxiZ2PhfF
MwzpsgLXitoETZ4Ff13Z+XDsibF9/D0BYDfYxI1f138GBtbHlAh0yP3zsRsfpRMn
s5s7kIYg+27EM4AyuN4JzW0xZEL2M1rmMAK0BDDp9tJXPRYH3HM+S546vorDawMK
T0TGfyrrGMQig+CsCHYWJabzYGQxNpFsRaFeLBt/GVwxNvDwTBNoXiewOSxeUXm3
WmO8vAug0OIpH5oBi48GeDxcWx0pkcl1lByvq3GTNu8F8FNkbeTZMKLWgBdoTBZ3
CtbK/+vCwE6qnd4eZmQrdSAGwG5cf8yPniMssYd3Vh0AGwXGCpF5rUkbyQmGROlW
S6cpz/tviueDh62YhmBt9WDvtncgG1+BY74rEnaI9zexbncfbdQJGWRoLYdvnveP
xRKj9GHN2AX+qiuboStMl5DD0MBs21BLByh704xmUxSiuP7R82RWhJwKMM2Cy464
cZTzecMppvIpHa9iTQS//WY4PkfmERgE2YMq3dAxaIjKCtEqKq2W1vkuUJ43J9nN
yFqMzTr7TDO+z7mkMAelVgzIWPe2HphnJHuMmEOzEGdzGRlVGBoVKeUulvqNiRYh
jo/hm/K+B/2M+ueE3ve20ocBMy/+MEmrn2ZvgoTLtVB4c6LibKzLdOpNia1ETm2o
C4jtF55umdV98w8t0Wa+CejGee2t5uLrAyxzJeufkNgJxEdgXze0UmiogWeEKYy4
kI8h712EAYx+PuSpKPdyoBK8aUQkZDymOlckiWdoJl1wMdLJl8HXU//QKV96G7e4
f7eJlPeg8Y+PKBQIKJep4FCaeNlPyjjjSiTShG7mTimQb2HSCwNLbg+UubzI+7xZ
YopCGq7NxbdZFpT0IotCAOQnvV8G1Q1xkIpQozhtYpBRKXur9WYiFEaqhmzJW1CA
O79W7BTT0/4C6dT2jtsvSSUpCJMEefJGjznS5UAhCYAzTZic1JPa9ssE1k+8PwRe
0pcDMYsXsZvhPIIY6k+fYeWx0e2TCTHdzNDryb6W5zF0rpgE7gh1aCcvsIWJ6bzY
6gqkWEeKX682db3xZ7fHWBQqFMPYSpQM3F7KPbjveCUY/wPakr80HYrKQISZJs/k
/fLtA4gBb5y20AJksJIqgcHxbD0ePjrhPUyXB7YqBqOngpOqdpKm6ibQrzoRlTxb
L0KZTAOcI10BfjcnnkdAyvz7J0E88InHJND48dKRq4182h7wA98wvMZ3PKWF8A0z
FlgvLFD3vjz/NJolHWmzbf8lEwKAWNmhiNvbGZQfGrIelisyQ7UTqXJ3bgWV2oYg
hhES5GSshWqfenFcNisyPmtYWAIyCw5+igRfREbLrTWhfAHc0wfF2iEz6Q1MKMuR
c8yvDLLf09GJBYNkOG6iiEUm3njqP1NvpNLPc0g6lNP3aN+YKu5QJKROi2craxIC
he6SgzPMdFeUzWvdqV+JHd9vYfQnC+d85urM8OLAFD/O8k2LQhfLWezkhoAbXr4K
pffjjrj9Lx7IZyYlus6s9ZG+u1ssElOjCztCWUd3oEhEBdES1kfa0jUVfjBt9SNV
/OQcvpGH6HcsuAmN7YYTKWiSJl+k1OCnWmRF3eTsYNc+lwv6hmxpC8MUy/Kd0QZ8
kOESO465qyBkPESAPC5ync4aPSsi1F55m2UrIH3N/a3qdA+BzIU1YrkSDoGrS53S
CXP6bLq6WZn1e/XIsZLSl0GdHuAUE0OE90cUgXctr7eivwVeq5dk6VUU8H+XJ9wa
JBIW9oMqmWeGTPmowWEPnYELjVdg8tk85Y+nhQGTQiGJxHe/yyWYX8duLIEwV30F
uKf0oGUsaQ5bLrizsDxmmrzs2p4XG4ExOyGHA2rr9qOJCM+8utfebE1OFcTRwuzm
XWvoYZO/aJUl5hOuuc0KOBwDzf3UQNMBvkuLrctZDsOFHjknP+2gHwOH+hsmBPRg
+jE+D0neLKIRdNNAmHlNSdzh46o8USWeo+izahNG9sVPfUkksekYtYejKU2MihKr
O+zkA7VTS5CF8SK1xwISVNuu/Cd+x+47JetQgT8MJUdiAt5UXwkojURLZCrz00tA
FRjeDHZGOLa191NcSvWjxPBjfGlamF/+zRzjW0R/YbK1g7P+Fa059UU8xtjlHyRG
mgZMKeDqxum7LqhFTdHoh7Yu05e0i4Y4wQ0wglcEpZuNBhCq/ZrE6OhiF8ESxa71
V7R+liK0SMh5VetF6PVnc+JNiW9cbCSY1Mz4E7ekIQglsNq4s/MnT7Z9ae1yK4W+
tl74NYSegwGUhRtoFvj44TFhfFswCKHXUhmms+mqpHx90wdLvWmipYiopZp6dJLV
+V/YCz4y5JvYD/E6eJt90OHk8mPBXIVM8jElnNoSXKmUg2dysccWQksbJScxrJ3I
XT6/DB+Xgw7yffN8H4K7L8YE1BAaHweikzaGSK2N2YFTZw1lu/LbTEJzp5ZXdIZ3
HJvG/75RktuVICMHeZJdW1Bgb42tU/Bji2MPKvrGCnN8lEzPGqYo5E8hBtZBnmEc
u2L/SEhcL4xKnUTH6bHFod5oC2Eti82qCMZamWAREv7NadcOK8/FA6aOSzYqe2Sa
odfnQJD+7vhaY7L08l0tYXEJJXpZOmmg8SqfyYQzHlqc0/Njrjc0qIMyurOyVV9K
xyx3fNPjx0PyxsaG9HqZzrTE99v679gBSW9pVgUpXU2rAGZt3UkRZKql/TkI4jS1
khJFzHMJzg1ayu+2TZLnIv4BvjswmXkT+M9GMYGw5kLvvA01rI7jidVIfWW0jRIj
gVrIljAy8OjvF06W/WnH0McCxHomsAZZyZXe6zEvL6EXHIh0y4ahfIvAqjUmrAEG
pSh7UPEPQKbKFGPVRPyL8Cni0mibxkT1/Sd0TYqzyinCy0jYnAtaxGwd/HoPuiBm
vS0HiUufFpk6ZZRWj6Qc7KUbeKOWnNGyJnV7hUojGxJoJbIoMby23GGpgfngTRsf
ZPUTEHWigo5qI39cAJF6dbwETtf5TofOcxCXUG5k5r3Kd8kgOG8gyrU7J+KJJ/h3
7UItTT6esZ0Qwfx6hMZOZ03kwM9RBnnaE5KYz/rJcLypGVlpon/hAEq8OHSswliZ
e9eElJSJdhtEGleWmLwqmW8Tvq8EFifXlWqUIPTksorXsZbcZkWNPBKUXHXNT/Np
ECaZqnWO6w/jwJq61Q8H6L2iIgCLQxSLupTRcfmclWqYbnOfwB4fotXANB9nT48M
MPfE9lfB4ePjTAMfsItludSboIzQ/ag0uQ4X44qqHF3RCfJv+N20MxQ8jgu3/Ngl
QhXRIa/yuM8W4FaP+1lZ6WYARWy11O4FJCywZTgZ/3OyHhELw9/TjGi7ZsqkuiWL
XPSzG6h2Cz4j8BWZrsBB8SYBLBhNRVGmu8ObCBhbKPy6RZ+IlXQ2tDatHN/nLrUE
qY5pGVU9C8UKGsy0Q421KbdvCWkH6FNlBOw4Fg2artuv8yffkwE/EJv6JzMv3MpW
ApggopbAXwFl0Ym8ksUD5mXYFM8JjAdI0nQc6Ls9H1SeKQVSglzHRe4z1aEB1FLS
dWsrje/irKpEC6g4/FiR6Az3Gb+IBuAKd+Zjp2jvdYac9p+lPLpxpPZOJi0bD6V0
jwlH0z1sA2wN9vIN7MI2/uOorh7D6QXUMMfOpvtda2BUakzHp0Sau3fKh6DxtIK7
qEukXr24HIiU7BtyahvAHt4bggAa+3buBJF7bbIvS/QnzG0z+iAnIetwJvqfLkEf
/2h6130OWLwdNMCjRxoRZu++5UViOcT/GFvF1/LZGYx4M1r40KU1OX2ft7tX1mzT
eqThMxXEqId78jCJ02gx6kCBF2BWnxY44tQOOvDtZyHXPo+E69H2CAzb9DAF501l
ciY1qY8/A2kEww5dpqBK4BYfRja0H9D0ULqMwbxcajitTZ0NRzcC8L9YwotvBLGI
3/gcAaP/48TY4Hm8tdsHA9n5Thz67YrwhXOGf5yTJulK8Ggxg597RnspYvJpKMjs
bNDtB2uDobrA9nT6Y8rZtFKOsmvBwMAqx2i9YdthK2cg7vN8AsFOSANGsLlIjArC
CyokQMQ8NzheKljILieHXeJBTCWwe0aeOJhVl/zvD9SfEj+3+s1ZEg/r2ZEvbLIj
wjqnmS9VRnxN5KPMf8yPayxI7MEaDN6ck5euQOltdGIl4TUaQ5Y71h/34abaAHcp
uhrZpkeEAs8tMoc8r6zrkj821fEV21LOGBX86XRRL36KgiYjKazwIRLCby1KTGpA
fhS+tCMwuAcREOppPP4SPMllvyUYCEf4ZHbJ+kcpeqYNQRWlFNQVzg0UBXtjA2Mq
VxzILIL7il0erxNImCRQEYEbWfqWuM82mbHnesT4hlBSrQUzf3y5hdITc6MPRLvL
dQ/BmqgEdVv81karHZDs3lpyCz5abSYN255OsZe/3uW9Wv0KmNn/aOqlyH2hR9HR
uoPbKO/WJZTot9+IdluJESgGdLFwYAuZBvzCFf+dUZ9cA2NgMGqFC0pXMaiic4HQ
sWYUFC9oeZGKT3XDry5zPHkbiiEPuRPhrML+Ou6UnnRiXKBc5MXo0XumfnxiGNau
9ZGnQtoVnfrDE+mfhhf3Se/YXOYjcd/+cowiEWMsQnZvz5B/r4WiBTNuKCRquEXB
0KImf8n3L5J4Q1g+YrEVFo5+mjbcpz/5gRctowKKB7x1IsYr69qR6yeyAyVl1itR
Tu1l1F5SnWIHJr5ff/21BjBX/uL3cAj9ELs0C1D/1Q3ChxW5IJJiCoj5LtgK/IJT
YiEVz7Smn6qUxYhN9PAt2wL1Q1A7ImiPyQcQoq7Hm87ce06uMpovolavSix/nwtn
LgKsVprM+bH/xXc4jTZOs89Sv06+q9ouRfwgYcYYXuYH6uJVnsWFZJuZ49VJCpdp
l+EPcmdaELwJGqnRRsqk0S8VpmXCpQq1Vjaf8WKXcukmmYwm2GlU/6lHT6pTzoj+
0XB4IMcxnS545juFt7xtyWwwp1dOCso/x9rvwcTEvqmKJKYoMZT+LepCJWXynKnX
dRKt/YNt7g6RlqlRS4xpEQz4NtAWRuZThmW0wa92MQHeMKvuwO5AyTwGn3vBLGNl
ARQ3bN4uBdfKocZyDclvU1/TRudTn6fmqTfIq9LEBywwD9SjBb3gJBV3jNnOe5nn
c7iQFeDtme+Zq6PZBr2DumzzdZe+w0fWV2iybQxyXjnRJzkuH12tNYs0NrvBiK0U
ZaR2NfNjeHwVzVQaPwk1kn6fFc7evbWIDaYbSv00HmNTNVPNmL3YUu7ThualEO2F
ffwj5MKHNTqSs9W7rYXu7Xrx7/FemWjmkwlH5IbcoLBf/E/7KdEdEsdRmwnHD3Q/
mTBAgqoGgkZi/hzpdw1vQ8tEhWM5W0e6jwDsKbkGzblfSi9TqeZxE0tUV4v0TM3n
Vq9J0RYkYwf9tQiqzBzcFZdRkxKRS72NmApY3gXyBzC/5MzmCCApxZzq+CGC8STr
dy+UGhUYXvemaM3jl9+RkFNaK6FzDgPWVHuft8rkvs8K1qkij6bVufC+OQCAkL9J
qlMmnJ7wlwfTsnFZN8Q8Cdopavg+3uzXr9pPCp55RNND0J8WCApvreXiZJt0A3Ss
j5mFEXRL/fOl2sui6zpLW841GLy1T/yBBzOY319CDuICaa+oPngWEzn+jJjkJ1q9
WInyuDyobLeHz6OZsUlEyDYmGVsidBakdkxL24iEFmGem7cwexLJokS1XzNmtvsr
CmA5KutIjfD5GVVpgfQ7cncuXXiJ2LdLv/gI9S1BJbueRz1+hIn0wzeTcpnXTR3g
WgG35TKjHA7AcAzhK9n0CZEXMH2Q8sin51glekuuoK6u7WfRnhO8cpLjJDqXV938
qDNHwlNO7oK3Axp6IviHMFBmrKQxp/tkflWUpJCmJCoy+lZ0iHKTkoyvwdEgz1mW
tZTd23A9CdPIhBUN6Kx7I4o/oXNsHbLmBx3DABKbpuW0ySSVrWaekfJ/xzAZo2zB
PzQTOgGLzEdLcRkxEv7w6I9AXwZtNgQxeQMBekLymTUg7g250eni4Zzraddc/f7I
V6CuZ94/E+77fmMu1OXav6Is38E814i4dMFdJIOlT3Ib7H7Hq477AvjsOPrKDak9
5a1nngAq8g3Qu7mkO6JKoe5UrAWpPvCVQ1WcSp4DNDhAuHfHhZghrVCXucVNJqHy
GRvDTfNTO7vIATG7Lrrdt4os5yLfvDM+X4rEDXhasyZkok51xxCHknWZEv3jWKsm
jKc1eYDy2CMDNeEClQ619yx8ioVOEImGxLywY2PkV+eWKwZEcVoK9h1SH1IXRrwX
z4AO0dCe+LzuvyJ2U3la15pQ2WkgR1g/0M60BRv6JAHVl7ADl82vKyMGInT9Ey6h
NJHSNwuMmDPISMOVKeaX01cukwi6KIh38xGKZ4yLQpSqz6WdDFrOdvC49Gu7acZW
ml7H3mRKw1lTHOFRsP35STLEa8ciPivYEHkvDIs3erMSeCsHjVR4aGPK66xlzdLO
FnxdOFvStcN1XiTw+fJK6FZ8S4JAS2YuMI5sElqK69pp4Q0i7dnl/TkfbJzM5iDI
YhRfUSyj5zhBvFjMMUWVIBf1uUJ9vrRn9CCh5D+3eMlevt0dCkkhbR9sgvqrJwHt
ygvUuNpHU3ThGvTw1Wdh89bOShzLeTURVNaDubJS3e4CGSjC+/iDYKzyzzlsV8PS
m5BWVXH44SmdbC6jY004EX0lk3DyMl82Dom1IaWfFsxep4BIYSZy6IE481iunFdb
chDnsuFIWnQRxp2Kk4Is+12UkwMyqC+5QsZGUzfcA67SNjYbIqDVgYAuEMOYG1+T
10Qs2/pgQByam9CN3k9c6QGGz3PboNv5ez9mDWE6mO4dKxafHvUZH/sce+6ZNxph
BXKL9vYlIbd/WQBQ+Id2ZOv53ENM6frrV9exQjKXYYt0bE9E1qw6TbmykDUGBq9i
B08Iwajcd5npmByRSYrpitZRvavLC0MFF46KUPSjw+k49yT3WVRySVP79MJZj4bz
4MWprhvyegHgdOan0M0rxbZ5R0QN/n/ldItqzgfsQ3jVf7/XmP+ObrqG4Gv5+6gy
BISsVy4ZqADxK0PJB/RJVwYqJvhwJy7w3a89OfAPuuMkt0ziM0ZgPLSFgPgnZIz4
A9imAIjAYSfkQq/pRCnF1R2ftA6ifiX5ETL2A9jU8tN1Fzd5LjIlrlfnyJ/NTyUP
UfrD0lFv7/tSPQBFAfXpzPYZaltV7junfZAcEofbQgq13qz+GUgdr8EHl3boCzrD
NCeovbTgdIT4xJzPpeHNk7fvnGrx0JyhYri9/Ih7QUVT0EYbkbnHhq3pW7DhVxtf
8M/IKZCUQFEz1LNHZdcKuga+xpusMGPe9lZihz+dFOmLnd2sJdcK7ONBCzPDQMpT
iemj70bJK+/weZ3eS67CXWdV5SSXinxl6H7rIW+3+xwTkNV2L4JUH0RSxTVzFnNh
UdhDZxCyBxbxMvkqxXBGHItPuVVc5/A97MjbH2d31HvBgKWKMei9U3BEVmUQPJMS
ONP2uBku17+SEYL7pZJkcxZz8+xCe1qpln0BRe9o2fdKHBup+GZsghgrtyda+VnO
LJPH7jtzkzOAFIAZseRJN2rSvLvLUR6Tycb4MnSHR0EEwrf3d+FdGRGHqrPkN73z
CVPp3BeN6Nk1mSPN/0pXPPCzc9g1hrkWAp56DtJVToSeEPx/vZnS2rBS0ebP2xZG
UlzdS27WbghXgpDh92w/BOQHWA0j1SSgC4d4kLzNBnKRsXCWLaRp3NaoEzfLW5yB
3FPVqZ8fzyVfefcRKAICV4xXStNzvvzvyxh07UVGSJp5gtO5QYlUlQvTkx7wb1LU
WhmawTw9vU8+yodTrKZD0hkvjKOFIlRf9HJ4AVMU3/FOnCdyFcG6dnh7a88kd+HR
2G7mKqXstVOok0Fnhhx/RX+yY2t6bKWPKUWj+Z2kprJaAgZ776WCKV94xc8pQuCA
ieaYVPEX2w1eK8WJOCy5tbjck1IMnRB8+Nb1kXGm+LOJMk/OlqueZVAUTJD3g6tt
8cbOGlaB8AHj3bYBipocTSe2cM1GLJ7QbDF3i+VzigAPlA29gLjhtov2f6cYV85Z
VpXmC7GFmCxIKDapUvtIap79XqKM+vgYkDKclwIarS/IwC+LfyHiqBtZcBUYV+SE
ZwWLDhAN33ougG9SEV3NGyvcKAAD4E/TQtOw4SuXBfMZ6CjvhtqfF+hoQkHmXsSu
rM+TFiIp1pyNXYtDR0l/PxEc21yzbQ2Q4/XTlEoU4AFWKGFuLilkVVBIFHcem1tC
j8JrS6GfQHBQmt7YDkMQjqZRfUbbEweKqDejhml8Yo5GkVqEuJyfaVS/zL/bTCMP
E31KniJK+o6hmcLX3q7+oedr1fdfoo8rfa1v8MoRhAdHtsSwUwLuRZW+KoOwR9Te
ADLozKpVu1Yd7sxBHzwJyVVAoj7ZgvnAMqpuJzcRUjH047sjXkWe6cDED8vpVb0w
fHCZEyS4ko2i/wf7GcX8gddVKhHJmyWBfKBiSgWSxZ8dnWvcXMmbB5zN8+UtxhNn
r+sMmEKmvMfOHAnr+9dG/0Dtn6sCVtZkPTliuvRvsBjBUPlXxe+fOh33HGWaU8+l
9kIdO/MWDl9iVhJRXq1ctI6diT+PQS9GGSuxDRUfaFiAQvtrHzcPJQr7xYcIQ2gF
g587kjRmLQT58dMzXTDW8LVDTzM6/VvNllqId5C3tVd24hlwMSQqD8qWayy9Tu3i
HR1uM1HgG6HaIf4tcPHrUNS9cCsNyn0vXUl9G83BsTTjKaZ1feXkl6Wy6YlZGFkr
NEAEDdjLGd6FBCgrRIQOhzQO3guf7nDR7TLljl9gKuMI4KrTA3Fyx3nxdMyzj/ex
ChWQghWoqa5olac+E+nElCASOzBMyaYvE6JFgDordJI5sv1Ftas20fBy+4nkSFkk
dcLK6LnuvWLllYkq6EGRxyR5wpXG4cmncWEVVxCZPTW+gsXawy7hZpD00q0tu4X2
0beafwNs4Yf9af2q/D1hojdN8ItDM5McShp2MJFoq83ibRblKp+QR63vE1JSsuHJ
Y5Dl3WdAMwoBur2nkSeNWsuXNjjIv47zcySKNwp3ILnCAC9XjXX26/cRBm1YlPvt
fd616wArFTG4t0l9acCOn8mXnf90G4z+w2ml3Aso21zxgfWAhcHxj26RW1+2DdPe
VjlkwNfuZDX66j68fLQlyZLFF7MwN8bL21PVwQOg6P2Y+bApqghBQz/BeWgz3kpz
iNmf2BV64Ti3S42qlxho/VfJPzvVNU33xY6hNimgr07RLmqXIKty8XjrstCOuMcn
M2C8U2Tzrn0YeCB8Yr+hFLNJBlxsj7Hia7bQTpL7LnHYmjmgm+BAh/mvCuzRq1ly
VlWvRZwMAFQBlo4vckLPiVk6xyP2ne6OC/7KP03dq4D4ZPJApCt0jyPtMZRW5Vy8
5nJ9/VEP5XJLLsDU2vEHEkGee+lrl0wXKi/2M+SrMKK0DuGdJMtLBm92L6N+wJBT
omVdyWj0nD/7Y00RuCy7M/1bamWZ5xEvW64fq+Hw2JTiWIiOkGktXmLPuCyFIKrS
TUGQ94GVp3GCzFzoTfWrQupzoqvWZnsMb+kslTGjQglFNNUdIgH+h2fag+7Nj4Jp
3IObPJjfwbdcdpfzheZoU7VquA9UqILOHP/9B05egUYTmQK8EFfWzv1pngCvkIkt
n8Ql/2sbNl5RSewpCcKAk7SXDx3rdKIA5Z9beHeDdLmsN4XfIVD4K7Sv6rv+YG9u
u/MEzEgyiX4SMkW0rHTgaI9KY02cDbjczxlshOMs6ukEVgci0cKFEqrXCSsWRx0p
CvHv8yq6VO6+XYWiNCZ8ndCD22F7bHlDA4qayjv0nKEfliyMKp3AKcQUbz2TfaU4
8r8gv/SSjrNcj7YTL1tPFBsYIu/ZKaf5dUS/RH8J0IAMpx2oBPZbROxORprgEtGl
dYZ++6Z3etzMcfUf8osYXiPnSjy1LulyWQB2IpgHf3jXE7LnNvX7Wez1xTam36eO
HsMIx7Hh6aEv5Au02T2P9/ZYdRHYaWxz3AfOcy7UnueKg2GthbahDWzBiSHc4FeD
1gWbMBVszrnVzcEAaFkPrNUldDBlJtsnd5szXRSgDet0+1K/RDVPzr1SdTEFWYei
m/eKu7ntXBePlNlOc//JMd0iMcnMnulNtpv2rl+rsuQrw6vNfH9reLbcwIoHSeKk
n/X3ht1JbQ6eBE/dSDlanYn2PSASGDGO7wOSwHfp2u4LihR8vEVxf16cDIPtzLTg
rEDryEmS5Ayo9mQYMoHtpB1tam9PXCUMUsZPzKwVvEJIJ8bVx40gZOvBksVP4E4W
x0KIIFgeqQCQCvnA9LQ9kfFL9hBrdDaWGx46DEjtn00mfJemN519CYy2vIf0xdyd
BDtrR7VFDQOZEkLnsesRzMrGlPkTaLOXQIat3rm7PpBvBwB9sC70xQj29m3m2vE9
9NHbfH8bBajA+1Y9eGN0pIDkXxG1xSAKVBYRlY+xl3qhH65BB1Vo9olql3WJlvo2
fy1HLIIjUwapzvOMxulr58g9NnNyBUUpr+wqksKzjpfjdDOiHrHVxwXJMirMm5CV
BQh8j+FFSmiFTV/QNGGvUK3wQNowwjT/5jstNABZFPKCefdfd4NpQrSw2QO7pGWI
VobJ8CQ/zdOKwFJboLKUsDzIPJ/zI1YkJpnTWYm5qoi7lsvLJ9V2QRoJJ1lRmxFH
I50V7xqtr1/MhFTyjkl7omhJePdpnb4hoqrJgqjvwGnTuSi3CMjRPbIDx8LBrI59
hv249TDcHK64LLo/23nzNcqt06ob3/s5URBvakly8MCXIRF+iK3Xl/oqi+CtRzue
yV0kxRyFzv/iBlfySjzx2wjj1ePtgO+wh6mxhyDuojNDkrdb/jwUcZxiZpWfMrEx
aVa/x2CqNm+Ymp1raCY35qHilGH9lpdV4OP6JvVw3FDgsjLwLpIsbK40dBE9bTu8
yH1JbuFasPYgURDv36z966gQtIROFtqaJrmf5H6M8iJ7qlye05sI6SB3QgjxvFHb
nYVQh40o9tP8B1hg9Sndji/Za+ox88CLW72ZjlfDso+Qd4hE5wkWcpMyplsqT7m8
wT2pxz24bM+8zKCExmy36MlbqwVIVsUW4Hst6UiJ3CY/QPM6ebBrzzjAXb7jSQw9
Mc4b/Ko2Iety/TShZN/5mhfzyPoG6cmNX2GRI8dCFlMo6f5/UD7ptxmbR3TBh/fK
pHuun2j9HHzOVosc7w1FaJzI+q/2cXkj9Si+At5ulK+EuSrnkDbuYgPFWyhVUmSm
tvgyXCoQuZdEIldVRslsWKFQ6ufmxZXiAGkYekfkfdgr1Z7j9uZMIJYIvLV2Ro2j
fj1aaWb5vnTpAdEdR9x0mdnbLLEP9/VVyLMXngY00r2JQP+bm9Y634O9E+LW44tl
RrvcecpdD6e+lmZKqTtI5fKjhNz7INgFD/Xe1FEj91Yc3ZYG5/LhM9Wu5Vh47iKe
X6RAS2X36C/OQlMjEgGDrMPLPxKrpxFqnZtRKMtEdf43m/1b+35rciIf0flLfhTb
kPnq9ZZUBKpgSBIh+VFbcy2NWPbujCImh4/ieemReoQArpAzmssWuWwGx9nscj26
h51DD6NdcZ+k+NCUdemERC6GGs+kabIjxTXsWIAEn73cWMEIw2lqdDzeBxKb88EE
wiPwp35NkICLmzRXEKfrp9MXUoWuEenxUu7I4NKtmw7sqYaUs9J2ZlMJuI4Flp3I
3DE7l8aLY3xEwdRg2r0eWvJPEU37xSBjUTOtwSYdTorW1VtTjQs5tO4zNPpEZvfX
rS6FfrhCijlMnwsXkOxecYAxg2MEU/nTr5eVrD10fKdcR5RasK6MnSyKBIKDpVVq
sDm5zkxhswl3c5krxyBrGiIBpkCTHLS9j0OlXNG2P5FurAYHQhw24d25nMlAxxqI
zM8p7Bzp2naQqQezNnKlt2aJ+zqKJeKX/+uCVn7FHnU7oSrNbBf1RYsTKR5Uks8U
rgT9pINSFuB9zhSTSaNLShv7iSwlZNd7gYZmIJ0t293TxUrvrqD0HykigGJHXPM4
kJH0l8ysX62YFNZlWhyXSZTAAFVChMlG4dI3yOff+lYru5odO2st3Mi50lz7tZxP
1qygL+q/Bsv3aE2Ubjx32UEGaR3gT7E7qLcY0UZNTlsdwMaywvZUqy5fY09qZhVF
oFkKEie3S+O+jKxO1fSJbkWmgSI4vJsju2yL8gQZ/TOPl9Bst1fFdnVsqaBtJJIz
SQqwpJD3CEcBVCmlPyrdZZdvtXpD07vnpydVW8tguxJMr02JuMhnGfjbnwa6Qd/Q
vXAt89QaL8i3LZlefkt44wlBmkVPXGBZ6PGr9zCn8E/zE4tksQqdTINqS7yGFva4
tchhMa+x81ijmXwlqR72HRfDoQwsoCE36aMKUT6PEYrCE0isRBZltz+gAL6YxsYs
td7bNGwy2h3LkQgPo2fAGlthuYXxwXiq5Yw5Oafbl5+i5hfn0ZAh9WkEQkC8cUHb
m3h7Cn0W65PL+NzJixN8FEI8Y8juBHKpLjrihttTH5fg+X0IKcmwbSfQPV9kwiZU
HHf0SuVzeECu7Ga3mTMmT1UQGxz/7m1iExvdldhDOv86VDWP5n1I4CmsWYqG07TL
grcJYj3b9O4F20BCkEVkVL/p9TTohHISB7+YYntnuZE9pzcZUtbuG6g97Tacrx5l
nTVIdCjUGpo5yZZVF22WlLDjrEZYouwtifGlnI4sM2kz/TEwtxk0dB5udGpIfl8n
E5O5jIxO+XY9/DfwvbFRGikrFJbY2qlvrwjlQaZ0MdUPvHky9Urtk3lxttJK4oz2
pdYCnJLd3P3U0ra6kJPy9LOOvP61sMqOboSantPBaKwHQxHZ2Y4pat74M286X4Ys
QISGzrFNL+dozdk8apweBC+IE7FgXW9u+m1Ju9LlLMH+2R2XR0btbH922sMl6OX8
587QrnKOoQlND3jzSJM6LzUZxiHwxNcvh9McuMQN7/Krgbu1QncYv9Q/TsDFsABR
bM6Jmp6WADUkSDdwJ9azp9bEFHcU8ZEz3UIe3qVAe711w2QWnmewoVrtuAIvHuK2
2qGKpxy1aZUK2vRVeSxYALf6VLakTkg+AHSK/R1+RW7Q6NNfuQzX6FITUFXPQnUM
wBFAZnqjlrLae4W9dEW/lu133jBIebOVeCWu9eK/YFRKaDmXs0DRvMFgBwn4lhCI
kNPb3RSk7O+x+IOh5TDkPwpn9CvNE1Qdy2mTPW7HX2bCkchTszf0coA/96vTqIZx
hH6hlWIMVMcd0JqxKOPZIHnAeoeSFfZZJFRu+A0r02A02sFkpwaU+g4XaSC2pEIQ
jt+yxQGtka9Cb+i3fHK3yjAI6ATEZeeMc5hdH87xBUn4hn8fexI3KsCDkvIkC68a
6c9RsH42AGgzjS6RC3GJyMccyH4qHYGEt1ITALppv3pKqqk2wgacWGLaMuj6xkPT
vyCeCDoUXI1a7owq0fbowBNGGPchoUKs6RM00+eTeHidXNVVZWStC23/pQvY+EiV
1AtWMnmkvNAFNnTyi0TjfS+gQHDqXQ6ekU5sEiWlcMKlgAI6AwLcOXCIxhht/zGC
bxgYDOC9Y17C8dlQ0gcou0ZalfYcjaaQduNNGPXD0SW6fbrpHtpl92eINUcK//Jh
0T8OQoyhw2pFYUb5NKBhtgm7ZcHGPZVJnCLqJGuTE7frqaNkhVHXG7pQvR4siGxk
LAUs3nAc3yXDGBF6zIMBLzi7/L4k5+W7dviOcjCCXxf8xDsJWyPvH/cl+bRhH7AP
FpqmCeX+xPpyRm9ZkJEv7qevloLzh8Ar5Ce+FsWaxNGgjtyxePr5/aIEqM6WGVXp
tgU4VAJcnTtnnVwcv9haP1LjJaRuiDEi+2hw4swjgwVlXNM+qbv9wn8C1e0XBeFI
E6a4B4V1KjSjNwVaxt8OCwuROuMVFAWX2zNltqqHTsDIXeQ+pK0z6nugMfCiS3qo
m5eXmIcRwvWrlm+DdPdoG2N7iq7kgjHO1r8wltOxtNzA5jwVri2WOWb2fCQGM22Z
8QRMs2QToQvmxffV4fhcpQYk5VsnFJhD7kfaR3PVRBtF+kU+K/QEDyeJDetWd6l2
WC59eHVjOZcGyxKWel/vYfqHDKc2r7hwCz79/1OwQph/ja9qNJa1I/43dKicy0Ak
RcFSe5rAVPuh56/h06Aw8Pmx+Y5IvNYpkOIXCosGNbCbBBYnQymL7gkwRpUecvwn
q83SJm5w/Hu6vMD7oF8QlKpaacQP+F07h8iOk2En1RrSe1KioHtdRFdTJ0ECx5pl
sf9PIBhY4nTMeGAn1EpUExLrTdohwlUfO6zLCFBr1xKdkrkISrz19J8W+xHpqDVb
KFQIAOBIYuc9DOl5RvDkFVP8cF4vY1qGUEytqreJncY4WYtw+uwBRV+/vQ9cn04V
ewK7e9vqbnFZHL0jTKSZxfniXTc8tCw7kjfSpetul/qxl2/VOviBpRIaUE8hG7YR
Aep08MMVb/I+RCiaFTaUoAFtkIYazmixAoAHRnJAOYnf4b9DnrgKWmwv3TZDDZEL
GHmh6UA2pV44BvveYA0QpzSHfxAU0NDtXEwTxog4CrLEgIBhjjPeFynqyyAt1SMa
VMyEEu4VHerqQkgvnf9vwSE7gqlfu5QsMqwHdRLctgqhLImeAqMcl1ZgzrJXffAg
iQxS45bynMG1gs+Ha7ytjRUGp93BhaxYI5QNGAa86QuQEaUVzabUjm1krcA1DQxR
WtRyHEIQmFjJo5c4SjsPDOcS5/WUWldAjBIkLiR8ws6/ntEoqjvGkqYLIogduEBy
QcEPJvgjn57VwAxVBxqogyRMLDBagQFEEC2OSnR6LSxsBIfgLFoAeIZFCuE7zmqU
K7knP4EpSqFIXcI+NoNrz1TKdfIpFnMZhY3yBCZOffRZ48zmYfKnScSZ7sEpZ6zC
51oL089FwH6Rniiuk+lfLpxtt/oUl+fqvicf1Dh07+y5upgpPHH0S1jJKMDvgeJU
tp7aurqG8KmiSlacEAbxTxqAihhZzSfylAHW3lnOTmzXXCjOqmoxTstC1fUnTUS/
O6wUZf7fpuKfzF5k6nsKmwEvMOUtWcUtyTXRQTgZZ7UF7VoIMv/UV5gEa0qj+E2g
y/gAPuiVtKGVVStlHwmg5U2OQzDmqjwa3/Rozuz65b5tYoiFdHDmsNJz7rKt7QqY
tjT/ZxkHOzGKWJjhLMbmIjBYpW8VFJTvUuyhJK5w8oZOhF9pGUkOEY3mWyhRPlwD
FnXszXtxOBqwUnw29oeYx+mQjEs96heeKuJpVNvDwR2WKqQlIVXz3m0fnVjWPUK/
0Hf/td3yUZhenxS3RqdN8vAFa7qN98788MHxR2GeEAioMREoKq++wU74O4UY4MHO
RrpeRAj4bukyBioA2ANo+6JB+aGJTWR/mP2WCkMamXR/3i6iPuNSP258JSTQIMVE
jXnVOV5Un2ipB6/PKM1khFEPY42k0P8iNC4lCoJTEcefcPxoSFyjmzfnMc5/sV6X
y9aL2sCnb8QO81GMSDWY/D+ZjOxXdKgyitnBtzMhfH+JAG5YForaSlGPhU4JWmKS
xD+/MHzq4HMdj8wWp96QKcpDB0FfANdFK/RUcR5z9d7QTi7HKAFM5fazY4fXJsNI
6GNPvfhGJ4xETBPc39hUQkqB/zXXkccq9EmXCSDk5ymykt2DW1yFFqjBYjTOcQoy
HjsKD/n19ZyV7a5iHbFdyzRWsJjkfS9R68yHifPC0SukU9/HNtIoKr7dKyIh3sc7
bDhsrWTa17ImtU2A2s8qUBCcetlg5GDI/ctjDVet1CJ+IfBOUcANv46/OTZq2QhU
JxhHzorYqvlcZdyTmgw2HRyoymN2o2fYlalqCJRyNI87PA7Odk3lodt9qZT+wlkS
EJEJlJIlC/GbpcwNYix25ca3fZAsJ2wFLEccXHFPDi9kxPqXwo/EnHzfbrgvA98z
lkuk0P3bDZQWvQj1wFC+af2+PVXZLbniQXVYAXrGJjeVMNdaKTM2Q95DccZNQ1Am
zfy9ShbJtSso+aUoBeux6zVb9PO8vYW5wwOfGj/h6DaOHKBpF9UTTvNpGyi25/2j
FRucUElu6+wpPumwFaNXZmtP296X33yijt5nb9z3tLSacu4ARzjrG5Is6cxXtkVL
sTLPtQjGj6wcCQmU7TFnwSp1/06kgzYEvEkTXmUD34vINJrkpaNw7kcw6dqiQ+gH
6eJ2qI/kdheIjEMrlhcPiM+D6/B+ZdRMeQCYKt3VdXd0Gd4RxwXDSnMNHte/DXKw
i1KfYjrGvXZDC4wXiqZ0tBN0omEDWSGb7Q7iBIloakBsxJHuUXTLGxpBIA2U1MLh
uTsV7gLpCaL7naGgJ9PEBlNe+CHwb0PNHCLffN24g0ngph4kb9FVqCl7ktnHAEs3
0ivJXRaD/NrUJCNyjfC4NkL5tIayFysfCiXF26nEnDT48uL8KSXXcZM0YJKX079M
v1B/KCq5kyZZdhROxvn0zgjNykkJfOdg9B5iOyDwplQ4JmWMVjteU6xr8XNL+wOE
sB4qFHZ8xX7uzGPULX/QPZ/7oa4gkW19+jTa5EoYo3tfsFtQmd4axbL26COlqKpa
/wEqYu179VOJnV3IDOTwBU2N5SfeP1+Lg0eFBVnToXve8KzbP0n9k27PTtBjIPoK
1/DC+CUYnDvQotgbzL+NMohIFRTAzvPNVXaH8KWnvCyifChD7vaHC65FAOOoDyeD
FLX0NlxRtsulVRY55CasPO5uUXV6hHGDpGZr7uQW4gLNuovBXBuagg5BXC1W0U/s
pZNCsuYBBXFbiv7astavcvek0hPYM2Ceej0dPJH5OD8HWjSlb/555KFQKFD3c8p2
f2MMVEntkaXrToIexxmR2Cv1qGw/zt3zB8h2ekQOPRdKW923MWzI5C5XkhHkJ6v2
6NRtwZA2FygOhrSp9Q2p6vLWwuopsoG04VmaLjSBxa1gRLGWosCOGgCPFk5OlzL+
8YJ+nWsT6xvpw648Eese/LLi7tjL/yRbA7kcWkVUFMMduZN7SIplCrfEMnzCH6N1
/pLNqDkVicqZCuWTtcPubG2BIDz+QpmAKWUuKPq5qTXio2ScdtJCz++IZFJ9ou7E
c3si/gwQ7sH91EQR6mLFjqsEfw4MdvetzFz5MPjJ9DT8XGTQ0z1v9UY5Kc9EPVZg
alrp8ryhsJIxNqDb4/G8apbDIXfVC2/1logiWTZb48MZrLRv60jDFFX6CIh9qrVh
cuAbD5dZD1tkEEr+a171huDBygUW+hvTVSh67Pav7fQWYisX41nqX+KOkXyAyjSd
6tD9cDptYFDXs9He0kRMG+vd44jyJSe9nIGAMe1PwgVYaivbtq63hG1ggeVoo7OT
AgWK98PMvLEWUfUa0iPrVbXb81DgwEIlQ/OocoKDyfeJEj5rJzF0ns28KB2S0ytw
VMDb5aNzmrYiIPFauuOR6rOFoihiino8xxrz6x/vMVXsz/0zEdehrilS//xntvKX
aY6Pjc80txF3I/Z1Zja1UwNGComUIhSL9uNJvzR/ga5JYJoB1uZloVfLrbk0gZVf
lzDrouG+jEojKDzUOfF2mBtJyqc9BL/kG6x8gB0VAe0ekipE//jZeHbCFLahpxVk
r/OgMNz8bbcBeLYV7JXkXhSXHRc/oVzUA9j0En8Yp3eq/QDjsNs7n7YPFXIm1lHT
EETDYqA4Bd1eIA7V9h57bwdpNkpvv35gmI4u6IDXE4aAV2dNjDVYbwZmwAmf3jhS
hF2I3PRBefiZ6q7SKRzMo4zKXkw5ZunEeAWfXRuwMv4r9i7Q0osLPgamQLr72MOR
0xYYQYMtAIqPLx80OqVx70DgeSZrEH1GnnYxAPJ8ef51QpdNSljgTr0AHHe99+gh
wMHVrsqPCv1AggUgw9PqwIuBCXCagLLGL99do7mcE5rSTqSZECS53Uo/CEqlAFw9
TV8zqZhsMDZ9io2MM2ACEJttAgMvOAF0B+bbQYjWF4tZJsDPWnqWv0osLXPEkjN4
as05YoUqznYXuS4QennasIRNhfTLTD5vP+guCXunAIqzvhR34Y2GiB4okwBPONNt
XWigwxKdKL2v25iP1nUInMoPCR1MTaX5qBZ04isDRDqaad0frulHvrdmZd4nWQyV
N9eCqtCPx82yOEekRaxxFJvrCfjEboe3HSh8yJ3b/WALiRF0qnwCL3+azKzVJx4a
l/FuTwHkxmL+TS26rqZ0fpCZ+xXNNFcYgjZwJDuzgpfF34QCPyDFqM+GAZFlDrmA
BHWLbytq/gHXE0C05cp/Ivdhijz++8mUyXV9Ly7KoZ8AmwUZGQ+EChAyY/VEEObf
osccki9hY+Z+RoKsKK3NVItSaxjMebSoGD9ccZZpzf51yW2eB6TiD6+znP4XmKfQ
y/6a2NT1pYxvBlF3k+NyLskL0jQHmkKE7qZ2ma3ouAo4gKXWNs6+cRZSR/OaNTWJ
oqQiIDZul8sL99zRrn085wcjXUu1V6RTILTobl0QU8ImJ9OfCLv0UnA4v3NnCcNX
/wZp3QlDNpHP8K779md1JIaaBAEHNVS4/GS2OuHN6c2TySPiWARwgsj7kmz8GWaO
1ZXv17873TmD7qqAE/n1GiYCjeejbXSSNcmW4+rUqyfW9QboNeXowzCWIAg9eXju
1sDSe7xURdONUkoOL1hKwVlk85tSHtuVyZMX88gCIkpcRa8G0CeVf9gRaC38+ipq
DbBmS0lC9ilZP+GRLAN6tSWLxel+ZKy0WSK+AjpMZbp2In8B5GiXXdzSdGCI83s+
TKSlpB1T0ScFAuciXiLctN7ANjMzPx3bc1hv9m2wn4rJNUuPOHGyGnpMmmtjd9ZV
eahpSutjBTxm3Vj7tUJP51UHgTgNRb321Fj9mpNCDHbxWDsB2UMHtZewB2mr4Ofx
bSS0SC74wkUE41QgrJnv7n2IQk7ArCDaK0GerSVZn7NmrC+XQM+3HRQRU5TgZuUj
G1medSA+7WjNZZICNUmrFbC5aBVCt/N3FYbmzhDfWnwivEOfA6Q/UOoogCdfWv+C
3t56r6gKF0mCx8HA5/pH3wynoKO5wrw2K32R87qQZVLvoerbOX7E02bceln9ya79
/mcOe7EwCMMnbs/vPhueaV6bO7R77pPam15+tqg/W6Nr4NO/13DgBTuVkpLmdr9Y
d+YNCwrn1xwDJmYT6T6J6+nuq6qM6Z9hSnDyoT9uIweebon28XypiQandEN3AXpo
ZwvJhNq0cEO10rv76WglfFZTSWXfq5d2GL0FBKy+mlti2jNk+Tf6SFzbKSoL6J01
+j6DbfKRd58OU+zy4OGkCkZpj0l5r1YFsjT4lnYrM57QayeTPrZFBSokHvSQTpVW
Ni2XK7NLMTqtqakG5XXPfe2LMoJby2YM+uq177Re7VIi2fhDyzOulHpcO3h11qKq
ZDIuNJOGhyMu6dUi2qzUFgLBUO04rA2P1SpqY/zj0JhlR81xoNxzieVO+/82IfUf
jRW3ESVXMWU5HNt4hQox61DoPUUuqF1/ojQsivlCrnh+jYaVz3to8bbtITKr/0Bo
gcXontT4dAUBXGLzKFFV6HWzTg7oz5uwnowVzm0c12UhrkktU1X7di1A/CQq+K2F
egWJalwNY42vMX+wikZ6Z1ngEA4cOIxVZ7iOdsbMdl5tkUK2QhT/gwDEDE8Y5VTj
VAkD7EafqhCr+MtJvBD06wQO8DFzpSeWKX/1ZCwekKImiQz+8kadS3wpywllc+QG
GSzYlOmkRZUrXG06bnqpTfQa/+zX270gT1zpO0B4kxha+ghyNGsr2kR/JSuGaLcm
mCzvM77muh9x51U0qGbrYyeb+TZbQPdiQt+J1XjWESZLXMhC8A8x4dsy0doTvzUG
lx0OPv303yXX/3YJ5xEWUw7j0ZBUFJbBwQiv6bulYG5BsBRaf3Wls5cZELhTD97I
eOVqU/4PsYqzlf6jFBolQ5rxEDZc5WsWWkBPzrfWpt6cimiykdSd9xUxft0iPu4d
CgipQgvEQony9MWLX1uDPbhIU3LgyQgOSfK31oW0wTBvsPJbXHA0csPBw+0PvdBK
Gwu6LWhNSLJqcVA5XSRs5GouvGJN/w7xdMZkduHCQmP6YkfPzDobyL/g28yoAZov
JG+Xwcy6+qfp3x+keCHOzNzINTLBk/u0f4UNNZtsm5vrlzQwvCqPW6YMsSdpidXq
fLd5mrkUTzChmX3tfEOmX4X8sSXCv6jbt/AkDmPAGOSeXJfLUMM6c1RffO8XSWhB
5t07fn4yPuNws1LDqlmaSzWKym3wISVgpWt2fsw9AdUE2v5f4iIQ4Jmu3T0NwA+B
ywAfygW9rA58H7gOceXKtFo5PC6fmjWNGNmW9Zb/7oNf2JE1rPqkpZqOM4djlHHA
FIyKlrWPyZAOCzlZ+bIe1A91CRTOGVxXvrxJTRhAQWeBvVbUfwfQKKmOBZ//KTPD
5gG4Ns5knjxUMwDQg24aNnRRgWUuB99wLggZx2PGhh6FvheqdZLODXdboTbcQst1
WF7L18H3eTK6ttWJ91HtkisbEaCPLLQqQyDCLWJbeBHaynv+zLfML4aUMCN3CX1c
HjMMhOCaNXcdCaC2k8dgTX/uF+UiQmVEchTfuubMCfFRBWqgbRpiWQ/uaELJxjUI
MtXEeMmMX9D90ld7pfZJl/3YEb7Cg266zyrUtYNpQQZFLlOoe2V5f4pEvgk/Wv42
KOUPrB3xe+eTt9MNCxqP58ydgwGSjn3UtFlU8s7hz+n9dKTqqyXfRtc9qieH/STC
620K0g72OAZrK6Xdl1W41/0pqDdqSm6M2P9uzNuk11SfAb5ImQRfLlYidJEwZWDa
i6L1po6Sc0WmwxMeZ+JkJ6ER/0zWWmPk9oPivdm2zcTfm6YF20HZheBjTRi29c6G
9DtKny0cyupJdawXmSUK/fFr3JKQHLrYL9JNEXyxTlEzUPt5RIaQXwF9PieAL3Oj
1RF4volbcNHJ77as1ijcR3WlIuLVXgQ8QqkfKRodbPskoKJXq9+qQNo+Q7uNNy4G
JuMhkjm7LafpyKLdx2KKfxsg5DRJ5XPAI9/59m78MCGnvo4FGROPtEKVCv9bniGg
YXl+bIHlZ4Bx73aDaK+0RAPONMYHGwxrkvVpGxsBkVZd850UteV0SO1KB0uiisCp
9626OU/PtJ4FwDGvc5FUn7xsBVtFxAu2aNVOLqP4oEf5SydfvE4syryBQQvSnw9v
j8luKCEAHbBOHDUYl/oYqIJP5APJNi2iBXGFE1GmAfWZptWEKorU7F4hOOf0arcN
3zqBjI4uqWegIB2DhEl+Pi6e2+Hwrc1UXvIPWsMukRt7rrlslililodGcPtdpCn+
ubfIRFucT44joZMfllD/YeYXVPDDThWuJL79llSiIH7pg/GQLUN1BnpaPu2CDsSV
37ZQJz+0Edr+S5dDfWwg2azYN2euTZkpJk0OiIrcJU/5W3ReTbXEMZ0p1nMb4ZI/
oanWq3maDRlYWNAXltg9tlKCj01WJI0zCNIefn2/Ud5MQ1KcjgwfdauKz6Y2NCUL
xAL+Vfjj1Kk05I3BlH4PHxPI4qOsQm/rQWYo+GeJnZgELmvUwCMoxqFqGw4YhOfR
YPLT5b4U+hgL9qjBNPvMEE9Kfo0zS4A2Eu/rQdlnqokuhZYCxVqpdOUDhimWyPol
GTmh56GKWE1Rovt/CxHFw54PEAXVVjhjJt77r2pWjc938loZC4jckq3kneK9/678
rF5eyUF7le5o9x56qNYWv/RTJxc7BMghUih730NSMrSRXdqt+C/bELo3pr2UUEGb
momKwga0UeJzWMkcDt4OgZPYC4aee6PZwU0lei+r+29N49KT4V2WtrUDCvZPqcqy
7yMOA+1JBRsrp2tXnFQRvQHGdeiLSik51va4JAXBBUooIMcKKSVkXwmr38AIJ8Mv
rejhV8lJJKu9uOxVGvKJrbd8Km1qGwfw8JKGbw/15T/37ZnsJ9JTRAJQBvI/vXFb
NfRwnWkHshj0TN7eC/LJj73dmgR4wcH1NqK3wSW8w4dLipy/uW+6UTviMEn8vIqK
tTKsqKcbTTGJbC4HBhMXJvaXEM8o3+0HgLkhXVW8jtpx3dKZDtc7jS6mtrfDIQQz
8XqiKYL48p7tmO3OfKKThqSpIY3sNZ48oDkeFT7ZI2CR54AvCZYjXzD9EDnRTZbM
zlvSjcbImlVnwm3qunLz/zS4Bp6au2QP2D5vHFxwGaBjEAv3kNdLAac7Jw746ofN
4c+cNUIhum9fYDfvAkViv1e+hUXEdBpl3slEa6PNLb/haT0jZehDhqnv1Cr4R5tQ
uK5aLya3h2IzLry5qvNy0CUWWuHfKjy1GEz59xwV2KALA+E2eVEbPQpWffnFczbM
xE8qN5HyVlMf4rjewlK003EIHUjrKs5AMOlawjs7fo+8fvBmklE1g2GrtyjbXlSu
ED8+DYbAkNSLyYRzs6yBo2rFx/zh6VcPedYUFFCBtvyYiRz1ipP8DaZXVeMs441w
Vfz8Ru7tCeiN8IIkNxSiVMv3NCY7XqPuAmIArAp9PTSclnwi3LAZ6q3DIpE6TkRz
qevZ70CNvzyBAypI3P24781ItBA2I6FFVfZqGhPfccsPAGugfg3x9z/DGu2Ko4//
7hlTuYAwhWIevKdTG+j5nicLKmwp6XvXwATWdP95oGeWjBWUAkbsiMA772taEGOa
fVHN3GMcykZtyaeIBzR6NDbEhNKGKOebuMEbTvDQkuu1olsevErGnQmzMpbTGelX
tMk0jbPPoBrKGGMXDF5WG7G2uz+8O0bV6gxKrqBDYJAAR39sGo+0R5JNiKGvnJyy
s/9f4A+Ldh4YFP/xPM6un7v51I7fYRp2TX4xSyw3TBlb9YeJOgu8j+w9UZBy/LWC
cicXPJuP19yr6zZqStWFLsCbh66VzCwTuPV/xWFYc1Arp2P3IDNbTqxDRHhxJEQ+
k/VlcuNcw/TZTyXMs6g7RQvGy4LUuTOWPcwVdI41K1IWhmDHjvUWogijwvi+bTJc
hNFrziuhhgEDKK0OuLk88gIE0SN3zCThmoyRlQy+tmHqL9hnwofg9dTOlCWzOfHx
tGP40OdPvlzGRGo2kL6xk+VMzbG9wzq+zE4PXdYED8HXXJFri9e9zFgEQYuBo1fi
ljtal5zKn1TA/+k/QmBprk0G3WcwJFFHlhRUQ7MR07tRZBfzYotvKsl3ufUornBB
/MgZyXNKCReinmCano9u1QWkAG3JBWw5aMbYIG4LpJlmdAR0cZT+RYeIsEdMd7gr
EDFctXaNGOrM+qz3dmxXx0SRAtQl3esimMiuORtRKXWWr5ZQspyA1BsxMd2Ov4QY
nyega4acnCOK8q6C2hJvnRVAwzlxVgCwzSvG2+6Tb5LX07Kd/BOmuqPvGs7y1XM4
JdRoZ4IsqKVNTeYpb0j2GYvDBNx6GvZYld6W12hh9X80m0iG4IlGFcOkfpibKXlR
NpQWYeWXRGJ3xhs3ioKonyO6SUg17BMaS9SURtvzYaHIi6SDF7RAVVFIvEjf8xxW
HGIMKrD1Zlt5l95C7C8vKZ4D8q/Vp3R983igLedFJ19e3xP2AUVcF+OxlF2QyBS/
Jjjx6B+i+HjbSlJmy4vJ9MYufsYwKBei/Mof0mpGFWw3PnKUp9pUz/dWO8glgSV6
k3pIZfQfxpK1gRMpA2BArAYKcdkyUVdB0RaclG3F4N1PbCKqj5ySJHJXEiIrKLhJ
00JofvzvI/aVcaul20ptvtjpyJtyaDrJa9USXfqMllStbFYZ2+TxuXrL83+1XjgC
vcIDGx7Hxwas2U7Sg7VeNORqI/hNYBqjQiUsPieYGe4Unld2CLmEO/gfenUSmT4q
HlA+HISNwcGECATgSLmWkO8UIyjqblTE+ak84YrGEt7AqV/2EobWfeqm4KkaUeln
tv6tHaA1LFV8yfano4R3eRsnB+UaJodEhaYJ0WHvW2Wkb5IGLvlsN2o1riXgMs5V
0yZUfv0NldU4ZKGDJsrk/PGsdZJ6EaIuGqLR7IXCGNwkDDZM87husjdEasgql9en
tmKA7YdOPxvNFXEkt6dFj8wntkW/sanayzjAYcMnE4FrWBMJ4x6FJHB9pcDapD82
2rs36cBdhR9q2JKDXKcnOJdeJ/utt7I9VWtnXR2OcjDBKjhuRNHDYMUUvPQHOcQF
yMSP40gr8MsX5GKHfQTNvAMJXRcV2salhZJdoiEoCVoUXIKpJH4rC1SpLI2Er7oC
HYxlTft5ccFZ2MuEaW268t0qe5CNymZ0xEyz1Nms/ypkrvWwSRJIAkZDrsiuBx+z
6n03DA3KcwKaVDdWlOgpVCa4DAEw7IFOydpT27TOEh7EsDqTPuExR4OEoaEHkaXd
YhP8w1VlyKo0KmM7d4C7Z6I/puYP4D5CbRfjWThUM1qItTO0DFGOJIIH9ailDKT+
85JTFV3yjE05Y/s8JdUFk4UvEnYnOEzasxc7jww+Szluwc64CmtxLY1VIVqTMqns
u6MzZsK9HiCsHOndcSpodL5ybYuQhzayUI3w53z7XRt/T7CnPmv4TONkv92pfs8Z
8VpH0gfII4GLcuFq0ica1siBM4XUUb7k69NNH5sDseA/J2vT1BxIctvu4XKxDTVN
jl9tiueZ4XxiAbCzCiQ66qLx4SnOo7SjKZ7u0Q+eiJyHyjjARUexiOZwfxi0GrBg
dOKprO+uDR1zlLtrceHfjQ8e/IyVfv/2edN6PKJY1Gii5+3Re93eMFbHRtpoyxZO
rpeyW9rlliOFMvHgUqfDc5YGzdjgHjv1aQZij9ohLEhm/NyO/W53zxv+StLBOnzO
oHjwZ+DaHaIgbU30Ee48g0op4v8mAX7rGnkEs3D2r9J3te2stB7jtnhP8CuEJ/zI
aJN0tCDM3KBbSqHoJVpEEep9jFJpS0OV+MInVrGl1DQ9rMB9BxP5ga1Dhj/CW0VT
79kvWfuI0pccsKUalaZFh1vr6iFOP2YcHJPGW1Q2yBvQT5kLtAKYz7aZGIvkcLD4
thcr57J+q+UvScen/iBqAr5UqHoW0OEwYGPZc75cIT10A4WbBg1ISF+1mNaQxEYP
PN0MmQjRRE1H/4snQUQza97Us3m7+pB5KS+Pxe2CzWWQsJuKtmcH5dYKgw5BoOe0
g8SS4R9KTKGOoTUb3cAtZUayDBDWWedTrXnwuBf7EwcQYHbevXJQFotvSUm1tTlC
3qN/v2Xsz3CdAuLZsqtEdmH6QbjUNZg8IxTQ7s0PuKzPHMnMxkHQrKshDugqk6nW
N+Lz/jbwDMt1flqoJKn8hLhCT3GO662X5G4JaQ2PJU6lsyz/uTVO/9Btk0KEo+mK
t1Pb67gsMAe8Jhs4Khi8kuAzVKtyC9cC0QIRb1O3JkiA/35uRTDOoknSHhDDbbVQ
zNS6ecs4Cienwf8xj27KyBqRYW0WdgdD6OAQm2BpCHgvLti2JVxOryibIVK64fAO
fltfEJaMcuEXeH664GgnvtdoiUTh4fdFQdzL9iN3xN+MNwyKvn8YJkxDhjR7HkPL
HhJdgLl0Pc8P7ToNrqWMyhUE6yJSiO9fWXL6JurumPjzxBV4IpnBZdErRWhi5ZKU
AW2TJwlj7XyowTrvf0vwfO3mgaxl2B1FJadMx1C5mppA15az+wwnNlh4bNXEacXV
39o9U2KaiHSrAOLSsZIc71IMK92to8n5UB1r2N+IxKWVzJ8H+gsnoUGKLn9wzv0P
ok4qhPOBqftBbSury91LAhY2oB9+Uj7xel02r4xWn9oWdIDQproi5676lPitnbQq
5qMPh6FmHibwLgYFUAwMXdIjv1TR45WImsoQOJHQH83cKlZJbtv1Ew8GCtiecHBQ
Fs8shNhGpE3ftq1Ig3GoMWQcesYjPMpShGKb66wYk6eMv2wLksvySPL8KDaw451n
BZULK8SzQ+3hqGV/KAzbCpP0e4KM5qdyhrnZNmKh7RogNFFagaeIYKTcTirglD3I
RzkT2vejuXgwpAPzGP4zjnZTSZ/pY3crvFzE9ZCbwW5rkKaxeLUyRWaYrD6QhinS
V+P0OTZKWTwiKNGzgbDWFXk8f/BlL2zcZftMixggJFchBqM+8pSHkcZsNzQUJ6kU
iuhNcCBh2JvahSTGqU3HfsC5aXLX01QDuIatPru9miQwDUhjE3E6XNkvY/Nn9s1S
XzBfntILHG82LKMq2XPsBMVAb+96ZIcnljdkDqGgyYGa3tgNM9qkqU3dNMV1mJgh
rEIKft+4kTD/zJOliCLm629Y4LpQF2D5jmCOgDKi+hRRqt2+EeB3tTv2xE/CY36y
Z5hScAFQCAOoGazuCG6f6GEVopYQJZ9z6zb4ApjMRlIfDcG/pyQJeDFeMRQ4MUqC
3fXpB8Qz8Uqaz9a4ISGHDaRxZvReNxtpvWUWGqjGGyq+AGNPZIynzsRG0wnFcwwp
WFc3xmy6Zchlnjaen0Mz8j4QxByEVIQDWeATaxVbaYAgxB+utMIQzc6yaaXVkv1A
nVbcg/MdAyKcwU7nBw+gLG5NzLW+uMvoP+hGL6BdzEqwwTbGNJPSX04R5Zz1Xw8B
bC0egV4YwlaT7Ar28fdR0zr+CMlP8mzIhX4tmfUuYV1TdrSQjHp32CwSVpfRlzBs
Mr1nGUnp5s9xGqT8WeHAzodRuOr3nfQeKS9vpaAzTAkr6Fxe0KUc/xcTOdl/SCP0
9rJEUldLZnJZtHyh/H3qXx6eJ8LIsn44uoBHCLb0adjO4jm0gpufFtlq/C/bTSYw
fnLy8lRGTWO7SwiQIqf9/hEx27jvgzOwcio4xAp4vkRDyKfX7W+yW9BX8masExv+
93lfCrkrB5p7rL+DEPwi2FCd0C9o3zmjiFJ1SVBDQEe5IoDt2HbIl0ZNt86mmxfu
uP+PfJgCnmmX3VYYLP2lcfgfp0a5vxmVW5mNl9OWIxHn4lOiLlnTNziUvzzlwNzN
CW27wqR5DAMSSaM331Sf9rSz+f0fRgSH7BLYhG9TIr+NAtI2bRxt6BChH7iKH0YP
lQu5EkizWsaLlYNLk43XQgPV2eKvLpwKms1UV7FmeNYOVYWCNRFX1fHQeeotiWcv
H677BKNxaaj9/xKolRovFcL1KFFuWfWfZ/JEKv5vsYUVnbETkZeJcPS62oE3QP7+
9zO4UUoApOcobzSxhybPwkAVRiUY4reLto55rdMh+47EqmGVdBjzrZng0PiyLmNN
C+FCiDlYWO+Zq6EwAmYKXtTCbqavgQB9QyBuCanIcGGagspgMSf+5YBDDDi8pLaS
/vQd/Ve1b8T1SvkX8k4IBEYrmrDzc11vAVL/+t9+W1os06BNyKLb/fySdwrLlcQo
u/mQ+7LeyGaVzAgSqJ43lDB82owiO1M7TRGAYKsk3heXn5h0yQLt9S/JoCydjjwn
yuU7crWS1oGPQquP+/qf7ZesnfJftb1jDkBzVB2+HR5ZHm2aqGDXVoIhewcvPG2/
HODdSUTWjuujYswtOU6HK+yPiVk/0TZ4S+XXOj5GAnPIHH4tparNHQyao8SzVzar
tdkzRefwuC+5AUiyoR31Iu4QVeNDq03ge8YR39Z+E01awDbpGDcaIdvVjGO/pBRe
n74XtwK/kjNfhU34JUppa9wlcxp6S/Yv9MgjY+C02zEL+z8bG134aXqqJjdJfpQj
nBuY9EL7MUEs1OS4f3KCecSC6ClMO8G5sNwHCL9ku39a/muW8sha3p2PZP2AAYLo
sXyacWFEOyNwUN/40TuPXzTWVuv7AoTgwNDo1Nbr1cXJolXFDc9pLx6LcmAKhQL1
I1rdbmQY9zd+mGtGY4e+sejw3qfr7xq+NrO26Fkqzmwe8QtAWFaPvFa6fQLKc4v2
/ZMb1Aw21ubQ2W1LLoJIqsD+eZHbMmnVLzOdsQ/RFTH0RRyBG6otaBW0rUx/KKQM
OlLKqV0H09WN1FrFA0DKGDOa4jKsV3U9/fTH9wQvQqzpXFM8e3le44BAAETvVlUz
7F3FYMDMdtquuaVrMyfzQN82rVujBk3EC/6c7lEkB4Pa5/IcPXPk7RvuIksC9dy/
oALIL48AvSGO1DzQkSCDn6HVnYsKvzPn993xg06U4pFV/LMGbgIy9+JjOuvFRSr7
nSF3BKhnRU4wcj0sadKsqZheybt4LEc3HGLBg7exfgN90O4PefX29f9pf1Uk+VLk
dBsRpMO22GaV0eQFhU5R9pQ+nX0NZlE415IbgeyF9oTnvWORvYm8oTUC/rMuBzQf
DXDR0feGmWB96C8+jVbw+eb+Dvqc/sop1d/FPIWsdJL/0ACofOwCGMNfr2+3Rwba
TjI2t/CYsZBxI77fgmGEw0ZSbDr1VddRooEz2MmbbJWvd+BfJs82MwwMdnP6keiB
E56nRtzjYzoPfZjIPFPLN3CPUmWvftXCm1E72ZrXSNZxi4IH2GActVIAcXaNx+Xp
UxMmADSdwd90gw8DUOY0VbTiVVGE9eI11Hyz0Ae7aHF5BvjeWcDghLWlyt7P+Vwp
ibJWhr9BsM4FxHfdkvhq2FwZRZn4ChM+WpGOV76KywZe2whSol235SLF+8aBlYVk
48z7YFSuRG5e2Rib9yBXVfUi7KRHD/Emn6tI0nIzRur4lSp4XLJkaODF+VrxCo9I
zOFeXuzvSFR6mk5+4JEU7mynkXeympUuugz33ve5Udeh3iNjP9iOpcBT1MFOLPbS
lKE9BkUBSFdlwnfGvvRzeAO3toiPwi4LbySEGeUGvkolUMNc29PLcpQo4c31SFsj
n0mdYC8PBzSsANFcANmOvQlSz5b+Z+1s30J+GDx7NknjN7+/A7fP8zN2h++yNSOU
0nOIYqGHfTKY/8/3xaBIIFgikVoXejQUmEBXR+0sK1O0EWemVNf0wqTTFIr2CeB1
2SCj38S6yabnvD1/D0g0DQUtz2gTbL3e5JyqjXB0n38cOouVcrV+2H/oi9KSWj/A
JYX8pwSbrHIqqMGGKPwNs9suLjrG6wX6W1IBo/o+JLB8xfSWiyEJ0iO2j5qXd1iJ
JqN/5rc+mIlae6XaEaVU1ke40TTCajdoaQoPOpFd0lD5fcTgnyZ53QJBX1ZKWas0
+amRrl7II0mdKTNL/pwLrXHW3x6MynJniLo0ULcAJsIFC6lm37W11gVgQjmB0E1b
V54uVaUsuyuPl7FXb3TsTskm1UX4hcDO5Rf4b2lR2o1a9EJYzqWuDhZGUCJBf2Fm
PmACgWA51GvFk2Lai7gs1njzcQZYFgn+KO3KSa/NSkmHmzJWF9df22kOj0tRfY63
xw6XebSzzPBjrl8VBfGnvpbyj3nz8ZCINdQF0tzgfBsbsg+OYo42f8l1QQSdXW8s
I17oG9v/Yzzn550Tt6tZg3qjorbrgTLAmGKTMvBrtpHaEbYzfvaowYlhgY1LelZt
eyZHMOyZExf8FFXQz02gNNp7XOdxEVmsfKXtxjvHYcAFD48gqntrRcywj0Rnz4p5
eSPmhW5w1RAtdvoy+owueQg/MfaO/vMFTM6a+pAPjgH44JfzzApP0AYBumAJ4sql
SNwsAIfz+R8SKxbx0+wgJPQ+9O3w3SBOWzWaMvU77uWgXtQo9+fYLcgDwl7kRWzb
61Ps+TCKK6TTQuRMmQwlBN3GoYUkkeO7rVrApnOnNobWfymF/gNV0fXS2VijHaOs
FN6op9+gI6HqsVZWrDtAkQqFfnt6umliImWve15xWABo29b50zpGqjvbQkil9TeS
j6POoZyVnodY4t+N3AnYzY/1Ixd3v1id/VD9OPq8VK3ngv2Ai7NTy/Ja9hSd5Fx8
tyKCMLRrgmVBxIjcuimYHDguU9oCV6kt75hi7dKQUWpm12MnaitUTF76B4c4zNQz
1DQpkPhqobweQ4So8w8ClnOdMNH8xh447XsJGrAf/X9Ka6iVc2PEAw8qU5QZe0gp
2FXIT8bizGBgUr5viT8tOCYcU4eR1Jamj8hnfZJMeDpUV8CkaG5h7BQMr4xK+XYG
7tBB0ac3qZ0qeiaCxawUqZYQNFPBDHZGqu8JUzW8N1RozyKfSmsJbB21PLWpRUyL
ALqGx57cCpx2fWqHZP+pRAVkkkYkAMROdueSdAJ1MKOvt1CJkuerrzu0qaX+uV5y
12W4fI9biTeNp298YByc14C6MasciK8jri0o1of9aJKYBSOD1G/Sok1rUAlI6cHA
A0oCzIUkNyC0fGIDM7HuwngBmzWwH/QwRsAKPKbf27umRiMZvIL97hN/jSP4TMp3
/Euuho7iW7r+YIRpWweu4c5qN4GnbQLuN5D5eZEXYPDSLx1DMRDpJcU15l2BT07g
W5tAg6ma52jDtNDV6Sz0QvK1ygy+H0B8UvYZrUmOQ/si93qv9RqZuZmxOfOl8xNp
Cdi8xo9ojiKgo1JF3WtI3+x+Q3+Q9fRPQNLHbPwKnzuGg81CLLcy7CtGauELMs9+
IzWVNQjofjUsv/38jlJp24mNJRPsZPGgBOtJNjABkRuERscAIbnc64jQu5oStlad
+qendo6u24TqWi4QMDnCw0Fnhxmb5RyNi7SVJ7v80I7TUbwuQKR7OjxlVPUwAiM6
VSpW1A9OBLlkx7tG4BbCRRsTM8O4T6M5B5+SWjIunCIVIAm8W0jGxCG4NyXS/CLQ
3b9ZiShG3xC+3894cOk6NQrQ5eeeUHRwiyfH25iLGUSW+ezGCePmOUr/Wiq3sSTb
+/ukrjdTrmsRqB2MysPL/s2aqLUb6zhYOQLRE7BSMyxE4KA+7jNpCOoBP6r11mA4
O3F8oGXYnlSOqRUqvPCH3u1tUknLMoqGNBRlche7Cmz72j6fJP6HNEujDQybH1XA
K+qKjZVWwS+w9jLamHk1eHWjgzrzK+L4Fdc+KzoFSjx4Mo8HoTVBadi2l/UsTfMT
xxQmlxbpB0vJJ3hzNkxJaJEaE29IZJDnbB5iaqEOJ7agBiUYyQvntYOsVm4EK1yp
b+xVACjUmJds9yqXYSkIObS5ApelzEqf+GLRarqjwGDBOO9Bv5Q7kqWxe2l3rZrv
BunoQ5MMKWijSJHYUheTmqrae9K+AkxkZX7E1m8pr2g/tgBxMOXbQWKLiueoKdrK
+hSaPgKqer+DTrGOFGyaSPK6ZKBu1tVFsVlRtRbJi4bX+jLF/1tuzLYJ9zuiVdHr
l+WS5GjSKg39ZNhjqhgbIFbIu1F2vXaTgn6YBVmzTmsJGxrmryy1eaQ5lQQgxzU9
syg0neYBMVuhAuKaNrfj/8SzO5XmggRMfWv1bqcGor4HEfFaVYZ8PS+zZq8e5QLV
d+zv47bCiZi/Wn3GReTb9b9UzT+umLrXNRFYOmsnR6rRUfiKlPM90iBnFMY/ZoTS
o0aTPMIenk2rvMPoIpbOq3HRvjdA8x8s4T3IdnOYaEL6aWhkute/Q3WI3vEHuE12
jreZu4YlzSsxO1vzrOiDe7xGVymTFNPEBFFiAkjG8fYkTzZwXALiLNhdvUm9d4OH
/1LssTh3ktohb/AgkfjQEBQ9ZjaoRW6NIwsPteP/TTMYdGCTZTKMnBlyUH7BpV+o
FbYlDAU9PSrOLvhSmxM6mv3rXIxz+AJkMYlcXzCtYjA10zuat10IvsmGGylJFS0L
vucKhNJFA9tRaQ/LqouOPpYXqLyQTLEdTIlHheDYeWm0FufIju6q9Kdt9nvW1GaX
QzqgEdJoc74y7TZCAF8nN1mW/WsCy32BtAGWUBSCp2hr7yaczqrZdM9mT7Yzl4QO
PK+/vYyZdW1wVze3Obr5bAClg/r5B0QX0yZA3N5L3VxPCaHK1THG43TlusM06IV+
ANeNnUgxy/pe0L7Xcs9n0s+HOYRQwi5oLDid9VWZZJfjrPtXRU47grPRl5ZviI4U
mhE5a+z3qDixReau62peejuZWGk/yyhaClmmY7s50dz2HTd5ai8YltCkBMZV5TXI
7hdbLzsJdMQnN2v7pArFAmbKYNFldxGFEoNpeWa5QlEmpWepHUTgmpndgBTHiO10
hgnIHvYJbaubSHdUKBFn/vcVXKYZ18aJfBX7PjzrXNFDHjkCCAc9HX0oJJFEPBaJ
c/ZDDEy1ZuWWI7QOF8ey+vB/f+eDy15v0iX8PzXsVihUchL9+58Ep4BlSInWwZ3S
I1u37U4yBvTcVm9zVMj3Ttt9+36PlD/9pouqlkKxAzfqmK5Tt0XgcGRUp2K2qnl8
X0d6W93nZvpjb6sA/2US5EjFWubnxT20746bdSBs0MTP3TIV0TRH64XmUExqt14M
uWlfAetQ8xf2YfPS6EIfCkmRZY/xKTjpCzOY0vHnH2qRFWIjxVgsz4VGzZ+govAY
1vF1N3vLpDTgl/3AdTZZzeJsVlCDa+7i0lau9ITDcoSXor/6og/zXpCQT+QclMIA
F4PJov3Dr4Ih5N4o2PBp4IpiWNjrnYVktFthWvs293AP4h1lJyNJmPBmx2DKfpoh
Sk3LRhySkvI4HmZ6LAYHOsrMD4vkCv+emHAashFUlmbYhsAtdyzWYetibJM5Os1X
EEzDt13pJS5VdWdAIcEgcqDUdSlbczCneOumKDQGGVOX1tHVn0cVI3o/omg1dmHP
Xeg4Y/C6uYl6n85IcC4xGSkHjEFUEwzuIB/XCZLkniImg5Dn8G3oYmt8Q0xvryAh
P1kDY+r1p3q+0PMZKpfjzVBfreraYuYyZD6GvgGqSeQuaDv7ukIoC44eNUIM0sPW
2A+LeX+Gr7FLUnCvm+tqj4a09tBq+GDxmzQospNyWKjqoJnvEi1qCbIebrEK7DfD
CSK9j1Kkd5uspixZ1x5f9LcpNlNwM7UQdoQ7hssHse8BtHDVRHdESQRbQsYg9p6k
t33jZ0jvnxontYNDqYT71htKVKYW6XaV10V89AnKmp1jTibGHC8lRUB1dOgqnYjQ
P+KiG3lGnsKr79L3kd3aDwoBIx2vpRvRXXneiZOgIsyETaMRipWMR53nOaqLhQXg
HJedZ2L2rK8QO5s2P4ouMCQzusZD4s9QbbKkm16HHZIm0jochPJebAk5FHFjQM53
fi5d9/OvXUKFtHX8SmPf2Iuc7RwuPRimCz6FZtfTL/jHZops1Uig4xIyb8JfEQET
fVh8fyrgIcqTRj3MHPGp6V5qHu8pqsL48PO3m21ysWWnLB2qNTLWvlSB5KE/t+ao
u3QRu3+r8WfkOvmuuMLxR5+imIISysHPb2Vs632RBwykqIL8qAs9A9sFcrEkA55c
varUUkFRhtkXfiX0xeP3b4FC6sShogu08HcGSdvWWTRRZ6IKwe47tfPICF4sDFPh
7ri6yZM/IYPlRJkg4u/VrtwvT09pA9BOssIrdpIzfUuqmzTwBbaazdLgZ3sqPzqz
nzmb3nOZvm0o5E8vFFZTJZpLGu8izpElnQf1EzJfX/2d+pczI4w2MDSH7MhDUvx4
Gv62tTd6gVneT4cYu6MbywOU8zcdOGhZsBL/jT+iiii10g+o7iXBcmfTPJp5Goh7
SqzYaBWLdTiVv3QO89ef6YbctR5YUXlNPspxuzGdGz+Q28Xcbcvyt1A7i+Pih5Jx
mAUChRgBnZ0C4OhOcqozZ4ZU7FkyQV74C5AyRzKZKjKtQtIToi2Ke/DTVWeWld0h
pf2svGy543N+VxIVDZxZ2cE+CIhsV42z5J8S3YrE9rgKyq0QuNePP4LckD5LjwhS
ELlOQMYnl1BLAodJc4Wt+6to0CSWxSQfdHEWoIJHxn4wR7LfY8oRB4Mh7BhcNIm7
LU6nYI5C0g4e7QAjeKzV3JIe1o9DD/EtX2TiO2uDHBJLrsbTDVHvNNH+KPgYvtXV
oiiQnPe7KgEDYUehjMM2zl8Ni7XDvEE/1o7/A6Oh3GBxCp5ebRperZrs1S0J4Osk
8ZemtiIn3l9faTRlqYYzOuFZN/og7dt3h9zxa1KxEfIgoOT+fGmELyUgzgVJCXjp
Sjy5D+Hy/CVdNcTQqu21EX/gEGg8q5ktx3zu86Z5XJl3PjNPmSNFI6ULokuFthC3
Dzh/isFAF9pjQhD17jGCSa15FGsMNinQHT7Y9LFo2oHpxz0+f6s1PCSntVwQqoZe
9vyp8ltezy8DaBrVW5u1eW/eV3SR29NCs4JESi+TjV1OVlV0l8uZW+IN7Q+driR9
HEPlIAi40zaDY+/y93lOsQOGuG7yLwj9WMyI/t3EdRtEU7uW84uPZRBsOzZY5BJ2
jWpi9XkPP8Jyt7b3STpm3oa+Oc+JdiqJdckoespBz00zEfIR+zm2SXdkxfpRMQ36
SaEWiZ/vgnjeQG1LOv3v9OVtV1gY7NsPE14ncyEsTMnlCaBaCkYf1Nl4y3oT97Ri
9Ov7Yk48EulR0Lsr8xvHSKTX9v09tDkeg9c+k0f4PMtzmI9/Jb7Va9hgi1ZA9QL7
rlolKmX1lb+ylKHKZzFEq1WWiNrSS6IVBA2k3gWcIVVm51timI/dR35eWP3L6chp
2ekbIpRq5Ios5VyPMdB/U+LH49/xSFSvOOc2rGSrChXm1HMa1PpHApxqStW14JfL
tMw8iESbx8xmF4voUrUXiZOaaIuTTS5YU/jOHswQvAl/h9W+vObAKIN2uCZj2GDs
DC1yvkFG0Kwt3jDthqcdgi6/LiUQP2OJk2TfxT3WsNX9sYeqKRnHQ2XraClqcUOY
RkynYXnIpgBSCJsFl/SZbnNJ//jWKs1201tmYjfN+yhYOPw+zlYZLTHt1mqyx0gD
hvrI/KVF+RxWQG0+o+DNuGF6Xtkhz45oCnTroHF5wpFG762qCzd3Wo8y9vC0MgpC
c8JGuABWZ8//alKOa/rNJ6zl3ilGWZQegULKvnlxl6DvteuDnEuSrRy1ixzmLkTN
8Yl5MI1gK3ixHyFwu/uiZywExMHo8aUlObM1Gnhsc0mHxBSoEeOXsLNvJAHxtPEY
7eCiJFfFGnPQTcQ2Ad7iaoQVYzygClETo4iSvuPcpj4pBwFv/NiLX3U6MZCHvicY
c7dAdWE/+e5dyv3CsREW+H9YN2uOgAnNJXePeaC9iutpgKJph8gmTb1xi7NkCX+t
t/oJWgLSGHpOp2MJR3wmMRJ+pdLtC45ki/QuFFkcpU9h22GdZCMwrndr37nl4HVe
2uS8/tpbj8xOJHvkxP1UQzo1+t5oHjZCVQYrAPDopV0sFMjcCpnH0i8nNfszfUWP
I/CDEBVIunn5U0FH3pUB79hL4dA9XRGMLn0wAXTZGI4tx+6X6WeBv6h1XvTFV9sf
yvvY1MxSIIDF7Eivr08Nbf5gijNHpMrQCMcN7OwH4quy2V8Qg6cHX9M23hz5AcPG
f3pKuAK/oEqC1x9DYBRO8UXlUorZBxdQQg9587vqaYNNahZHV4HW2r2Lc8XfhKbc
UDbeRu8r4Nomd0cVyyY1PddPMRCUWF+gQGTT+s6MoTgCW0+bm0C9oYJwoGpgjYAM
I/8nrzbRKAtuZLf/XQsJWWBPMrld/xWiF3p64GMZGpqyajiILGhXd3WhpT+O5rZd
/G+EfrEsyJHyr1GguFo4Wr6Y6FmGqz2dz3/Dmyj4GedMgOm/u8E5JtfNR8kGIX6w
ETL/psWB4x/bCy4WAVyYKkSx9JuMc2S8pTGDRME9s+ejuGo7vBa/t/x+Drlp5TV3
vGJX7mQVeGpwtwZ6d01DW5AvbAHesO/wm6mxM1irtaKdvl8f1vtUe1ZXreyFtH90
drL07pIqCWUSsqHcGCLqgnCw99vkanTLRJSTGekk7M4wLGUqhr+50CI3GWc5Egvx
OHOev1T2AlL2yVSUFmBVrqTz1bOCMtyyjo9valbckpLq0HXMRrenK1tpFgN2YFjJ
rL3kMr0JVKyBUIP+jktx+yES069T4ORx3KJ+WlTlM7weBwwBCfHutGkwpGdLThaC
USNMBSF8hI3SEA/qbGwfi/iFFwkeypcK2zRbWBMpyAKgPLdxBdfzXjocEFKVDJVM
pizUmu4og9zxW5vVeZeW3DSiihfWbsab3E3EKV1tpvYV3HB2IJyPqYGAyVX4regL
3L6RETnGwSIft962dMZF2ygeBEbYcQZ+o7kHA3VqDD0vpNqfjRfRf/cs+rS6JCed
aLbwSNzTEs7m06y1DOGewt3nO8iiYm2ZudNi7fWvpwJMjZQSmXfhBOssNaHyLNU4
LPmJ0v12pEXZVQ5CxYZzWw5VQt7maE/JI6z0BW6Nu7nhIBgVk+URiESEPoRWAQ8u
1xlvLTEZpge753sfhSQ/ZhnSjLGNouIwUyeZgv2j3QvWdoZYjlJoj9sakDGe7NfB
r7qp3aLN5axEeISq4UZ5fpEmXtF/83kgSX0TnzApr1UShadB52YyVe5mfPL4SluS
DhNSNN8Rx7SR/XlYdOGieDvXMNFidMflXmFxf7Waafm/cBEQ//s5J+9lmOggrr9s
IkQI7aPG4Esm0ZiKHS8iZx2zFnwovcbmcIRhzQqwVQOk+e4HpT/a+9hcWQOONWla
BKl2Cd4l7FXh5d9y+wFMTmqSuTiAI9xrIb7011WhuWnLlQd/1FpLCyjJ6ZwAC09O
q6Ro6S6n15nxoKe+V3iRWpMV5yfzoEVJMLp9JsF1BiyLDcFWwWnPKECZqSqnntTi
d0v88vrVbBsjJa5iYe5abPRWY1SwZopIIP78vFe4g7NyUftg9vjBKhxNss3ZBHZ5
sRjL9ACeRdXHjbdOKB3KIPNc6s8JfoaPCuDuTgumzBTFaG5SMQGue/LM+F0JBS3B
MQjFxQxHndNzf5TfkGzOXsPcZBf/gSfyhXOScZYQ3Xm2Jg2M5JzmKEJmPG6qoZWp
CqzSRsuWhv6Mk9EpSG0fS47sQIlECtKqHOO6wu/ZsxGDbQ7W7I6pv5GfGjD2gmHp
uhMYpfgF2abXh1pIUNkBdFjru5eZ0ijXd0RSZQuZmmOcB2rkF5zAsC9qIvtb/GtP
R3gSroO7zDrpvSY2x3fAykoYdfj2kJAlfT08/LYjcSu3uA+O+YR2qtJfz1Yj9yBe
dvmQcR2rrYdpiQUEGX+XdjALfVYLcKUnlD4vUCvX5besVbqaAUhCcnCHIFEovMEH
CEQdfeGvsnQd0/9s9ZOnPDwifxJWfT6KjQpHWFtyp54GuN9MnUA8yyEPI14BZyPQ
Hbac9n55gbCu6APLWBMV0U4OicoXCezjpCDf8vk51PT1/Za8Zu7YwZ1GE5KOhUMz
WE8De4nHyyzyy7w2hsn3cTRXZqOJ3M05brD/yfzoJXDzIYFPz2xh1E+9Xk9okC97
3eDRm4+j57CHeyefoiRS+AABYqb+7W7Mg4MlrR98W9p20XGimuIIsWRS5QL40EmC
8V41bcKaDzvsjf0WqqpKuUupK1VORrrzNjMReeqjl62X2pS5SGUc7lJFcuAJCKvS
hlHeZDLF7yUDY0G/OVNAIhhLNhAQgAxRo2JsBl5o4P5ZcxeshO5E6hy0ReLWi12Z
ObT+B5ZGbprxKUWukwHLJufiXGWc/lOCZCghLwXuRoLHBQkwuumrdwSUZI6r53Yx
Ab/WUqYr0mRpoK8GoZJZb78qGC2TZgUO45QKzOeNUB2kk3WGcp7WZvK/QfrAZdO7
emRtcpnbncpGkdMLWxh8XZmhQQ/4ejVXoFUJwmeW4Z6ioD5li0UwRXUl07uLfMIu
Lz3At1tz6ub+NH5G2Xyp9i+btuVaS3aZO+BDf0XMXrIBWD/P6HqiAyVPmAjglwRG
itHWukQZ9kVzNZI7tmMuymkqGcpZud8XqnCvu+9vU0b/948UWXU0Rg9TXrLeT7Da
f+cwZKsv49yy0eKetWG9I7XRaYZqKIdiS7jV2mroU/xSpdL0OUQKA1D24aohLjJg
YSyrNf5j4ngXO4AiKKDNhgp0aNd+U26bqD2Fzp01GSuGPoq1jZVfUGu09Fw9GbuX
w5PUycsEVaDN3MgC8odJs7I6OovPS0Ia0UJn90J5ukWQvjej3ZQZ3aH8GPCyB/Wg
+19Bawof39VhsoI1FQJzqZ/ZrSPQpv/L+Ch+1Yknr2Lyx8CZRFeikbsnvxh3YQEf
QadnWEBudIUqrREGV83YBsWn5akjJfXbfRDfWGm3J7DRyv2vpEO8vsJl5Glutkab
ui7ejWZh4iPEI1bpfXOB9V0h9CN0hb9PVxO2KuTYR4FVE718rdo4L1Vik15k2NNH
o8f16YlNx4heqDVj3UDTW7IcSRYr6yb4Y4Zt4rhnM1TmEc+/5ib47UQl1i1tBeeS
Hb5p3XNWIothGNvGu/N9Vf1SxXDDmjZInxeqhb2hX4x4n76esVdSBJ3ybwyrvO64
fjCErLUVdA9QiGQYrJbH4cluLq2R1hU/fN/owYCvke77aAI8wgZx2bgaEoQ2MhAA
4Yq5ZpIQhRg0NQGkcRKkFq7hbbT0UITTELSiKoL5OPuFyPeGomCZwQhuX6sLlNFf
q703qoZQUhD+b+iwVTGGMY9VKCkyjqMPsSq5RQcRqCAX4sI24tCRjFYjfejsvG/W
8EHtmvBCcOfNbWuqq9fAccG9w/Q5M9Ow9ZwbjHIKDfqBAj2Zq1s7p9jyCSXG/OLl
kvMgYL+tyPfQ4SVxLuvlDnMUnEYpY/cyja0xTTEmWeqbvWvl7q3bB3b77CWFGb0W
WVy861gChP0jE4vxHibyW3XbqrnvZ4HPXFHxprejG5L+WE+Xp6HeDnoqe7/IEbqY
zW0Ss9VFEfi2SBv5CPoEzEoIk1xTB4pWzW/tjVTeofsubRUFTJzRLwKGjj1gdGso
mXIzu0v/4QtLJddXKfY8q7PWOfylJbt/OGsbGq/2Dg9NqqEBzKAdaDr0mIzikts1
ylYgI4pYkv7+acN5glTSyOk/umLLybTcGPOX94j4jvfK53eZoack/YYgoyRIGLhs
5gtkr2rZ1SHSOs4k9V2Jo920h31VJllEkcjXuUbVa44LtNiYyM0Xs06N54681vaP
bQUralBfoJg8laVGn3hiHHc7GOQzYgCWb/DA/6fDQcI91Qqu7NMlSR3IoB98UFmD
TDSIvDKQm+cwufTx2AH0w/3/4iAykqHsqs+Q67MSsenHsQgxuAEaLC6LdxjacbDC
HnkYSWghnGYSvjg72BPaN14JMjPzr8drKX7F/uIX6gzEgGIHf1pIhXidqOP+h/Nm
xsXe9HyCkzDrP2Ji3oZRqbmdDq0sLd1VEvhUFsd9sbyM7xbegs1tRfBfEDlo9vr4
oAWgdSv1UPiE8o4sC5OzIdBpReIeV7KGwW77AIgkR51VOjX/ly1hkb+DNtIAfc0P
yYh+lUqdTAU1gQOdC8koCeCxjRWJmyQPQrac3unmMKxd442xBZKHxwkk56P9ULGB
8b8noQRBvZZfFxLO1HupQtsxrrZZfZ/I6m/Wm8+VGcIpaVH0nIm9OPnI5dorAngX
0j4n2qavIE+sH8M4Ju6cQ3H9gDEkmcpk9O17xXpY/CGEqtTYiHSPEVB/2f5b6fi1
Jyn5S8w8EQhLENpNh+EpB4mx1wgdtrB+RFdXWx21Mrpozo56KdGwgRk5KecLy4yg
oksWdA3YT20It4QH/MNHp6hUmf7Glmq44RTL+CK4YZS1eNqo9VZp583n4QJAPCOF
YesimLq83BjuRkJp8K6ea/zitMSVkKDoQ+BnMTc9C4bW7aePP0/OBVYwjOTRX9SR
B71YOFAGFyPudMoHGKL4cjzuPhe7oxcLGsCfQ+JfLO+HhoLBEsxBo0xaRgAYJ1i4
T827sj2e4UxRFFLI85oKuW5VZVGPyYT6x7SH2EXODNA6wRvs8Js5N7NaH7yBNRPc
nD+DNoi1bTigy0MEBZnH0R3L2PoB3jxjVonh2aJ8dHJJ+lkJ+MJMvuW4iHk7l8Qn
Y/iKRjgoIphaxGrqpLvIrWd2ZX9dJvnrA7qAlXagoO0ROah/8r32Pynwf/uD6Ug0
si/MmuA0UsBJ5dW6gIZeQtDh2UFSlHJSkYJBKvNsBFo9t6laR0ooeFL9f/W/uZmN
vgCQI5X4G7z2hGT21PGU2QTSVmfh37WQUQKrBCQDRZPwnM2z9LBRD9QX6igADEin
xqKuTm4NwZwAOdY3sfnEiBzFDLvNUStwiPjoYfSp7+nyuzWla9DjAUjNQMV6VrkC
YE9wU4+Po0L2hI5Y9AK3xxYDitsc0t775KFx4HWef99JL1kDPgB1wTT/VzPpMUbY
eFrrmt0NNZX1v0wF1JPV4hUohQlA70EvsYah5wgiPLdYWS8U13zfdiNBe74J/pLN
vjqtT84WvbFdcnMMlN4utj1gaBHN2UPpvWbVf2HXVTP81JqtxIQJJUsv5BWf3ZYq
wdGql1b78fthw1aZe+2cnY+1Yr+UpmCoolWPiV/dCwDVJeHJlNPNBP5UUI1iZCb/
iJsLURJ2W3el0FnWOLb8X6z+AVBRG6ecM0EgJkAJ9CG+/Q3goOG7u4Svs8pyzsh8
N90C11qh9AAxWfnBlM7WrUa8kkaIOrxj01QkytfzLtQis8snBLt1g9lkfSTQDg3l
UrZBO9+UQyskMewt2P7OdtDWwJJvwXFBAJOO1UH7O93xXzPQYBm+yHMBScyUNKfk
oas6QnPJI7lZfftJQhjmqkU5udWHJ8vbTP8zIKf5HT6gHB6W5zky4se/W9+LkwpN
OlPj6hGp3KRZb8PeMmdLiozQpvrVDCMKmeFtlkV4ITyWJOxceu0wp4p88lGMLIjN
8BTjIrl56a6uGafJ+fzwKB4w05IPT0PDkK2Oyq1Z5SZBmvfpOBgoCsat04KM7tIf
j6qJWD2yjpAOgcJMh/ZKnXOX7nlPofrVLx4IlViqNoqGSwzacLp8q/V1s6YvZknq
eWEzdHOodsdXRleeJDaWCFrSK3rMkxg+TQc3nex1bjH24Kc5aEbX9j2AyyrF2qRm
1kh/agyHHoDfZ4m7M+d71KpvpIW2WaQRrDJQa1aPTCrJaHtxTM6uIjLRB4jSYy3T
uYr2R/VPoOdwJ7BD+isxHs7A0uC+++mn5kXAZKk5/M8YaqMkIC1s/NRmls+hFiLG
uVu1Z4cbDNRLoCBk4Dzfpc5MURpZFtO1hqDs8FA3Pp84Lm27wFn/x3jOF3uXSgKe
zvi2qBNzno2NIrnZwBpX0YuzpmOMUqiSXW4w1yRrICsUsba1U/+6NY9TlPYM9dpZ
h6AdWQj+hei4gHp/MHlWahvmzW2vLSd0HXXjiAcPB8gRYsoNV8Ut9cnWJL/kd3q6
ZOPOAS54I4xMGM89ydD/qpEn31Qp5zMa+H28WQwPuxfNoWXQyVL5Ca5kr5oW/sJh
ZCiwVOob8HFVnSCTjWQHhLhuIkzxlkYynpIdG+vj0OJ9meM6IJrndIJ2dufkN9go
IH8fGEGVDNIDxIglbWu/HrwJhY73QQiF9416yLLNF5KM/RwItwYmfWzRe8u2KP3g
rhTsUK/wTGqKbOK3y4rKclXQtz9uGEdXXpf0tlIBBFkrXZEkl5J6Vwdpz+/hu0TY
3EX8/Zqt14NYPIyq1NFtUGILePWFysOArA7Entc6sIJms8ax5HrFh5lN0CguFWjW
r5b5bc99Qv5CLRLf6AH2RZ9bVBluTI9nQdt6LTDudJGFo0X9qonUfrWwlLHQJA7F
FpS3Z61L+5fCKkQ+lAN1V/nKjgSYmiGAHIquiu5VVtC/IjS/xDx2CEv0FAe7sKtS
fk0+ZrRT1zuYZxWpESp8L7XCSJcAuR3bxqr3VtN0D5vqkBToGsVGiI3Pix2qp4uc
FaqirbitqNgUXkjDyKxq7R0jyX7wWq4Qn3SKo0D32VcBeekClktKP8ZtTl/S0NN+
ejm67QGLFF7a8OwktsHmj+ROjJY6d2fYrU51XLW78surREZsEPc74M9sTgiHqSmG
ZQn9AbX5Myyh8LuPbITjLInY7EKEOtg7kTYbmXavk2mh99LiHI3MpjYkJmwXfRse
ilT8I2ZIgICdSSCB0NV+o6rMWGAx/EoMovqHOtTJgPcoDddcOFf65TLC1ah0/aBB
2ourFIhdr1czseRr7CAoUWkHUhbjne6xCr8vMLHUlFYtWiGcU/4evylB69uyLlXP
SNrINX5dH9qq/CIa+4gqHtw4CCtoStKmw4FQKx34U7pUze7EEafTPtfMK7YqedUi
gmZCOqxS2IMQlrK2ntvssam75yUfXe+5XrbmKyu31BqI+6i8mZPJ+sO9xWeHmsp/
WHTBa9gd1suyP3w8SCPNk7ar2k+y5UeUI12ftlthOSFkQNXIDGX2X4NKJN0Rrm4s
mDgxv3rv9Cm5V5ITUGjIjTj4we712aibueyyq9Wy72DBlslgO2VMQOg5k5HBs5CN
OYRux1fmFo7WUFfkts7NVAJRI2TIkgKp+cRqPJFu+Auvkb3EOoa+X86LAl7MpXNg
/13xqda2D7tLz9DgoxA0Vd3lqxxphk66BCidV7yXEA166YWsrsMxyJg+ZUPJ7Z6L
Epv/4p3ZN04QQloOccsYYR8zwTycyvlKszAZ0oLcw63cxoN1h09bZGVDn4CgRZLF
7hxGGt81xCc9GqgECZg1nPpphYvB1o63VQHHHjwzc2QL0HFJMSQj7RbHQJ+7CPVm
Ykx2KKl9S2XgNyuOnenIPbTCFrYUwYHllKNz4d950D9zL2MSGbuArfDVYzut55rz
Y/yXIR4/H5JVWjTbnfAy4kuAmMTaLGA1XjjNS7lkuOn/BTkPcP5kFZqcr/pld8pk
A1vBuO7Q/yS2RRcSKaewVXRfNKJt28T1cdGvnoQGhpginwk1/MOIf4byKeQe19eC
DFP6plRukZNX6v34epXLsBmhRO952dEStse4fO9XyDZ+75iGPOHDhuQDv20SlL/Q
JBUYNRG24L1IaUJdtdce2Cq9cu00YqK3pT09l93Ka/Dw6J+ASEOUeg3TYr3OQHLO
ReFePBRfd2RXK5OIpWcg1FYd8V+61qhWNbn7PEphOvsSPofpvjMyRctwj5VxGh0p
sk1+zqPQAyjUMHPCV+Qb9l+4c1OsGcrE/8EIu1UEZPv+GWVJ5ArIe2MT6vWipg19
ojla6HnYA3+jZ/+J8NmnBoy6PgL1tORkmD7MptN2UXAIU7AneIZ2kO3JhojDeM3B
1irOPkClPhQ+0BCuzYDOZOwhod0TBhL2CMFXibQb0cHt025t8Hq2fBp3Q559hhxL
tVKb12F14xkt5Jc+YMgSEpf92lIlnMRl8Ywe38aVL66f/Jvy9wmvcoPAZaWTGVLt
jwbalmstCuPseTvENXP6Grq+JgCKc37sUCujgC/OmU8cHMG5fg4IpcGbVuX1Fuv+
UDOQjDbQc9E7wXpU9bLOf/i3MCwoBJTT16BF3dQESgDVlmFbyrG+pDSPEoifYN/H
nY0XAVxraGiUdCmTDYNz6S0p/3VJ00rhUkrneM/KH7GU7KedGkcpLUpUoxqqts27
XuYputCEamLTyN7sxsZMrGf+NlfWofp0xyvbNY4GVqMunlNc5945bTo4APNFJYcE
s6TqHYZPu1prWI+1N7X62EVCdZ5vKMN4sTOyiAcHEDKAL5vJO4gAZWnBBDeOxpH0
sv6yExpHpDJ/V0rPg3d6CJOVXX2LQypXHbJMdbFZ1B+XKXRuacJSyvyecjraOhbg
ALbacVZ2x3FgNZLyuokB4Rkq68KbnLElf8HSHwjZdGfOog5L3zJca4uc02YwNpo5
N3rLqF81Ft6KqQSz20BHx0xYVvgcB9qwcdPhzIVsJEvxfvh9aV+qA5SVPGanSwP/
AujLWehJ5hbX/aZp4EjCpuwDTCMb9mZV9shTZYt91WZOvwluqOVzPkbN7/I+MqLn
N8Mu7nJnGZedAlFImEQ7lXF3MwGqYoR3BlZKOXatR9D+74AnEIm4DleCCrmTWIJe
1pgeHvHv68YDCNXpfKpmFRbobX0EtH8azYuDMRutA0CNDiSCGgoa3CUhW7L7/Iwl
ycLTkT8zYqzN+BdhggUbUXjYv9JEsAsr4bP98mBZ0Yzyd6a1bCs5JIvWDRc27Qhs
+P2Y/OT66zU5mEsRRf7WBCAhoZEOO+kFeaQGX/tXa3W0/uhydQkbWXJ+M9zve12M
PTlq4LT3WWMy7YZBbrEnC6lx97qxicV2wUxYiUiV0ULSpzU/pGT7T6I4CKGxGG/1
ej7VlJQSCB2z0O9BabMHMN54Ey5116AVvIK2biGpzfd/zZXmUcZ0UO9NCmK2s49T
fghmQrY97BqbszoTVqZSeRqiIFiB5SO6kv4FIS6fXizlP6NICMh+JZRw67QIa2sc
c17g885MRO8Ne3PuQWBCPtZt3QNXe2/NPPlyFIoHqN2fBrSNHBPFL8WrCakEphrq
ofGKbvfTp5K+JSKS/brjicdKctM2NIEqEnsXNlIFgaGY7q5VVUlVwxjE9b5B/JZy
q4rDO+oCS06QG04u2PSG8tE5NHKbVbCysaYDoiObYCO1h3b81zSvMgQXSMctSvfB
UB4+p9+4TmSS7TrfZSgOQeqicSBbP6ZsYn1uOPkHqX35GL+JcH5mYNc8+P992ZAE
BIpUptao0CnQKycTvW2Tw+RmRcIV8SWgRtExcKxgssePd8UJP/y639+EoI3BlFk+
gj3zBUu7uotVhddEUBplhHVDDlNZmc1b09TqgObB/Umnon4tXWAzqXas1TD4bY5p
f6srl4mBIFAmS3tbKipQffJGuKJSkf8minrNg3l9+cyDAHOvHBdam5o7DFS+9WfN
L48ljuqE2qIMCH8FPCv7HEA1gZcoQWDRB8XZcZEotaK8CiKyIilcOrMlRhli5Vwe
hTi/aD34OR9oGPktOsS//6Uvjru60cYfGT44hU5d5N0AylDtyv1eexRdnHOaXB1B
4U6yNSK0LdkYuvGhdDPcP4ukGFWmz6b2qRaOA/ynodfAqrAAT8hKZk6deh5oRCuV
7ZhihLMVLavBBLk7DnsMDAn4zCbAviY5jrfn100zOFEXryCMWZQrv6e1qpr4GiJ2
6eZY9RnMQ2GBvT6YR+7AC79KB+TK2v/4ld8kLIIZXI0tssKCRgx4AHij+W93Tgny
8+M2I06QubZr8Dtqv5MyJls7h9/OIPg42a0eU3QHZzeJx+OaulpyeTY5RotntK8y
RGYGRuzbnjK9Z8SbdEyTh8rH4AyQ8Lktt0gOetoasEo1wAxQZSxyf/RoTK6vDjlS
P+94aqGmpwOYhWj9cO3UExDH0IT/2hM7TOk/UCEU+7rzqWGN7Y/8WuYtYGKa3RWp
toG2+hWfB1Hse8lxA2VO9/puwdhxtI8DkymoUIzea1HSe0IPdZB3NSJs78WsmKOG
lqbOu2eNCqQOnPblM/TWPLYU4n5eU8ToW6lXiK2LgS6mV48nEEpX00RwQaeeWSn0
8L20q9pf6hZRhnGDLYI/wSZftBks1WJVXM1LChOoo+DGU2BruoDXJR6SZWUPFM6U
melLto22x3PbsjULUOO9AXO0cuUjF8Oena5UaLMGJ5EwyCquUG0Gc/H8ILkcwF28
+atfygrf0T4bjwV20HKKQu2HaenlsovB6j019Iz9j7Z4IKPXw18JHMiVY8AW0j6H
wBewQQbFbmpu82atr7N9rTVuHkS0ggNh6nyq0WgjxZcMLBktuOfUX+3PTS5gpe+l
44AxOYFbOMgj3BcoWPvhtSSjH2BRCI02GG7w3bnh97LpAXDmNC/YTJyzSFVjSRP4
+2pW/MvnZJzRtgO5I6uwTUR2Q2qGgLvb3qdSsm2AA/Xq4BBsChoaySnTX8Qi9yt/
ChC+fxhXexjlznwm0G+QhGm1JBi7pxXKbc7xg6hombPwbRAPeLfTp+8xfhQxTiKY
VvT5vOJ8DJBgjvIR1zqRYxMIGp7NUP1TF4shtlE5A8zqRsf/QY8d61LGXnWvhWdE
ZjPWgCsBAu8TZBLCqxO++W7gFgYFtcAFkPJFa//QqsQzFeXRnfsV2btBC56hgT6h
Jx5uYt3Bod0vwuE/Zwj9mSYCTH19cZ8MSaGfzi7HCKtaVDFNG3l68tLDO5y4iL8F
Rt016wVr2laEVchFFpY2/DkOLv4MacGhC841ri3Z0jR+Jmt41Tt9z0gHRTmR0bEy
gNjRPsSXrR9mHN1+F4PuKE5KhDkjYMEEI7w5CD2S+iKG1cL4/5mnlRtQaHn/X5f8
+sTgjokxQzlHVeUUy2FJ5yMtEfkZw+KW4FQm5qt3dzVkdCsnCL+GSfpmJ+DXoXeI
EWlJh41cfvf5E+Ta04g62rLa3G3dye6VA7Pks5Y+BLnB3nTthfXO+XA8u54otRRs
kSNcEdJFegN2B8xtqAJIRj6yKcGVeDX2f4vF96k783J6VyEBh8BCm8x95/FDxnN1
ixOpWMF/tcWBON16OIul2SFgIy2P7gZklk30uHsHqy/E5duh+NqyJdfDdnJR31By
Is3yHJnq+WhP7Tsnty6Boka2l975rzsn3wdrUbtLGCQsqzUiXR1k3yWqvb5sWASU
sxh0hEGZrryRGNIZiORCOsPxW5vyxLkOjFXUburJdatfvQEYNcn6gQ9PmyPdoTHz
3jvgZHtFLYx+SB/+AwvqIb52GfHugTOmBQM8+TsXJ3VYRaU8oalivgl50Cx/J716
qHWqLjXQFMv29ETAK1IBOP5o/Lv6/3Z5kYhdbWqpAchKZ0He4ETPdCGbNvBLwpag
AZLJKkdGJGuXGOeZM5OtOlAp/cseFmPoIuYxQ3kMgBpVpVZ0AZDK5w7jTB1YxfVI
YAbmsc7zmpv996Lm9eB0Uq+ytGrjbkLBF/q6KMDapeiSqf6FOCNLS3MgvG8xC1Ml
oiB0hAwuYj1fWP/D2xAcpp3Ja44gFsa7JkoRRTJ4Uw+IKSD+5ojN293LHIWHUB4e
u15UvG1q+Ag5HzocluMukeGbWkCzKULIXYZ6opxK4qM5nOnxEG7QJK5iP0+rCrAG
snKFdt31kEK4PMIxWg3syqenvpMLhN/pO32MpPCHxf3rR81uRo7GH/8HG45CyzB8
7l2zsJ0lgzrGimGdjGNPLwn81v8NrVlhMoQP37n3IO1I7J6dmAc3rXv0ao/fGBCS
xrRIciI0tNtOWoISHf5ZadKHPCt55xZEMKTRnHYOvsau3c5Q8r2m3+WQj+3NHJD1
Ecvi+ny9DYoFeOaFBJZ8b4CsVtogjrXvbqvXNf5Zw9cQ3QfZsc+C0aqJxC7YNDrR
sRL79xeffupjmdtZvOraTvNAGMsJd9NAYrcou3G+UOV/f0YM6yhiZjhre0FM8Pc7
cm60QEP6yWbjrM9L5ppyx6W/L9TPD/1tjUyX9ddFzP3TQAJK+p6RdsCDfcmKsNJT
o7YL4Kls0QXs1lNtEDXiZfY0007saDjl+pbAai9XkjT6DOfG1wsmzn3IkFCreLnX
LogpMg7rxjm10EaMYwvVc3Kvhm47uXxLLQRGoOiQtdeSeVkEvhXybs2U9E49foLo
1W5w9mpCpm98IX0+6E75F8+PVDEIwMKXTTEQyjAdql8ZpDAxJV5kFbphqdSmw1+h
puHfrgUvAJO5pQa5XYpD74KxXVLv2TZJjSQgqMDn/nbCb6eciKaBtdkqlYiRQqxF
UUwrVu7LfkYYMrWdHJ6oIgFAr69ISsII1jcvNsoPm4V1NyWgfXPz0dpYPHKPQQ+f
uOAeuHZXkEbxAIdTxXMgRxwCWsfHReOQXtKWY49olAvFDNNv2uV9d54d2gukKY7H
buzlYsNPkLKlNuRkvhvlmwTh/bIqr+2hyr4UNlQwV/0B0LISlRPUYOJ/lCdh5pE2
z3qh+2zaQhtsoMLQ6ddLcOZdP2X6LFTWcULW/mGSNngLkBnU21+lt3yq/tYc41LQ
5vJMIECY7lM20Yz0Xyp6pvcPIAWWrXf2Xr+GTTu82QAgpvGBehvjc2ja/aLme+G9
8yNa/3LHk2LIuiqrgFBeC9SfcDGBuY8ol0SZ+KwkpNywiBZrsfbukdgIfEAgdfCu
WQvQZn2axycq6OTr1MK6ggMfnwN7hwUhuZw+Gcrk9KlCFFhqAVmygRyl488+u+Ov
0xyGBzl1KjiA0gqZFLN8dCrXAs9tGmhOt77CXcVA5p5sfa+BC+Lv2GjdPO3Ji0MT
okrr1OexYf+pi7jQfMnpfmECgP1GTUkKYSPUFxtfMg383/B6FPQ2ZFqcsrDcq2wi
e76sqPp3KqHCoLLeGixK8nWRYbu7FrMXK2pxtPnQ84X8T6ryRRrMfE6aC9qEIJVY
ksvSfDfi6k3sBDBzWqSmxrXtmrI6B4DsZC4o46n5jFucAg0CRwgk+nud0BKK2RCq
ucmLlIYjCOTwOlICBy0t3XiTyi38BYKBMC/fbxYYvIzMaRf34l5GWH6b00iPhN14
juNZ1B/4BcNnegg9mfGDMr29xvl2OFRxDohTos63mL+17k5kShDZYSZOvdg4OF9i
93RcM/JuakTMbRM0SgcXeufNL2qv5PR+2GLqDlyO3Jqvoc/PieoM1gUFBrkftPKb
KFyLLFH/dC86oUT+gg4vZWaChCkTvfuQ848EboKwD6ABoouQj9m/EbOvaJtTYrNR
lXMbsU3/GYDdfSPraTrb1WyNyN089JFdxRaaWgnTSsMbx5/XMRjViZ8rpRYEct1v
cnET2ALTFa3MKfrRDj0dGVgstTodmcoQTt06C8U5GA+J2B2LjonX4atvU8MsJ0fq
KFwx53nSJTx9A+q0XCfeYcmpyYceTf52kWyODtER7kKroQ7YMbPGuc7QcdH7aFjs
j6Bljo8snuXCZKWPDZWeod00ZwCEpn9/L7OUnlTgFEsPTM2y3xD98SjXFS8bEMj7
ovEbeJdEhyPAgz7xC53sbEQCAfbE/wntpXDC3y95R4qqXEiZZV8v0CTN8KBMYJmr
5KZd1RHrvmG5EyT6iIDT3bkCd2mSQiK8czLQQ1LUpqDBQIfUoZcGx1YvLz3yoI/c
trzxmNLwlx/02f9vbIk2gGoUHF70YfEGi7KTH1OeAY5bl/OaYh4B47gu8Db57Nzp
mlaTw7deXK5giEe+yHbpXb8Gr3PiYVTeX1YolKHLRIhbhEPVUX4HDdSDSSUPDQcC
YrxDvDA8onoilD2HhUe6tue4CQ8QyJ8icga2PESe1F6qn1I6KpjDLpeEr/jR1KER
IcOQblMkRVLndt+XazOJL6bFIxX4qMXTuzP9+he3AbfOEze6+ZvDdoqUk1TjVwYW
S6BIRwevAXUHGt5YxEfwBI4Vx8CeHlTh8/HyZt1vKnsS8xk8Hs58x9NcGnxrYUZr
T8cBMIpwFyy2WCEWEc7SstVBmo41QWnMcsSP6S1wsZ7d+Bk5EBLoeHD9KtP2Hnq0
ki9Fuud6VPKfiiaQ16kZXoI8TLXGPxqTZpLIRCYff9d/iLjtjQ0amv1IoIkM83r8
NfFQcafRSfYOpi3wmeAFYZGrbiBV6FfJyNCmEUkZdbUplvu9jLh7dm75L4aYGTfM
eIZbEVY2x3eDfsvR/OYZh5fIFffhB0AcppIZ+gD8/fkH/dlTDUFCIS5lrIiTOD4f
6Ixs8mD/aW2m54H1mtZGRoauQErcW2xwpKIkF6E9rUDsxpz3mGp7FbA97LdgMvg0
gBjRSyN5WCzlwrBXus2mI5fGyUXdhw30KEhmWBQqbmnpkdNLglhsK2C0cDMUE4FT
equuIlFqIeStl7mV54KfVdYoYclip6aMXMAhnqnA87qN2cSvfuOj2OPLLW7y4A1P
2qTdhAbLPdH2q/Dddg9lTSiJPl2iOHsc0Bx1MuA8ppn+IqzwqnPCUNHvySG0uT+X
tYAUeHYbL9ABZI6f/e1QbYNS75+HhD1yZx8vimprYGR4dAhp6eObN422pX0ZFqOg
e0hPSnX1QHN9CsDRM7NM+M5WIAjnPbtI0pPoBM8EQDlMQJwQ0QVF74DZeRt/m7nj
Ep3Dpod3Iicx81HY/hJEqJzGb65AIXhqPOcz+zyl4j+2BWBKk8wpmSZt4ugQ1pyU
iYK7E1rBrzmi7U79h6MvIIayZgqxbvGOU9z2gW0Kq2oZrRe7CpPfJ+YVV4Lg/wYa
AlmfXCAukH+Fp0sdiexPADLNkDQSd/2IaUQOBXzx7bfR5LQEZ15ka1hMnfa8EWJi
34W4QDxJ/rRxAz3jIgrQX1RnD3CokfP3V3U5xN1ckAwFkLAVDX4TzTSsEMUWfyn9
JVKauiBV3x1KLSA8mRrGPOmKAmsdOCtbFkgJ9Ue0xjuhOtEpuWWNUHebVts+2Hzl
ovryARFjWbvaKiPgdBNisHfMJPU073KnG8HUaAKfkhwglMDMo1ExK5C+xVCBA5ne
Uhg0USjyd8z0jidxbcyA7pngi/NsOcrspO1W35Bm+8KrI5F11qqAI0jtKU1SvukY
LVuvHAobLYkIe3XfDb1UHcdmcN6qf9RoIZmI5+b0bC++vcPJbSCnSMcEqAvV2nLs
8Pd/dBEAohzguT+00Bqgs6RYrkT3zpjqV/rHPPZzDLlz6dEOeZo7RMQT2IytMBLg
4xu0IOWcDhvtTiFr0LubcDsOMSXHKky4TXsO11VUH8Yib9hgRixSAWWkDE1JKmE1
yjqk+8IAtZYiDfjgpbeUNXCnhS+LLALl786cSoQ750gTqe+AN0iwDLk0QqCEieOe
AztV3aqhzQCJiBRwQaJYhEleT2M5tlF6F48kBXC81tg4U+ofgnLQjfz2j9Jneqz7
/Ma/rV4y4AZ3xy/S7gEtYDm4lj3vf4v+unrfo1gSKjynf+5bTSaV2aiMqTBE2h4S
Pw2U0DQirXPjP+9VIoYZ3u8udX6v89fTCAJloXAv27aK/S/3nes2BU62euj1UNgN
0DY0OGFFx0AXt/XNM12OdFrJuh2DcilBX29YoP6qMBzAxgDiRkaciYpNfX1hAdc8
u3+3tV0tuhl+sAFpS7fG0vdlQFRIUrO0BiWpqwzsqjIJatAZH9Us58mcS2xQCEDe
OPohJMeZw0tCA0O4xRmKALHlPR4Rfb4Hzk2X6iP+EGY+dtxgxCXUarDGwOom2OJy
stQxuVQZ4njBvgTUQxXhFmZwb9heebRv0VQekZE59xTcpOuQ1KHA7f9RGfepyI+Z
DV6NN6abxo2leNlZ5btuW5KQIwc3IGoo+sdclbJOPSviOZrSnMy3XRt2NhEtjuyg
A9tljw3YQaurJI7ewcpOuh/YXJuD7iumZiQnmspyE5NW/uMhJ3eI+f6Ki8dtClKQ
iVXyq3fTXmsx79V4AkEJ76kcbux58U2muxATwvxou0wWZGni6+mAoqwrF+ssDQFb
S8ApkSKHpvwQCup3iXvGi2TIwmDQ86WfZvnZOiFhOdqP0YXnmpovu6UzcEXc5SZA
r4oMCCKpgY1bchW+J/IgvsgjD8UBegw4N78WdpWJ7Q4volzCMc77ERSEh9fUYJtq
vQ9JV5/k6qafdXgUSYl0z2u0GTau11Ymdj9MFIzzsvGYP3zuiuGIGZTcrlLu6VN/
oPR+HPv7HdqnfcI4gNWHu09LzX7hUy/vNZMU5UIUGTdtcY/+eB0NuKmNC0DuYVW5
aB8usYkQJF+wfUxs8y2eQTbbnkWQ2tfqYrIrDRLfTwD88889dGsFuEgB2AZM8/VQ
aJ7YT02t2+x/6RNYUmQtJNGB88erLnDGnXpD2KN2yDzTRbo1zTxB4m2JVpCERTLY
hEY4e8/Y8hIzzVJsGgAy7SPqzMb08LTG1bZTizv7c7iG/kmULJ4EVf/75wN9UnHB
zWKSXo1Us7ryhQ2VdD9+Dg8S56+TNBMaxc7FkjV2xnMTzTCS2nLdkI47xHXugF2o
cB23J7FWqipsmA3bNDbpVbzj5Y0SpNiNo0J2cVLNJIwfFv9o7fMkjeFFJMbL6sfI
jD6p5RiTdQp9T07Ob4WXJn+26sdxkbi/w+b7vvs75LE9p98Ton7vErYIGoqrVE05
HrWFynmtxmZyoL9UMZve7rlKbjj1UD1i8bGtjXEew0Ld7m0+k+AVptFwSi3Kv3fP
B+X0a5SfpWSYmWMxJO2FcutxgyYS+VImcihO8wMbrDYdBePWOPZkNLO1pb8GqjXG
VoGJ0t+wJj2ACpuMdsyLP12SibZJ2ZxpwynKu4el7RMyefn/WPmrn7DmjhOSXucl
d5q4xiZMygcDkIGgQAZSD3I7nwf2KRuIxn+L3rUYc6gpOoPuktuKnH8mENZq7WIU
fB12ALvA3T2zzjGo48e3hZpSmP4K9H3m7ruCpcoUIszazu4qBl2nG5p6TFS5tVqm
w5rGuvM02aYXV0XsVuJgaTLq3K72i7CHQocoftaHCzPntdpbUHZlCB7OtT/VZoCB
6wDZK21ktMX7fWrCsgr719egKxxJWBWsHzPavsyQSBsnQ6H3gj5yb07TP8Spvt8r
DlhRq8kznR/BQU1hseSUwK39FzRcE+ouc9QeEYhWyzvHZwpNEh+bf8iJ6rr5DCxk
z6cUYYA6TruTXltgwQFhnTqqW/NJGNWneYQB+b/W4I9nCmq4Ze1rpF7lQt0MijUx
7mu/NG9/t6L+tWN9AHxR761k8/Yzcd/bhzpjI1VY6PmZbVBKcWHayilVFdLJwYZy
Tz0mMgdi9r9pa8AiiLTxyUJEQU/gvqyJYpchnpbjyzwBvZ4pFc9DcNHhrM55P5WI
dNi1jT4O/Naph9BwMk8KbabhLAgi3i0RLsPNGA+d6dZRhGn9+JdDFbWB7ZVi71UT
B6jf0BolUm9QVwEkjTXJt3BiBLUkHhLkBw2SKs8Gi0c7w88lcEgUmNhIGbOkqrCL
IMPozEO6HNnzXKRIDHQtqHaLC4LysoNLNBiiMYKfBvL54JYGqH/qiQnYwlcGUTbn
Eez1/FWoEzykMhS01Mk2cFZ4HwYoCoC24TEdgBsyTZW+EbDP21kItByxC+1SdL3e
fdyC79jZeABfoIHJnIKX5y6MQ1LNySZPtpSnPhlAf3tGqGj7w2XO16vx98bnawiU
911pBw/J8mBqtKYwnNeCbV17I7xVMSzl7rUDIpsLvS5Iaqp6np62Zu6O7gONywxc
Z+JRJRZ//9ayFtZorUmvFAXWOLmdIExo8DHf3huByedbhzf+ETco3Wt8cxB3ln70
zMxzEkHFZff/r8aB4cIU9q7ovv5BfeaPgmFmiFq77M4f3v+jCQCunnUg0ApQe1ZU
HqFUvrGssmb7BDRg5w4l7UajU2iV861BEDce1UHzOcrQPQ4JFnBqeNc3bKiGNLb4
Hnpz9a/20xFpNZzAEDRGznITswuQXH9rICCJ+P4h36FAAtCYOL4+r6gqCLRHciTo
ahcNyOFMk0IJzRBIit/xbeCCn/mybxi5mF/GVmbFfBx1Aw2YLuG8wC5b+yyGfTin
Br2e14kC6rDRQOkqFohKRWwOT7bkrjv2Ef6W5PJLwUobQJZapy7+hTS51seVJvxj
zoRPRSZOQpAYQsMgAhKTCBglpwbSSmQuPeZg5+xqwx4ICmOu0Qq6ut8odxRTap9y
fDwa52yvy2J6xdhT8OEKOpykyJYawVXc6dJ63FTLo8d7xgJD/3L0Slu+TeRXLdAY
p7g5VBDVrBUs7UlVx0WGVov04NcTzAFJwVtZg1mKmf/8ZBMf6Ed6ssyWnSUhBjGF
4LJ25fjgelu5XFCzqp+NNq5O5Od/N9LN+1JWjSB0NPdjEXCFZqAD8C87YmlpzJIA
6GVQmHDjD7iewDUOCB6ZT01IFd1FRRI8GPmZE8OPZaMNIt6nDzZdBtBl/xnFAh9d
k9FbQmehgT0Dd84KmQMH2WlYWo34+zvT2Yy8q3AOo8K31B7wZL2rVh1S5mu4dQIo
qlMVnPKkiAas5gt4pLd8h+j+33tWZP6Q54q6j7y40Ii9+qdXp9eDWzKwAd/kGfGm
QW6czFFJb4swRI2MGqoHvPuVDNPhVKVhH5FlMHGMANZpx9fn9jVrhLbUfl8w4JZI
L0qlCvymjYgwfbEbgXPeiuOWqHIaWvbXDGtJCA6HzWS4QDi+3ActUVNwRsnrbl8J
u8XvDAFevKEZF/ZP65pemZ1tqdON70E/RHmjtdw8wyIzPjtS5PAwTVS/QzAKYLM1
BC+glGudmA4z0PgZBGLUtAC/xsLG0tFuz8ksT/nRqFMUA4smXYqRUovYh0S8DNcC
FJyeixwUv7Z8v3lBSLlt+33ROIoNuBK/eFLMIGKq2ee5v+W4KuVeDveGvzOGdztf
3xaLWBwjCUip8c1LBmxBE25sX9JtqYrq5BdqIvlmuBwFNputiUVBBKsFPYjsqLBN
7wxGww6Eq+IBZORjLj/fOrgdOKDFyvP1TFdaRtQxJZIqyP8AI+J8+faQ1KFguxhI
o8gX7txYAQHU+KRbYtRpS6gN7Hz/bmXASe3LgbGqimPWvMWkH7SPRVUcZxVxnFSr
3zOJLcngYgbYAsaHlA1eTBaTJhzpp79099JFTVw0BGoS3kgvQxkVeR9Kqt1JULRa
HenXOMRWdnnm+lPdBXctY9kNzj3SrQFzYdR7jMrXP+hTyjfyLC92ewh6NFRv4MYW
OjMy4GM+KHktK7M/fLSANhTm8/iCJv7wNc53sBY+xr6A2VxeidOL4gL3O2XTKrZ8
uJRQV5din94q5Ctm/jMPTh2EZzyUYcm1DxL9+AeUymfZksI2fzZIMEtUFDNL+7ik
+qbOkqPdWzH2jkRFNRTeev5Uh+gCD0Zp50OcYr0n0RI3VAnfzQDdDlFVBhBoMrRT
o9Xqlj24ZfsdQpHTqiabOhZUOc02DoqoXlVXROpl4ldaZNYGvaV+Ez9LYyPKiRMf
LnfaHlVcJ1HB0nDl7M1SxHyIstWQx8VRZGhhhan/wOL3IUhj6C6z/7FB/QR7k+Fp
FjeiF8nYpYU2S0pALLCoxgtOTyxjVUC53ZIsJlpvD5HAOdeV9UZ2sbL2BHBMetcN
A8x+8vLBGhlngk4MPwwYgpHPrPF/fvOqXB64ai7FBw//4BDmKuqIKB++E0NaaMuY
tpVf5XsZ6m+ekBK7tAHWMkzPKSK5biYM86M+klIXoTUch64iaqJaYtk96ardCugj
rHcsWNl1ZNwpM9vuSTRw2YvOXPAHy5j/A7D9jojQcJemdXUMfyyCo83wk/WVieDn
3qplm3NWecmzE1v1KNB5BPXrZZ89qxptT+0O0h11Kpd78gqm+KRjg9ThDDFNlan7
ezlKNLEWBNfAil1yqptixPog6y3I8wOCQ/8UMM6KxqnaZTXIGNHHKP0Ox+UzCMqP
hReAnuTCFzqDKa1i+WbuRSLUBW38qR8hXZqfno7mCBzbGByptwhksnE+Y5Bb/spY
1XZkf/HEHNREccxOihMgb6FqVtpq34MUWZJtRnjTmM/Qu8bcBG64g29FG/m8QxuD
+mLtRRmMBpOIiBj4kMrj6y+R7pp9HO/u+Z7NEafXrTQ4GAxiNHHkL6ydR7J2Pyf2
rNmHzlxYNnqnGLUEA0UANWI1lU7R3OuD8btxa+YYwaMErIKK6lTguDptGOVPsqd+
WFPCnuOVf1EU+FQoY7UWTgWFcoHQ9gr9AaWtC4spAWzcZJM7GsxP8X94Elr0DR2z
e/j+Sr9ew9FjF3mQrjtU5o2uPOlSY3BV4d9xJYfpV29K26PCV5UkvgNmlCPi6ojn
QL53ZAiXgNfXjlmXX6axLLL/J8GzEHM7Uek8f73HkW3JP5U+IeV7FKBM6N/G90Qe
0FuRjLVtH2o7NQ1vEzKSpAaGu5qN4/y77NcRIw7ZO+HHlOyD/cKeC3Y1jGGDDhug
YsVbN0T98yv+KpgwijOFDZPoD+M0/EoUIPGuv2Js69cknFydog97AYKfx4u3+2m8
byWUb0A7OoNl/hiqN7fIvTMbyQ8lT1MlLO2K4AVtNsm7WRnUZaPrhmV1uDUbSE60
mTuK9zTOwp0fLT54efANAsMSQ+deORCazq1dBe06/RGRjDDnS0S54b4OSR26dQ7E
Ha4S+CZJdmCDXsv/nvF/9+v0dN5pePeHkyWEmLoYNK83sGmnQd4XHIzouT5rkv9G
sbDQoiZf5qkjhX0wgocze2sHS999HqCSuEqP3h3JLhF/O5ZEwyI7C9JwO+IKJG2Q
8pq0bZF0HtuCs0pZdPQNPjl22XXXeIyIsMIlBTrIAFfqc83JRYKRHKJAvaVWdVhY
XooCzWHUdAFpbQOhJ3IqcK7PimDA8vT/yvKxVT5HkepMsWAlthj8GPi7sbmlSxTT
aCggr2rS+Pc2mmMRBnSxEpE96cSdduA+h3xDNlKgC7gnLpn95mL1NL7bab6OFAbR
Gw6K+uQftTxGWdd1DqFSFXQU9U0/3nXErRBdx9xgiygno/u/MHAR8H1v+lIp7t2o
Q5wd88t+2IhuIW13Vzg9Xia3opsNX3dC8UrQxNolBSyAAzwSTWjoPVf0m33clsVI
94irHP1EGzu5wleHE+P6q74YCA9ByEGD3QPXBaYJONSyZm1nbTd9thh0Du+4zRdA
OZxft0pXoDgh3JCWt+5pyzXCip5pJvCEP5xXtEgxz2JHQSdg0gwK/ijxl77wfZMs
LflT9qFpeIBkhSIduiBLdS9dR4EoqjhAFVVEQNM4tT6T6gM950DZAsTicMaLdvLl
02pahhecbPipsAkhRlA/ajSMjGOHYuEb9zpJcAA4cxJ+w+5l7a/r24oKqdqWF1mP
DNEkdM82b/cMVU2Pm40ImZRMVK8KZ7ZmvjCTFdMCZsAbNzhdUUAPV+rEazQmxRBQ
paRV43k0nOicbBskz7iLST+cVMdX9agyHu8H39AahSpjwr3K//CecF3sdOC1A4Mk
auvnVS1HPLHDlFPQ7ho2bdNfueq+VD92bYbFkkfi8aRkt9MVXdM5/fyi1kelaT9T
Yd2DjTnGjqebeBwi9iwyyccQxqskgUzB1dE25rlTBl9uvju9w+pSHMmy0xLsI+/l
oBV5WqDZqpISR5mtU8RcWnUBqx0VIU/oo76opi2z39Or4YUXwS2gxUAWwjgZEzAy
eVcXD1fqfGb+rzqOEkrQbsFcgGpib0ExpeL0/1gabD2kUvPMVRQqw1a1p3UNDYoL
acDb5KHBrmwCLegMZfyXWIMeHXLnLPShF8g9npJD+DoUPb57WPoioVESgdVjdPmU
0BFhIuBHpHXTA+/q0Y4uZ5anKUVuaBgapmByS84G+qBZUuLsjluAGytBihC+XFLc
n2ae53yEw4SHCwV/QZZeGjnw4cyeeO8ZBCqzZ6tgau8TaYUfkzO95T9TvZqsJL0s
AaRw/c9O8r5TIaW5AASXms1h577GkKofzjWWvifF77nfRc28aq8pcmIoOnJDfntj
jt71xkwY6QXabslJOcXs1n+EkorOQTPCmDNR2Q7+2+q0D1LJEyhrNCQPuR3lYjBT
yl56lSfV+xfZmR9842Mfsq7bipRCCNEL/Nq51035/dWjBcyscfuiiIpXYW4wr9vu
F+2UQ+2/dGwazoUJpgu51tmjoVsAcfzYmoDTy+vOh3vdP/vYUenU+adzSEaBKUj1
eya+AYy/lAgaEMC0uHykLLh/FatVdF2z0cvr+8lpeZXAeuWeL36M1PSY6LWnVPnw
TAESVFTH0aI673n8F8nnrIJXwvu1/jHbC1VjOQ/otvtKrznNuEtTNSoyYQlsBq9Z
CQvy9yMGNnc9gYnsS+vHtvaWiAXgfchAuGqbpu28gBEjAiTnhD3jgw9R1JL/3KTi
4bIMPwuoOUfQ/P2eA4x4GFqIUBEtekXfgMJlmb6GP2bhtH2DQFoGVCBFeOWimsAz
695sbX1rPAOTNcIWVtGvToUk51I9rJ8ydJgrJ2UhJHEYTTfb5YSXTlJ8fytQTBCx
khbtrKaHhiSpjwimNPxyHBuQFq1hxK0WNQ8n+Lm02hVrYQ3audM8lj/Q/8JIdd/v
59rLaif5e1Q8WQHdYpExmNI4RPHUnokSpD7dnCrNULVBBx631A3OlvZSD3WM0g4e
K8TZjpqIDIvPaMoiJRUuu1fd96Kbyk6yoTtXJxH5wmVGJcI8y04/M5xLvoZ5YFva
Gr8m6QWDmUsyKFI/gWIxOWQy0V1rtFWAEuxjwBKIDEEKo8uZPMF3uWJsUTtFo6Zk
mc/eTDBnBdkGjWgA1Mrl/IL9eLEj/uNM7J1MAw63cP4v081OnxITfSsUZl8Kt/P2
yWvnnKeZ88VGvZBGwGkL5tTv6uInwg6JcE42lBvRs5MJnyY1Ihe94zeGu74XlcQG
b396W5FA8oVFXbqaZiYIcHKulSg/HT8R7GZpsLy+m+wfy+HRL41X9Z63u5zFeKbB
RTOAOl7nQHNdru0CUHLKCA0i4aHz++JKKxcvXTyhUg1mVQkfk4m4nejB2XqjVYas
9e8Bevufur5xSOsKgrBtIpqkeFfTmbeiJClCzOtRMfgmbxskGG0RDuN8BNlRFxIn
bvctw2o2DZlXiJkGtdHBM4xybo+IIuWZ1kgkl3yr/gUrmjQ0p5bx/OZx9SiSQNME
OhoyNmgEMKtH0RlU9o4622lCFHI5ZQrGjbpU76y5TggNiKceHOA4LMEMGty1hlwb
zidEXFRivlX57U2MA59HD1GUyYc/3MEJWnLgky4DT7pvSr2y4Ou77yOU0/8q+5If
lxcjliFGrXeCN1+oMRvLz7Q4q/wJLoOtkKhbSX0Q4jYtTf2apSVUBQ+BlxCwPqOz
jGaqv8MI6CRtk9tmMRmPbLPbZauP8ttMxb5pJk07yBQ1x3y7I3IhP5S35ZqC/A7p
9nn39m7DIYSROi61oKfgBpiuIt97QccGEgxK1JHovwBn+vHPKegXE9dHrKKYPCII
uts2TK+S+JX6gh/eknjn8rhxcK9W/uoADZ88D+Lsp3ZqyTkybnV8HTqWEreA9dKA
7TuyGKgNWw7VlzebTMN1+gGHY8KM2VEPE909PBiGwwQEVnqaO6XYRTuyrfcz5YGC
AUTdN4cH97M9bc2X7KmluVacUudIiw9hlbuKonNh4Z8KFGFdZY9tc3UEyfV/svcR
s2zZ6XsgjpO8nyct62zZBfXR7qRksHyHApT0iD1mOeMUBqBO3Z3R2Z09vqe4bs1K
tQTBIvJp/hDr3FZ017jqdLsN796lQGnXao2NouRm5xgDAQ/ZztPKgpw8yo6h7yJg
Y6hrmTo1hIGW/D47o8gfggx5QFCpv96FiFdlP0ZMQYYo0cPPBUizcXyouW48RoZN
y1zIuXyWe/xpCVE8Q96y97N0xQ1kXF2hfTCnJH8PlH6zX1X2yc7P1Zu3g+oespxc
put9b2TOJkAYNsFUdyM2rsqcaIvHmI1g6RL0nT5q9fAoKzcTvhhIgHhq7agtv8Ch
Lu83fg18pqQPY2QH35bafa8HW5d1cYNGGsNT7Jd9nV2remqTssoXA3Co2i6gAbF3
nApfurRr0L4+o7z8Qk17hcHpF3nfCmZtDiwyWCSm7tzpkeeBdZdozuZPBSwsB60H
GNGxsqHUf0+ln/cnbFMXN4p3YHwkGUIN5hDQapBsSYNebaepHLazhWA1IzaYtzT+
lk5hEkqaW8MFsEewZ9htOz+oulD3vcfrIzrJOyOU09BWpsys72BBF86/iydgmwUu
ezlFYCohj4h2GE/QUoCaOb4+nHzpDPAfU3gmnojOq+9CMw7RCVespFuthd2byIYX
fVP0sc63BcQuqWmJYpgRqUbZwS/AI77FqCsnCXCDG/uZzcmUAFV4IxLTv2ZkH6wk
SigSeaOUafSCu+W1z/VF5z/l31S/3AfU7EaAmj37upoXxSToBD9AkowsAL+bdj4J
XrrFWlcmDJijWQwBAEWTLR6egkmmYR350Njirc6TGLRnVVB2tbss3LW6XdhAyVBf
760nrCKxGkQKWKRucXyzSP8c3/N43L69BouJT4sohMuZ3MpXY60s1Cph9ALTkvCO
vUuYKC2Np7qx2e/XQuDxKULmdGDzoq1WE+ZZ+J6U6gnsyxpia7Xa8wfjTRoMAxpY
Be4UiSWQqjnd81mH6HckpSOtmhD+yOVrLMpBUAQlm1c9y5im6FtkauSwj5lN7hYZ
Jo3lf/BNRDzbzGh9mM1ALMN43nylVwSUqZ7zgtKNKZIe92b4soQA49evgBcOdxf0
WO1VODcowV0PDfy99RtZLdq9v4jTk0ZbqbXST3V2df1beuBvM9ryOehkSeJ1WpFy
zXf6pqQkcGGOrkiV/u6CVOTTbT61iQHstPOL/yLTdluy++IhIZaNqNQQpK7nGFJf
p0pqjDmUc9YtCjPDnAqcpvF+x1Oq0bnJvT35K5s2+DQ+BY9qC9QnogRHTc/PBdkC
Nup4nfM5gq91qBcbrARxX1qNEw4VavFlZRzai8r4qyGXWtqBsl7Qh2mdl+HmJv1k
H4sB0k/Crh6yQdS26effQUjLGqTkBxxejon5PSrx+eOu5PufgQr6eJkp6HUgVsd5
TJTaV4SYTQH80JY/oOHqVwMfElHowVSVsIlKIZmWqPMURfd+8idFg8LQiLaeMr6k
kESwUGn0WTz4O/guFfez9kjqKpqT0IEcAFL3R8TSjkyWRXjBok6S5y6k6h9wwGlu
l3ig4cXteaTlpr30rxMsfRXmdDT5TvnhlCEIeFeQJ2HisM8VSsCepaQR6ZBDPDPs
DSLmRSW4fMu8LfKwesb6IULWoZC6xPRqLElQRj7W8gnq6BP52+JqDzhZ46IShjAv
iHpbVmQjXknrY6uPAQca8aCphIG/7yzLAkt8Ub9TkythAEhCgBM78oWWyLy0h+Xf
1143mZXav/ETe4O8CZ7vPAKZ5+vx8VNpxATdB/PNNgfmd3hyqFDdyoTxs9Fwmagh
XYHFperPoBFFBX9NHAYDNf4eiP4H147UpiVSYsnVqkG6Qnx1jdS+LSFHi7iQ2GA3
Vv2O50426Zei9ibBi+E54hta6Xo9vPfdx59n9BZAXlt9yA2ePShsMC5uDPWvQ2hf
pIeY8slsgPROskhiE9oA+qOXOtgvT8ASieFSzyMPv63XSCiSCDHuP68k9MrKQIvJ
xWJegec5W7RCUDfJzOC1bHNAUbbr/ZzJZU8D1xx0CwXY3l+ckS4HH64QCP1CWxHp
6Fb2/xvfGBXP8nxjBjm9/KZECbNswwn15bSQNSfmNgcP5HcMAJoKfkPXI+UzyCOG
kLOCW+OkcJ5XUfAYF5Ui816GFnCZLFisdw2vqQLWZ7PCwf20sPEqjixXqvI4TIWQ
N5e8Ye0azSC0RC9ie943694+q3m0tBqKWinzXJE1zQEbyhubo4wpYlkrMDDkieO8
qAgUFlZpPNR3VR/iXtavdALntQM6t+VIN46oFTwpzqAxhCVfNpOvzFSRlHtq8A6T
n2JO2JWa4T/JsyQaRReo3duRB5TpsoRla+94lS5ME/ouByoA9WINHmiGGDzJPZDL
U2cDMHBeUcoCwzTC4gq6hhU7V9mxjf8/oYidqALHOsCW5ppOz+uIHU9i11lglqZU
F3D6+qkZOBABw9nRBmz+D9cA/sCjB7pu7w+aNp9zR3Um9+dUXIKXtAGt2oCdUUAt
x5npQuywDMivy24W2BECCC4tXKF78FDnEwBx+pbiF3PrdWF3SUcBsJVP248Zi/8u
DPMkuGqVlanlyOKDzGQ9Bm37XpD35OlixPGUfJMczzlvcCc8M9S8zKOWkG7BuIYC
jwyZLmt/E1ePo5307pgYG5SpPDoao+yoAvOiokpcs5j3IlOSBSqmhHK07dZlF+i+
yYvHfwCbY7seGptawPpokazYDxNJzgD/8Jopc50TnAXn9MKz/gvANux0xU9nNbxw
E2tZPpmXRgK5Pw4332xywolHPgpUiYSfPO4oDlU0po1d8r0RcolSMryxPBOKDUOj
tp4/Rf4ZlC9VL8A8ltCZSBiPRRnFtFA+K2KAhle6NC82+ePULK5ocDHy54wTBZIG
+jIZvvdObqEFgmB4eJpCCZtlwFQC+LVcRDD1Cje9gvKB+MbSj6e3IDuSgOkszGfF
bVy6VocJdI8tzOfSFlDvzKn3Xjhc8Ved9tLlvVOKQVxYWUEar4TLWmbQgKs5DK3b
ElE70Ur8Dce/f4uqL7KsnBUbEqAstwwuCt+FkRH+uw6kGGvSQnI4Wy2g6Qt4qS3P
evKdv5IhTEtNApQEsfMjvYAjCV5ktVHdyJ5Sds3T6Zs23PY5SAU/zfiZcKdqNuK0
JUj7T3UdTU7t0WxQdmH3nWb7n6tRPjd9WAkFH1WbYaD/RzHJlNpn8iGxNaFBr464
qMQxWgZCdxg05MrIfv86LTa3a7+qWmQJ4zI2qoFJEWFj/b3S4IjPBW2wjjB65vdE
G6dd8IGTdZzsNITVinusoJUabAZCqwXn8xQbUNz5aCJhNA50IhUsjD8hShfiE9tF
xfovUkwjv8mj0wnSC1QJbLlRd93RyWOJRnzf/Rxmh6nbO6ZQdK3atfgvl4HSXVhG
nkpAc9b1ph301zj/l7hvVt3Q3J74Y9rhJs7VY2WBzDnxhhVgFRDpWc5lhBm3yxw7
0mNMdlNeJvtVLohlPTV1Z9bNJA/Vth4o5x22snggEfBNi+sadyhq5UzkvAwrkPXq
0srLGw5WLusr8q2X1qLG+X8FYcj9vWdHtSWtPYty3VtjCD8bUHWqFg0W/2GOW/ca
7Hl0LzI37x0p6XIGK4f3laWkkPVNQ6z+LUANtDLZ63Pm7AG++OiQna6QXTgPBZGg
4KeamB1baM3K4Mwo6Q5nUhYuD1eUeflM3qgfCYF/r8JiGxEAQ5+qrXHtT/Z2upXs
AW74JnMOZmq7iSaEIVp+q7CzKMrXQ+r1XJPxc2ScK8Y8W8Dy9+gF7mXltpAE21tc
Dm+NjqfsunHyGm7ob06DEgs5qMj9yFxg/34l/1p61MIvO9rZYK9fEIXbHM/Cgap0
1c+OD3wfupZoM2qW4SinFLQpUg1Y5Rz6Y5ggDT48Gcg2B6zjaPyhGjeyqjh7Ugw8
XlxBAS85tOLwbxS40gq6RJaVTUQMwSkHknx/ZMz7KzbQxxnWiDOQ6mcOdp9OIs01
aJqc2i4mAC7Ixd8+OaNeYk35Pc8hP45d64ksvRGzrAX8d7rQkpfIa8j6QIETx8Jr
8PbY6lfZr28LGWrpg7wqwuMSswG8KC+3m4JB+ZnSDsdKrRLvidlfFeBd+oDcDwu7
fWNeRwPFbc6csuewKcripkP8di9eSazR+VHvafZ3UAHQjwv+1kI6sYQBrJnnBacF
Cyerryl7iZOfDq2v51l4ggH4XLurMoTFfRJ4B6maRRFIlCnYqn5N5lSCSjzQiiaB
bUV5oupZNinm99M3eclWMaAc5o+3XHWQSKa9C9QlDwD+P8HVRBgTs3M27//qMWgE
0GVYZvDmbecO4oOfhQok5Xm8kZ4P8wdyGZtlZSVT2cxwfCypFaLN4oTKQbR1Pt8F
pHq4MC24XxJsE6LrLgyqZzqbkGqG5+gFBPmg/85U9hQRHpeWB6UT1C0g5nuY7pWA
P894vQPy8ubGlb0y5kM3tkNEpyZE2YqXCLyzdisQT1qCTbj7Pj6zH+DG5MMC6bp5
TXk8Ug6/2j5yL5l7zhZc9WJTRUOK8ATn7wIFK65vesJzmE2MjkWxl+UwjqDg6eCg
68AztfhuhTJoDkURDrYFX3Ts5xQlZZO6+t5s4Y3plVr0dew6Sx/phkTzPkPoEPIB
J51g2xcHySKGND5fKiiFE3qMiPA7pItWKuW2vPngoSu5B4Yk45pz2Jgyypr+GH91
Y4FzfrjDvDaCWxN/dsqutLQxhoA8QKAi2lj0L1y2ecOx3X5ZUfhxcu9ynPf5pzU7
CruB27Qf08jJu32SOnk2ttMFPld6iOo/+7gdtQNwR0004LAkZ07xjPeyJIcyHf/L
G0VH26HKsTxpgQRy1+SRO6AOWZfgJqaMtQ6ukJsmEODE1hIW7OCCBJKsS213JtjS
5qbnImwTnRdGemQa7WLBcj7Uf0mY/f26Nu9yAzMfetTow6Ye5rPvfYvbqJxoWI+Y
N6BumbP8hgF4rxE41UlR9IwtvLmSRH3mdsx4fcF8GRVUiCRfn81csOGLb1RXaZCu
gltZ7J1wp3KGDAClspnffb7+AWlNUSY5VZ4dawAnddvcser+YozzeG33htuNpw4Y
5bKXvnlwpkUovFKPrLdS/i5R7O+zbYeJ7CyFsQKZ4ZMIJ0hwTpdIJqYQ0+JVMas3
3m7uIFgBX4wHcZ62Xzo9oJyMwY12VnRwme5WCDYosp63rnQeqzhNzhH1BWV08Dn3
njprQmzr/mSaXtxZpOZNv+k3NxLqRJVnif3WMNETPwHKVa7cPJLZqSSlWnmV8CA4
fW4M3VNEBt7EjA2Z7DGXAoPrSoXq805O6XyMxrAfOrXz5VV38l/ydsyawNghhurV
DjP33ZYmyxCfJ/lmRp9zjyx0mZDKeXJ3zUbGjlB/siRwWNxkYvtluajD6BY+F3DY
j+wkPhHM9gFxk8QVFSkRHFIu/P5sZk4tMutPirE4gIUKgzgNTnmMsK3Is+U0y4ar
6iISjj6xbvnQYma63vypsEexIejsvJjAQ+ED45rpuvdfPmSGDDB0c4W85q/X2jx5
TUp7DFdO3IfGpRiuFd2d2buBzmr7aepnSn84KEOEHUyDQy7mA+b/Vn98ZiHVMU9T
YM+Oh2tJL3tFDTJpKZKb++6xqYW+LWq/G+h4jG9McnQs9m+JzB9tjZ5mijqHWKgX
yfK7zjdeH8BiEQjwnTvSSU7tuGmFDyulqz7SDztbcC5m5SbaAE95K+Udw/SqIBlM
JzLvsfQ3JKou8XwRvrtyhDumqPwM3eZpOiRq5ljRSiaW2wtzzbfUDlCu33Zh5Dy3
eqtwQNAtcVnMa0vyRL6qfbMmQN6BJN8WfG/uudR5jvT6RXLYLuWrro7ogz08xtMv
tgxSEH2/XypTNdMMuv1EcMTb5Hm/X4fFoeVVRQy8xEV9VxkEgWcnGow2CGJFC4pX
/OnIl8OCPMypKwlb7j/T/lnIc4wCJ9niRosB95SbMJpT3PqreJaVZbsaepnDMfcx
T1w8/dAj9OsmqbFjeROlSooChxOySSKv865wFQyeXWso6sWbmv5ZQEStY4RheSl6
HCil/Sg5hGXJhWLWH5K2s+FZe5v3xHEoKOSTT1znJC09mSE28I1M7j2WJOaNVObj
e7aTjt9zo3oSt4hQsC021WiymGQHI4ZId6sMypMAhpKzI+fdIwbo48kFWb/ajD4C
vYUuMPeWogE11v+dy0/UQmWarEBTPH6dpzTgQjMnp/jU+YXhjFvB18ft/WQYEyfU
9vzUsqWTpzRWDX8fSAnfpk8sp2W1ZY0FICWjjMLi6DlXCVbBJVFfdbcdOey/RsCV
c6+zLhXKYcCt4hmBFyw8zJxI8FfRqX00+l2REKN5YWF68xJPuM1JWuNkl6RhvA4K
hzgs2mm2ZBkiWH8aTErtXDkUHMX6wCK/Sp9OQrcHWdswR1qpzWzwN8vp3k3HlVh3
2M/wJ39ss/l8ZuBEbrrcyjCrUGqHn7wxHmYTzuiw4eYauH/duYi1sZOH5xX8kB3T
vhPXsLzS9XmsmKPo//BmvIreTYZ3lbIgm4sUn+2tlA/3WL8utGor2emgh8Lc7b23
oA76jwQOEsmUJ3xVFg+lvrFBSqqQEg3r0g92HAJ+WT9XNVlZEdCbbT+W1zq56kec
k6q+CXtkgzW2PABrfvQjlFqiwkBKTcRop0mE/A/BLJvnFL+xd73Ke/ftpDnhJx2H
/9pipZSxcKzgB9puRnsNtBid7O57SSpUf7/YkIfX5vSS7Ax+kh2NVw9Xks5+gKHE
352ugLmezZH2RFTntbMDuq6vN9iBlKnyXwqU6kz/TFGTClfA3Oz2QNSEPrfwjNPS
dY5FmHu7eX/h5bs09WQ2r6n3cOVKkgcJ/pYgtOLmogQov1AO21oDJMAXng3QphoW
/X+essRR8vRQqXPO6nCAGLgFLtA6wL7+a0nDu1r1bPmiBW0jezcS8kGr9IGta0st
zicUOmkZ4+aZQp1FmIxX16PinybKtQ7bGGRL8dKuES49ccSMj6VRLFpIC+7pmR+k
mlpO3miyqp2D/9qjOGOxFa/Y452iJ3X95lWyJAjpnvF80DzT+VmxMAKqgpsKG2b2
sMQWv1DSVP8yIQa2MltCJnyz1HQKZCHxCOI6FyyLwrWynKRBfi0QTEcHlLxEsFV5
9bDtfXU4NPBFRfmyaezK1kB1exxNZ89gbSlDeneUjRUuM9GrHnZpOV6fhW6fPPmV
TukiVaPmIIsqWZaIjfZb2C/gb9MjQpAM9b3sFtPLguKYsKzA4YtsGajIRmb+BL9C
QPT2Mjy7F5a90JaNT++WH183GqRBmSstTyIzEuc1XuADFPRRlsO2zybK+x88T72a
EkdglrhENVIEht1Py+IxoRVGt6hjNSkX7WvRwXHwr2p2ZT2Qnj6XqFo7FAzJeiyQ
8RL+908V+XR5TbeCjYN0nSrCwlRZ1ZjxiolhNu/uU/xsxqgnI2McW6KFphbK7xSO
3ohjxsXgFHmaIflLIj/pyAU94cW3eJdMs9q7lNqFgm1AaD0WKKsujG2cnw5AniBg
2uOYTFeeDw0NYaWsmUEtIOnei3KnHTWfpGx1vEzLdjpVEeFjH/F6p3P9GQRMp1Jd
3PlINqWBqYqVTcXW3tsaPs2Vu8cBBhpxFnVCcdu9ESxkp4rXAiLO4bYu9KYdOeUb
4La7aQINvsFf00HJ9zjQs9m0iyE3tvozeB9J67Wvqnbcce2FWhmcTt0TdHIdqoHK
9urBQmaSNcJOPB+1O5SEdByd4bVU4GXn5AQdh2pmcrbW6cIh7IjXt7jQ4tc0ZLaH
7S7vZIIoXBuRt6B/aclqzPdlxs53gIQncMEXjUJX7b2aVPeRPhzd2GGsMe+RmZVa
pkD2w1esAU4TbljaRJMok5/onh7+IihHdHYk69kQhCWV8boVfYexHn0fSx3GKayZ
9Cm67x5V/yQLbymSTfC7reYeXP6+O25lJoM9GQmJNQdNXWEZf6we+flOlxfYVoTt
MWrjp4u8yjogcTWIxpMAXDzxmHwcqoo2l9jyH9dvAdyr+LvACADDKQN5H2WPj68M
FOrHOqYWUJM9Yjq95vD7lQkfvrbJXScDCbEFceIegiriwCI+AlLaCCm8OFPbF/Ug
OBLqQDAbfCvIcb7arTd25iclNT4sutp6oZ7Zhz3M6JQOvlE3DyX4pV4l1tJWy3GP
MValeZL5QfHHErKUWscE9fNoc6PvDMB6Z2fzkOxQlyVsos40LdjTtetdhnkF5xXD
cZvBepOJxRmeL8O7o+lOcfQLSwWeUUfZNN91c1HWxJQWxeTloNXJXVr0iJjY8Pl2
ViJBj5tmYNYas8/YdFSsJOGzNoetVJANTbGNBPebI9Z8D1CIGbw2xvIMAI2m5Jla
bE7L353d2BT3TZx/YG78FxKRKBIVKnfGSuPl757Z4fauj815ipFnhMDNY0nTTJ9g
sgrfIsQa3Rnj5VNebNKufrFN1aDJsl2IRTacVn62LReSWsQBnBh8WJCXc3qvcin9
/un8OmJ9+u3aiU+s2wXF+MBR6EEMlhKlBgwdxt3ChVs67KquQnTfbzb/KBP/GcGZ
6nxqFvUTQwm7dG0c5vhYQpiiUOgVGmIlUcHTp2yFTiSIzpEepLidqdjRT9CzPAZK
wyNIHZK6LDLAdMwz6ddBUFL2xYOBdC8XSGL9I3R6cItCjHYrwwhkSLd1LvAV2qqZ
O+YBMJfNpXSQDNa2asgtlHaFQ2i4VPLv9auhp2LWBlXq/4DNm5qz8A8L2F3uSKOt
RbHnz86su1RzNC0oepCqCVed+6IBJo9MmOVft4LSSZgLRsIFpUr/8j+sHZwDnaQx
Syiaue2f7tZ3TQBs67tYkNld66U6NwVCMAKrDiUiu9oK8Wll/HdcM18OlM1+iytW
0+BGoSaQzCCSZUBBezfA6Vswf/Vu6xVI7I83xMws8SzM8cmc2OWXBVqW2RFJdUe1
IV7n1lgXeWw5cZcs7pb8IBVwHQRnZALVBdQ3Pbq6013FFnz4HcPfFm67U/foEJXg
g4rm7mTXucgVNXOrzlj9mq0ekm9j0AYKESlUQtdCVBvFCzzyZ47TMVFQVJBYQnfc
v9kqliR0gKn7NZ3UJAu4kn+qUg2kD/hbVNCwoxYYJcaeSG9+zvrT5U7Kokx0bAM8
daysfXqyYN8nNqsRZuj/Q/Z7X5ITNKovjUs2imJvUvgz8zhyPLYXqeyH+vFdF3+Z
9UuJM+I0A1xFcGu7u4/dhdpeMcHulf7BrIwytj9MXtdteFbnU/TdQjqreprMfNKd
Mv8mjxvi+4o6OXF19ykJgv43ysLHDKa81nGxUJEi7Ra/xs+hU+CvXMMMVbfzKhC2
P8eXVyxuzr31m2+qjKtj2rmb3ZA09dDGmV7kgtP/Nl/kMuStZEZz6DZ0rEDJOAn8
2/v8sRIAGchycHL4FsTcdIPTdbAaqkhL+Wg/dFZKzO2VbPsyv3KWZmhnwN/Bl4Gm
RUykyYBBG7herey8ezSO+ov4KFAXKcsT+zqLge54Io9eui7z6K+YBDmP/TUXO1Ck
fP8osr8wC01np9cMxgK4tYOkskxaFr6ligXKLHGP+qk4hQgM4g+YLOU9DUBNpqst
u8W8T/nVtWlmwNJ+S7Md0hokkV5Y076IyL5PqMB4IB4yrc4mTIIkbsl3vvQc46/2
izWAL/609+6W21Pfwm4mwp8ttafP5oxBFlx0rL7wQFFxnmMoItgcmLLUV2jtEdAO
btOLKkF7S9e313heL/K8iXYcv8+wPQKv9KqSxaSaVISd3DC1wtaxL5C7/AoCGDXz
DmI+WgphM3bvx0o+5FwSF8UCjZW2c1S8yvcEq2RNmom1phfTsK9u2HciNVaPLbpa
hiQen0ns9C0mfeIjqaZz4C67Na/cQWuGKOlgn2yAz3COignt3T8h6xHbawDyFJCV
P82Jx5iFlOM1d/Uq81nGi+/qllmfn8TpNayuL8gYvoZcocpyfPaMVv3wKFvG3TIY
fLtBNdKdANnt7orSc16iPYPOE1IxKGaDT9X1aofBTK0alTlO4rkvmp4VLnOK5j9s
Zx9MoskNodyj9PTeeD2RUr9QvJ4DCtFZw23ZXqEE02j2g1w50czw9w/5/q6mWebs
EokXreY3h2Gus+V36JnpCOo4fZ7PYQB4vNlhZ7EJ8qfEBKMDttOMuwZMXEGw2GAP
bVYnYfqwH7SnraM407iHS2uFic33is8EiqLmZe96/hmFhyFVg/EP1OIG+xL4SJ1d
/JNLEP8cERRq6ncEUpgVw9Go7PcxyZTxKVvdWfGi09g308NqMCcKbwb6adHaJ3+0
3StFmVO3Y5sIb5QwDN6fjhSOsIAhXppREkMKk/y2lbQqVJi1rHeuGwwHvVSQcneX
CORmPJqR10tBMiqF5/hnAQynW9jsFEzQ6XqmZkLfKXw2tmIwAb7xGQ/oi3RT9zRP
5Bhqr3Y0QXwpcLe9q/DMsN8aQvW+gLUW7r8pDpjODlEr8BDkKjU1VZ0heH3nCIew
yfS+PrWEdCuvV4+PNSUgLw+Tbc1SThiLT+DAtzN28KGwQijoCR+AourYRSybPUZv
coy19alr7qCROerX6JYvu4yR7/Fs4cYzdFoxXhWquFLNT5QLnUmLXbQA41gCup19
fezoxmV3WEHt6wPzfy3obC3aB3yqyYMQqI2DjL0eefWww8Ik491QO40+rLa5oVxL
y8GddBl9JZNBXFwrbthi3+NJRjTrKiQWATZUQ45cK/5rB2PR3kpNMW/fZ/qMJfdB
xTBkBpkyHmreKrhA63DLSomx/HmQtFWxJ0oG8LIxYzZ2uItIOpfq/i6mVZ4RCWn8
wDgU7pFqfle7lMcStuOAsqNBPuhwVZAVVaqO0lYzzBSGgpi3j7qHT6DcfyWQhjLQ
4DZPTPiGb7FBDBvae7x5vALPNsGM0r2CGzwnfMn3TG4wEl8d1PD8jRLaJjRPDAnQ
lpX2UMS/zaxbrk+UM6fZc7QYUE20w/QMlhXglx2GHOONPZxZfr7Yaiit7fH2SbuX
ksyUh2Lh0ueK4pj22a6e0/+mxceUEWLRYh/j8wharVN5xmSVrZr8UexAX8Pqtesc
GZ2eRZouSls+pVRFagw/snh2fnzn1NVFYJeKVmMwmSynphCeGu6V6YzKGvaEFnmR
/BtqDeMLdhvU8VqwDUreFEgXuXlOAJ4Gt8xcb9oBLxIMhFgyRJtK1Z7N2bRNyBKg
RGOjJCTBRY5fjrqPaMInxd14/fuxJY9jBVa5ORD1UkfFQoDBRn78TBUMU8lzc3UO
rBrpgZ6r0avFs7X/+yUZ19a+O3UgM0Xc/mB5awVn43ovvmCf32408X54cAS+7Bu5
T2MoGYpWkxdN6nchzePyFThpQ8xuzxlRS7zmwUmIi4Rzc4k4TR9HIy0xF5Yk0RSR
3oddpdNxVwfBa0Rsc60/zxXqrFSt0JsmkS659c/jiRs11BZOBPRMCgnftlL0sNOx
Z+MPpYUBfsn8rmtg2j6pKkUYAZ1X9kcxuAvkxH1bbXUzbn0VSIfwZEqhgoFUubVA
jF8LoAE/iQ/8lycXJBF/uOWkcdVehx/Lg51KBIzyH/1Ql+BI7dGv1JvUAf5E5evN
Sa8etCw9EwijpDoYG+g/gGzckskP/HaAvDJUr4fQ8e5OmH2TUuthHIVnlCLFi4Zq
2MtemNZaIfJubWZLAI9Rcjl1QFMLE6RNNRlp8EVZxSV1m/9n/5sOeSwkxw+a1GYs
Ox7WqlVrXR3hjmls5StGiHHDaqs0MNqj6CC6h12LPX6lNrKGmAkmDuHWhk/eJXOw
tQ8lXG7EIOq2kSyOBxEjmuxdAcNc4i25RXHJwU8/1CHk8woiBP+51zDSXXYnM4/v
q9uJ0lbb/LaRBGD9aWjZeuh00VrbJi2qQgb4JLEqq8apgO9eov/QdwkgSD4yRPTs
VXpm4KbsO8rC0UY48Eumgn+Ps1mpPP7XEK/sM3JVrzaMX0McFA4TcxWDvu+RcfAw
HjmbDfK91IchmSY/zde4LzBfEkJOVMW4GkVmhKBabLN1m64064VnaSye9flbFs33
jSF9VtczZ+qyFzT2iGtdzN/SmHHuGKRt419SOBS04Pr7VI4wUcjzBJJUasGOkIrY
RNTgv9dHWKzUsFn5BBkyMTt6guIdtZsbW1pwcfz1PVZBeqWQvffdRp/kqksbzazI
vEZNoraidIXY2K82iJlJfoF4GVIgojzfAnb1B0yNa804TfQEUyQPget9YlSqTM4a
Fu/b67DjaMPENUjVQfeOvKrtc66RUPmhntGZ94DRUU/GF/J29hR09yxvGfAOtqMq
Ji6C/kz8bInAZqsDD1Ng6MipXYnXP6uRltc0UAf9FdJ+IGwT8M/lA1yQUU1x7mLT
1hQ6LzFKIglrCf2E3B42ZIcf95nNB6Xj8sLtJ5+Q+073agTdzP14rDZoTHjJifgI
L91gbEY6cNncr2Sh3DCTJlqU4t4XKethsC6fqqNDyLb4pGt2oesZMaA5S6+6zC7K
0irXdE/OA/Prw3xKuMZiyly7SYjwSbiyJScdFYWC2+QagBCuq7PHmb8sdH/ksRdI
Hz3575+HQs51YZDItLPFwPKkqu2wp51BbdTlQR9E11mKhvjh+a1cBEJNksGJWT8+
Of3xnc4db6h4kw7tdDd+1J1KitX+HTMHfdU8rYV+qUenK/Yy9PAmW2+WskJfNa+7
iGxAif3v3IQTAya4QrwIiCT4KX9OO9LAt2MBzsmc2y4qZYwxAk0bHfg0KZf9oReW
mqWQ8g6NOKCdHM3553Cpj9ZchgrAk+y3gcQxbIoWNVOEbPFksRDE/oOsXbKsVEUW
W2AJa+4ZcmIkp5Rg9La8tZQ26DFXvaTcyLhJzoYcGuQbL/ZbXuh4pnYpHJEpE0L+
xFGrljtHRX/LUV1JOHvF2PuJDCOTrDUuxFfnqvwUg/jLHkrDAtQWT9411RgurpPs
Jn7cx2/uRv9FD5+YVhdmFK2KT3k0GOCvvUKuc8Wym2gELLwLkcqMov/1lWGl8al2
RTj72zkmB57CJOp7x/ZL4SVeNNiNMYDwGlvAoWsjrmo1uXROzg6eKkvCYLDzGM+N
pbNprPweucDtJIcs8UTGof9lUE0fpAcikYD6mfqabv+83xovuFI6VIHbscqcCMjM
XS4wqPoFz/bJCrrLgjTRoC2uN4rVcHU2rEeDqsZYn8mQhupPSdkxNwEygU0UV1yx
gr32jdJouELMvMKm6k79Oa8vHO+NmwhcqCZEdgkG/OiEsaTl9oVc3pU/sOulf6rC
PoEmFDV4CeE4UuzDlzi6N3gMPtJCmlAKG4cg0Q+uLG7mmLMiF37KZHRlpcyAZq9W
k/R2JthYxaP6QPc5RS3B3u7UdBr3sLaKBKaBhUUCwIMXy5KzGF9NEy4kvxrEVgPn
fBk15yvdlNt2WQ6No+82Pc0jwKzM6phnWcCb1WrpDNrXGFuK4doL1f6Gx8OU2bgq
wcF9OKRmyupYVnR6YwuM7GaxTI6RTTmARch9O1IXO4hgMCzbizr5vaf+55G0yo2Y
cAKU+HJHnO1aU8GzFIWlZd51G2sasSQ9TIl87dfbFGOkJFqgMV/POvZlrJfkOO2b
lMhmhG8REqGgCI8CWkeSNMNtqc2LIwfMsJinEcQMYPwLTcLC2XeX6BMafB6BiTl5
QJZCLoEvhFVZMIOqk+IbrTpzyZThrhos4WqJVQWZ9F2oY3bM8dgT5IEhHAR7Acvg
Fzgyrsr2ESnFq+8wPReThJjyYeEbGGj2HQGsM7akfpKytpvPMmSuAhqGpPWXOTD7
TehEWovigzOOAVHz31Es631J9L88XQVEtcWvccQVDzJRDxC33wgcZOgp7/HGEN7Z
TBE8EKPgGN9GDInnzEYmYqbHG2PdjI3lhJdEfhQ++NOSBiqgtZM92EtQcwB/0t0h
L900sBu+hAXXprya+kgPniHg9A3mSBsMjRRl99FTwK5bvwp8nOn3ftuNjMYFhdYh
Rhg8qXNVW1VHqfj4ocO4TQkIEF9+CfKKN2K52yW/pbcjIwxobKBXmvHRfCtdK3y3
3kXjJZhU9/ehfZOHq+UGmR8dtdcepJNqDU4le/LrqnwcGDo5PAoZA56Eu0MyJM/A
eJ588l/wqZ7vS5tqXnOv1MmSXN64aNOMCDYC5FNvMxpBHi+/Ybkg0dYzF5l6bbZZ
6QYtZG7qyHzAvkeLWZZvV843VyYLT+i3Gj3sfPm+LmvnVjHrj8CauV0ksS4F5up5
n3JYgrNUrbttJTUrQUE7WpPdLAJc8ya5/eqInGUsu8S7GnLc+6MLJF6uUyZ49S8M
Bci490hSYBIThJQ2RSOhVxyDSDmdSbez7Mp1z6Py9RiEZcNAYNM51fX3+SUhO0Xy
CHkZz5ffnKsPRdZL8ZbcAF3SEVQnu2tg87ta3UTJd9XGqenFfuhM8vIATJAx1euk
GklcS2U1dUCRmbjHdEPPPOYscYMepcww+vZiIxDfl29ysM8764zJoy0dQstojvmP
f2+Fzo5VSb02HmgVJBe4JdPjo7yLyxTeDNJuVM4sjWX+opjqym/d4JXWSAgYW8PU
bdlSQIf2FmW65R0TLxDVvytz8h2nvzW3VRW01HPf9L6ksmpqxXFH/ERZ3wM93p1R
EE4d2zw/wRzDBdoR+f+/kT9eMXH7VuhpcT8qR5kaglf631sEUxXqw8VLB5G07eSp
Aui2LAH1QW8N3xiDMbvOE5ncHIgdWJgEvpDU8dVacb//KaDa9NO0IY1jrl3UCRz1
/PhGg/SrUz1m86nOQkDn4taqu0bO0igonOWgBq4T5JwrTuHNmWqFM6unZaSPrEom
TBhg8ylpTGDtYfgJFblsS6+3VjPJxk5nJ6nA19YKadlHfMplG1mFyVegVRXJMvXp
YBu/4Ti0BTSEjX1Uw1xOOrjnaL6RuewuyBZi6FJpTmuL3VtCe6cLpHvzHQ2BZZEo
w+uGOOcPFU05yC6WYr2AwCm5Q0Ne5b0PKvaPsvcx0M/IYvsidrkdOjPQS1LyeOwZ
rDHNSBnnDd+p0HB9XVNlrCSomEpfF0vjxxc4/mUc+6lZrHJbhNtA3F5bypYDmcRl
T2s3toxKRnac2pgiEPt9KKZCxFaoauHKX2P9YHZBZ69guAc6/rjMQI7j0aVMjsYF
9GLY+yLtgBOcnhhRjZ+X4kxGY9IquuktnJflioYlYSaaQuycONe8Qrz4afTpUt0R
Y8hwTUYxUrnCXYms7etCZQLYkYw9LCl9mgv85MU6fe8tReyUXHdfrykG0sA020lX
3uB+JhRNIxE+ZB65ygoy6ReI8BzB/qZovQuy85cm+e44qhlA+Vd4hPDnm4Zud3xD
PWeB3COypgHqpxihFWvAuB1MEsBA2tLVs41pnXB/7ILCYrhVMgDgqcA0hcrptm6f
llAQnUFOBsAEy7M5dxN/Db4zmplTw+jHcHOxCS4foIjzBM1Tj63NG0vG0VVNabSM
lQIY/dZCcWfwBykUqm07V42JOs4XJBSWxqq7NggoqTYgg2m1hKZ/5Z+iP46CxGMr
YZSbBbuo1TLP2SziG4GJiAb85l5gQ7+EQZairm7ArLpD1yoTz9hnjfVNaLi7asAT
mhv63vf9Ug5PTH8rmNLki80YEBYrazlPZF1lEu/bDF9J3AU7d9JSw4t5YXNTz9n5
RbIKiTtScy/13m1SE9kIPkmWuPHZTw8BADpcg2MvUsz4x8lRu9EQvVi39fH+Yn9K
6TpYJ9ZxlD3s5yuP/EqmU239FfrN4aGbHHbYF3a99xnzuBTnr4UvdOE4rITFQQ7p
mJTukP5lLlavR1nv742k2/17RrjxOoPkNs0bcZhIsS/AuGQRnHP3msjL3viqCj6E
eq7QUs1FXFbCjKDVHjxlN5NlOOJzk7C5YTzVBV1rFzmSAPTIInHcviT7YnWMlsga
+sBg0mkgghkZBTSyrtxPJptiMZ9x/ZjyxdjlORDtAIuihgJ5mfGff201wNwml+RL
Iksq9zkFe6L9xI1GZVaExFX7Hkk5uKsuqdDL9ULZHSr+pgdjANvvOcF/ztw5uo1S
B42GymCgFWVXqsixJqOAdV21g2qzQ8A6UM/oR78oyHtYnR8jdVfzIuXF9qawCX+n
CeSxMNXVzVr6CCgDGlvMLbk4P+w8M1ImM2XjV9ZT1UQ4H96iv+19uhT6a/dyPtd6
uUbXlPw4RVemAl9j9ayuoUGwvyEt6/+kilPqpN65EsOwEdE1PAp2kkvfQwkzfWh+
CYX8hixdH/XeWvofn84OT+1obpWSGUVz4EGO/Oogm1Z5JCBUpzH4OoOa+JS8jiZ+
872RdCmF1UEqvcP5B0pQXA0xGMzvJJao+1iTE4P7QHqIwtH8ETXVAZJODsy16V5d
ZR34KeQDDwIgNoW2SzVS82RiCREvklMPD9iR1cUrWJFTiEDsXTVF1e2Ahu5VqSlz
FV3mfS3Ts5lRjp0/2JKxvy75juyPsQvUofyBcFyINQtBCp+CYqouLtzwk9tTwUT8
k0rNtI7aZ4p1zkyGANMkvQCn6FOymEHCiUe4DS65SbnN66n5MhwxtKz6Ycrl7yol
fPPgRoR05eI5bxscXYrw/zmr8032aJzTRwW7j5VgwD94ua4DiXbP8xA0fQOMBIij
4l2n1XFdtA5pCP5W2zJWzavVEBRtAJVpQPlaKqnKSdurIe4jdIxIe9clYOx9f0zw
ofYXnXQpewMTtHB2VbPlk/yFNw6X5plPKPDgsAAUvYKB0Xj+mY/yBghXnrkw/N/g
i0W/7ibFpj3HuR3tJVpy0hiRWZUml9qYjkNWfFA9197NxAfGRgaZYMo8LF7SWfzE
P0/WVDKDSyMEktMhp0+omlfvbMJjUv3V0Vr4ycdYwyCHXRQ8+dW8YYNeZbxnz9t/
Fv871AMHW5AqwJjds3vhfevKT3bTDFbxmvWixaY+Lv3REVRAwstsxweB3y+NieQx
RxYgg/D7Lc104NbU0fz+QL3lNXlraGFSBodI842U+J6qKYqrslZYLW+wsowVeKgZ
yBLbOPUPAqq8meAwrEvPWEciQUA4XWSsaNK34avOvzhsafMitLXZTpNYlbhWIpc9
cTL61hyj1c9QClquiBkHZ1wmdiNNIF/3p5c+F0IhvEc+wVGqSUJ8MJwa1bZOkb8n
sHH8ToHA5tcVw0ygnf6NwBIGLQoFgjznruaCsqkhS7+GHoNHTTP8AjKwJUpe/f10
Vu75uZdtv5rwE0LHnAd3TbQLYiFq8nve5SwomGU7YVbm6F4HwoGXGthaj6eE9V14
ufo8vFtbTxaQp9vFMY1IZYi75jfPlcHXQrHfN5AknKBi+GOkUm+BygMHvnC6Skks
Fps8ISoq0YyYNDF6YS+Z1SHHKm4mdr8sUgxEHYwPgfAq/Zo7wAS0YGMUXTLRBGLH
FbtO3lvIO9/Qo5rdE50OFkPtJ8b9P+GlGiZ1oTmbZ7BXBdilScg++lzfMHSGpZT0
VfuZpyw4X0z2ERU294W0TxMmY+L6zaM/yti9Mmyyyj5VFLHjm0Od+G5trS5h4Vdm
aoB9arjiB2sbQpNj8Jd5+x77zQk9qfS/qfr1RQEyu5dsWveKNgDioV3ENBqpMO1a
B2y961Zd/EreYT9ceMhkI4Q/kaCHVpwp7lqcJlkN07e7j1l/BSMpWCY5fD3OtFw8
qkwpqsDrsG6xumxWzH1Rvp5R/hmibYTH7+UiQiwIN+BFkd6bvU7n9drVPptm0C5D
d4IAlIXHbDk9BM7XSCav2+fmMK9ykMflBJW5wh9TsK1xXfN49G0i9ndIYri+SG1q
raNszzVRwJiklILUaHyFbrlidvPEVqsxbK2JZfzduSJDaXoZnV86LhguUearpCoU
2lwjwJXseYjzVb3205yfGx+Uq5j8mcZ+fTXXINinDeBF9xbS1s7ZcdDA6h463DNN
2xZUuKXhPS6ZYuhHjtaBfchE53h7DLC2Sog4N6dzET0PvkuiMKm3d6ydsnSZay3l
XUdd4K7Mqm2rX9qJlIPRuB1gwoOqU9vB8sEu2O/IlXVzgGVzIu/VDhZsnWBHwONz
Ucm7rjEry20b8xC7V4q2m8/xzJ+iRwWQQp1uIKtfRHTvBtDuHmE0TpEr2xfC0ON/
cE9t0hlziAdiDyJ6OK8ZDS4Jcpk0n49nbRKjQZ4mQuD2O9jYZz8aIFyEvQjKaPzR
4s6//UqnLm7U2Us1/McSzf8dIbXf+vnMNWFakRKmCEB4NQexbeWAItSydkEUV0X/
rcJm8JaW/kvxi0ZJ8WH544eUoosMqeHU2noy5owO3NRcqSmKo7eNvwHHlxjWdbWn
WFVQs6DzYsaMnctQb8fYdkFZpURtsu/XGzcwYwtUGHnXgU3GDU2+6RmU8nW7V9Ge
jp5ZSmDlLCilB+zCvw95h0Tb48o66msRqmqlnSfCZFDGaJUqc1hmz4uBgG6BkGKi
HON6XVOR6FnQDISEuzwZZXHaxwuNeNaERHgpRpPVxM/Oo5vzzErAqXzAfiuuiZpK
VsMH2CMFJKmbpf4cZO47gz843pyhVy3rExdcKhwTxA34a7ori3lZMH41KKWabEnQ
v8Ttlqkoyvtb1wRhvRCkRE6Roks9VPjBi+xCUeNjSVIYFCkLFKB3ebZIw1U7dHZg
ZHRSoxraTc7GJfTo4UiN8GhZ8xRbj8DMSeabLXF7XV6Qxh1T39cYd64HMG7F8PPS
u8Bbo1/8ZoZ7X4s01aUyx4495gUtlGHwzRiRHB9kslOUBLVGshzrRrlt0wG1l5+7
lZ/KtMWLXeROhAX+W+dNDQ5JWFCZEifEF2fwSBgO5Wi9cOz1/AnKm9KuonGn8Ngm
MbQ7TDIdmF7oSNBssn2wU2xP/s+6zKaGk7+jK1MUzKikZcFkIhb/dQR+7k54H1ky
PpMS+FE8B1xylxVYVkNb5ayinEdtzjqPaiWeReScm+LA2oeo43U9LfoYgJKmJF/3
le2+5oIPUgrncpRklqYfK/LB3nss7elkri9r2RCcvAXbJ3HPuXmZPx56Ifr5xyXd
wIW4y/V7Rgq0NqsCtDG/Ie+FOoJr6DqN6WvYeClKgyydaqyieg6LL4RZPmEq4vzD
MfZW4tlr3UngXoN9/ILnNNvJHi5p/RMqBQVk+SVmvIFTVqeFSDCQsGJiF35r7Ea2
Su1LgVcTVY99xwnTZ7Ww5WGPbidxm5yT4X6pvvhdaFYPNRjegmIpnFl63A6lLjXV
7/0T6f/HrxuwjiHqZ635cnCoXbF7PZVSM+I5D8uW5hM21VvmOyeVL2GMtNU4SUK8
SBAUVZRN51jAHpVwzoRO7is5YO8pgl4lCm0U8czr7n3dJTtMZZOnV25ZdOq4Dilu
mDA7hi7AQ6SoUAyZEVptRn9IqnQGrKeP+g9Mg+LpWaiXa25b0M4XbzAcjhCyS4k5
mQ2xR+fP7+F7NSWJmkytrKc9d1+oPuSNXzAvudqeb195K0rIOcKsrR++tlSBHO8C
PNXv7pLWnMPoZmajGFTT8dTUWuuPh++eH+ci7hSnnKu/mdLT2LTYH7SlAZwq2dNE
L9wWnbQyIrDjnodyG/3z4MHPXibWcwtaxcBbJcBp0Gw3hAnsNmB46Qlyn7u5OUsB
bJkP2t5bZYQaBK0DTRx1T/hTgFH6RYn2V7HD4ydPqype6rk+9Xc8wzYJa9QomNGq
BLMepwNf0oVKx4j2MVB2ps1tFW24iM+j3BGHmKbFgV8wwN8K77uonuDNEjlXGB/2
rU+7mLjWwMWc2LPPDRMpjUQ7F4JxGeXdSroyaCuFvglDDFmhaUEa71KvJqfdu71D
aNCQB+5tB+nSeiOB8RfuakIFQyazKYk3Xitp5eYoBNywTYRb4l9HDzZl+aoaBK9J
joQZD1+PX+Dg9v5U71YrS8+iqx7qa0zBzm7AYfEP6VHpjSqt+vJVNMuTfHhKlzJI
9o+YR3ga32tBUGHJ89q/+Bj12btFuwLMdq1TOHV1VGyw6joTzneN40mHFUWXXkJu
aTmwJO5o8fERXziqGQ+Kll9N1dwAoYhnlMNDFM9uw3SopW1won1/vX1JWBpYUnYm
S0FNO6dRQc6b46QGRrAfHADjGahpQmpAw3RmuOvgAfQomh/THO3GCftNnPTNHWtn
/sl7f2O5qjtKkPmHaqXbirOHIY3+YK4W2UWpdN3kF8sGwzbc/SQFa79TyORmTMN+
/oKcrMObwtjuGKIfpBndtzS/Knh7JYCRv1HjY4SXM1HAAY3mjsIhuJYs4lxukqiK
mkSSXNyuGdW8RO0NF4ZI9O9PsZ5fiLADA5eRsyXAUThN0pTMeuMS4HUwEvBOTKzv
Ri6YCIhPca2kHgyX3nv8J3ll7hL0idjYoZq1uJjgFsdXkJWxRpPtW6GWpi6KsF1H
ZfGf/PIrZIEHfbUyhlBY3cRSE8OdJ5Vwzm0YfRctekS7qZPzCjSr3eDiExuprwXY
9zqd26OPXAdCNPEUvD7MB/tjve4UZAXb/tRoU6ddaN18YhnA5dPICUyA1MFVvagn
du550q+xzo+6s8doqQMzBvNpVJGmnZ7MTYT16z241UG8UfsDXGP54glZTdehctLk
yxyNO+v1ibFDiteSIpsS7Gb4gcxTu9LEwFPUa0FbO/AkclxhGxih3U+uuBb8cb/I
Sk1DobBSq6TRRGG9HsS85pjggGA1IFmaWeWfWQKwapvHiE7YbaBlvT+ywAvvizeS
K1id9WAq5paeb88lpTlUjb0+YytNWUDqvT6KTMgYPb4R5iSDQwAbh+zDrRyzTixY
KpwzxQ5dDQ2eyxTKK5cPuRDIOQpmscJhpLV22gqpsvpGdrJG9h95zBOTAMkI0ZEs
uZAgVbuWfG3Wv1c5lr3LkSRQXuomq5swN3VRzmZwRWTnH3i1jlgaljTYkhFIJNMg
Z0KGjwQufbtBYiszguDjJ+WotVyf7QylWfFRbHJcwt/P8vaCJDhHVVy49SP+jcYt
uI2vC2D/wNC97wo0OtocEkQv23Ozzgt3e+YuBHgK+yZqBKwanKv07WaldyvSaWD9
jtmgs1EIZidg7C2rPvack5h2yLFO2RDscFANvG81kuprN7jZz/9eXD+S39XabqNz
6Fk2DAiVl3cDd4HeJWH5EZmN3OlM1zuq8KOxA40iIbrLDV59c2SnTYNSh4y4s432
1hDafnqtaH8I82UEL/9L+GVi2OHnZO6w2Ve18b7zWQ/i1Cd4BITPeaLlF40LWc1R
tLfNTbh8PsSvjZTViPd0wxKUx7tae7p68SV8X0fI0pqkrk6WQAhhathW59bubmHG
zpOuYKICmyuRhXqWCh7vuRpng7YYH2Uch2wAIzoHP8nqQj7KKuOokWuB3hivG/39
7nV9KJH5BPCZqevCLz10vdiWX7vfjjsx250Gu5gGiUxpgTl7RSm2pAJ+srs8KACk
2IEIJsJVAK+VMljJK+asCSL07F3//R3a+T2lZ3RyHqdH8ejKGVj9ncbvHeZR9KPA
mHfhxEuKIRpn2LPXvBSjMBdiFEu3Nuxk6FNo1thkAWaub+pguFdsLOGZweaTJTWD
rKZMW2XzHEjYnRj+UJ3k22XiptGnWDm61/OdtFvVpCzmt0ihobY0Q8R6OyIxRkw9
8p4vpJVGM6DKB8fqITO3JsEzW2xra/Y52CVAcU935RA4nLzrzjE7LjXC2fryKoJo
AQzlF3aDagtVLsq3i9TBNq8FXBTRR6tMTi1FLhGM0soi5i6vcDh6VsWrVv0mc+k8
dV4qi2UcTu6XbdAn+cONN8et+7xRGq2vhSz4rLGrnehNtLlpEFlk1bImdS3S6FIQ
6JH+eZ7XQs1JGDZFSC9TT/RVlTEi2x2FbV2Twidsnm8MW5OfYxVmV1/d/Ryw5Vyp
QYNGJfWmrnQUPvEKRf5DOxLZjRQ8c7Q6Mxc3KEUlsVBiqssbJcNKm2UHcdTS4F/t
FEOv30tgkD8tSswIj70MmpWxH9vBE0nBPEBNk6DntV0j2lPiNFMZvsJGyEUnZXca
k1R4jF9DsyawuYA0VteSqTn3SBeomIdRslIEPZCyUoTXsG9brgL56N+IDcvsvYTN
aoeGfbvEJRxJGAhdcuPjnDC0yzUhyWjtT1+641Tfk44OC2L9RcTnWjkicK5xhlEa
kqdsY6ZBLH3LkCtxLhjVhkGZ7zeKl2r24tB3VfA2aKGiz4X1IzpIyK2yhEX4rviw
DdKJ7rSi6xsP+kOi9uIi8/HvBVSDMF04uSDcpj8TsUJfDfoxr/gzDVHRZIlclApn
hjHU8HtMqLzhCQsZ3foZeQl10mkRFwjCwC9fvCL3y5toFCBlj3U55Xtdsx0t8myh
dBzrsEBHSab1pBiWqU4cKyEbHOmBMuLxs3Wy9O4cSEiFATseDP+JkYM6jD3eTyfZ
xWDeOIkK8KYQvISeGQCsPy+PZiKCqhW8NIbtsn2CKHmMGR5fZRRP1EnN30IUvfBs
vtzgJDzA+r0PSNUQO1lXgnSUTBoTE9MH5O0PKK8gfrzLv8WTh/kaugJWF4CcdB7a
hzhvv3xddbWr0gd5MpxAdVCHlx7frr9MQigZ/sKEgDsJBJ7jCXdr8Yweqb4pZeW3
qM3OqAQivYKdp17K6IzM2xrY3vHn9GkhxZH5/BNkYB+Foq43pjsM34i9OMxlRjAo
NZ1rdgwAr+BMl7rV29BYUIPCIvu/B262CNd7Tc4spkWoLcvlk2EEDYDCsH3dGK92
MVmnlxk2YheLuQrzNQ1mmqbYcMHKCQseniCbsHJPgWTeKdG6Mc0s0la1gZzWe8+V
bEuCysVg0l9OhcLr/aRKVTkbdnWcYqNCAJ1ztUFwCkfhOagfvlMbggP6hLcQrlG8
Draa0/vEHOUUWVZ7fmj+qN5xs9qOej4NiHduSkAbsLEIyqMSXpyHOPV2H4oMGyZR
4D+ZMCHwVnb31ygGOln4gei0nIOb8HEW3qlS0GPxa4zA9m5LZ5yId3ceY/bwRNWU
eWkQLWmty5S/aikNUkMzOvAdBdYsTN32/dKBq7iUeprFdOztwGmI9j89J287kPIe
EUO+vaL8KHU/XFc9XpaECROJflhDoWKyN9/A/0MDZHmpKD1ButliHbB5RUcUVDDl
GIXrJYsZE14GJTcFtXNuJXMVZA5F74uJH/0rB1XNOaFCwbECz92AbDSvL+84/uOF
W/9yOh1djgoP0RaLM+BYYS0xzE9hmyiO07tA12CGhdukEeYbX2nKTZl6KXCwc4CM
M3QRo4pUjr4oCLNV8LFUfNgN6OG4DGRhXGhNRJYhym/wfcAJJkayWSLIbJ3a50GJ
WaPAuZwjwXzlaO1rCo1xO8uS9LTPbCCfwXMkqUbHHybjg3+EtnUfixSE88hFkh4N
4kS4NHIZDvqyIgkzfobhb0DQoz9wIvC4ulWiqATrqFkKdm6qywk39D6lF/XxgXFv
0ZrY4dWRTABpSxZD3VgGJQqE+HUNyVtD2JEHGNCCvJVBy8pt3McZqaEUEDaKdN5N
OYIkpLHCAOYw0y3e4j2nJmyKw5IYWLMeFBNdPgWskGyN7hZa2VFgmQhH0x8EyxpW
gpro8s1PDmRQd8eJcFAXXyBCz9JpDmhB/Ax7rXMz+A/18qFNmfuEDYkDoRuLnv+C
+8WBm2RxAOYcO0oDgntSxO2HANtDpbKcq8lQFEwif96SSktuFXmlFUgc7jhGdaB8
XBwH5yybN49HyO9trrwC2OyBxYgU1CJjL8CpPAmjjjeW8OXc8mptWeSyVvxrnX4t
wi2DWnprg3AhcSn9Kq86siAYrxJNog/F/MRWn1FggZ99lHM5ij0JHgKd3vm5eaiK
dYTrCAu09dz3NtYVDQ0a/IKj5aNsWWppDIDIp3CZEK6KAUG8+qcuN9MzGtSz0fLl
eY2dTSzYnJWlgdWsc+xr+Wmoj3TlZLPLuW2jkG4GLxqltHcQkZ0rW906F7++Ww1Y
u40KwgnLi2FDsPlkTD+SYh1lyvirwIG/WWKwbNXb5+hSGQPG1CY8KmgUktFLYkP5
a8V75DVkXgxGHTWzoRLaa1OBGGJqdj61hAsvXz1XnuJ0/QQ3NwTKdDl/WNU3kvOk
1E6jnsxjdGQ1owBSUB4tYHfjAIHWdNsZpnKqRYtv43VNOgohwJPiNbTAvlopY6GI
8itTAQxSOX00s0cF5FmUOvwl698Wt+CperGdJ039WAV6k3yDwgEba0AWtuSSegwV
X5l4xK6xYQh+yS/u9dvXsnkCHlzXXQvO8rQzzoPBKePS3tvQHnJVVf3OFmMZ2Ns7
/+voMMzEC9ZtGRxxyRJo8fDADFAYFq7w8rU8VAZowfua19xAA5D8CPblUbq+icR7
m5lVrIb/Ql4icaFx9/chhAJfD3lwBtG1Oe7Mh7b3Xuj9K04TJ/FijWfw0Xo5Q19h
Kt5O134St38xjC9/xCFfpbbdE0rrkY9cSj+Q8cqdFbKPpjrUxjOYmw5iZnBhC5nQ
2PH+3myc0mwzp8lY61fXPpL0HDrt6vsO+bIb9hh3XbLOBebHicjxg+HYzJ+FjUKN
jlRr9eWIPoj7xAduv8pT2+jxRCWwMJfkXvK/GfcLE95C34ymON8+a1Tywh39mFpr
mUBW/3CroZ3giV3XVGHM6k/80YL/Pge/4K5AYr+dtZXuoOW33I/J1Y04RAfjq8aS
7zHVX8CQ4CjgQ7tMk/0JTedDOVDOkXNNYMd9N+djF7BUqwC5sLLwm9tdGOVcvXVG
gndSie/akpszjfFVW/RnzvYrwYH7rF7AD2RMPgsYgzwaVLKUYcsrfcD4XjT6scRy
ep8PPWjI1T5kh58+W9P62yXSwmGUHoyxvwbNl61pNw0A8vSzBJBaULBFbaL5R21/
J4wMjEoujR5AAFh1gxijgV5bNFNKyRfHbuAExgiw7ecE6SU9I+xy810oQFSdmUtv
U32OpJGAI81yesP79ze9LTleUl5QY3tdYfkwpaCIyIGsMxvgff1vEnG3mCf89faV
BNRvYiesTtuB7y3t4po7rihqvU4I5s3kzXHA1AmJnjGm9Jd0SLqxMPiPiAWuAeMb
Fna5sQHYW9t5lzHno6n8ffdSGnNikXmHHrJkGPPdQxsSmgIYxxESk177VPPkI/pv
z8Dm+JiFlV45aRYLkT4KO7yUVF7KSpA3k2cPbER2uVP7YFHIk4T7u/tvYj/tApt5
whxMEkHpLMDyfcMCGHuna2I+pt2/SBMf1aRppt4mG9wPNvmuOHhQF7AumntLheW/
Xth76HNh6Ts2Z/rkxzwMOrg+kUnfixf9IWH3mXUgLtC0dG34wmo3Md9DUYwsvGtW
JkrdGzQwbd+vzxckB3h5xpNQNPbU49+x0BWjKTrhOfjsm2MH8iglmqkmYCfHp4BM
vrORo1vbphRvyoOkQQjY8KV0wH198ahosufOegDTIP74ffrXrNSmkQrAapJoEujy
d3jLZCF97rhKR8kDt4T3xXsNXWVaViJjB9ihsio/H4ytxc3XNajxFGxjRfle86AW
GnbFYej+v411BFv+ayzYeV68dhQ9B7ju0O1jO/L+Nj+MocpYtqVkRvbOTt/pjXdz
mEvXjyFp8+W45uYa6clSDpXfc5MY3JvRC9Cj0CK3AWEhijx6y4dx2jpFY25KACGE
RWaCaQ+AkY59MPasZ5WczIFA8xdCvGDQNjrfyiUoMl28MmoIodspblFAwqULJRiy
+hfEAPTYG72l2Fb+WI2ieNqANxs1YYBRilFeDhdzufk0ueijQN3wNDxS6jXrlrTb
yw1jMr1QO36yF8Bgnq28N9nKHSuvQ40cJB8APvVzxbKoBlhlHigkah/efJS6q36j
PdyRt8B2RdHgIJX4oCKE8CdLs7OOLZD+BjuH/U1aCAwecSbMrnqZBujB2RMqk9Qa
L8/oGW3N5biujnEUI2pB6ThafH2+sYuYxN58Z8e4XNyTHJslSTk+qcsrotInzNJE
hVrkZ3fWtg/weiztIdiMOsD/xh6A+yvKvZZ1I3qVa2EYu8YB7RFHJTti1HKm68Zq
BCtC8TkFfh0kgUNmk0ma1Qh+IrYTTUd1e2Uz3sb/DZsqkp/A3CWdjm5TZar8jGKB
TIjnFIYgzqF9SoHWt/rCcBtEslvDGwIyiKhHIGvkC9t/2+ZoFpZ19reCHQCTLbXm
kv3+mFKBV09yiwTcHbro37iij/tZutuCY4ZcbIYjFSbjIw0tB6f3Vce1jmC9FDMi
gTA8MsPTB8TTHq+ZQzm7DJfWgKjQyEP89LVuv+B3oA5lIrD98zIWSAyB9lnLEQAj
uo88NpJhItWvu0a3mW4yPY1bnOfRyIb4sanxeNFHuCjdUZjjAx4NWA2vktcHpESG
jnXPTdCckpd2QElz9qzNHRvuCvOKcDf3zm6Ec/KpYpQjBZGNQL99g3s8yEKOZE74
AFQEltXNCQbhCkppdndgQKLKafmyyw7I8d/QyCmv4eDyG0U6dLZE9RGwUvUZQBe4
0N/9HJ6p/dAtbg/7Cr2mkByA6XGjS5hL3eIE48dSu98uu0+wQSasay+SjWEEWZGm
XuvuRBHXV6shDiatQGWd6gUWdtSEMOcg5Od6md0T8ZC8j3WmRzqVNB8HdUVsNrd2
1R8qeDLDEEEbaxpIFA0dpTGF+R/ST5RFIGn3HKzUbxKOSm+UaquOOqZvr+LBXIrv
ATgU3Izn0SRYSnBqtPK3xhhEq+r8JzHeRAZk0ShtOFp7N0jI+AWruvAv6wiFk9cu
gZRVLuabFGHnXaoE32eRnng6phib66/zqSwpBd5HsnQQoFUaQUjt1qf+sfyvMKrc
GEu6J5JijtYcLuhy8v/4LgHR08+VGxXrocpbFPUTtX5Ruu07nvCI71Myq8qzs+Pt
dHHalHHohHhGpZ5rBj/iT0v60lgvenoC/8kyJt9wi1QekMB7KuFfW0rDEShBtLGw
twR/JedoSFOASGd+1mxJDBuavrducFo6VZDkkfK501tS30W50I+lhiwb/hyaFN/l
7LHFuQjXeMrOeVc0kbqdu1RswwdXIAa8fzX+bXWVUVgOYu5H/rVxF4Nvdn3DAqoP
CS0rfyGQLV1OJqY3FPH4J48Nk5yI81hZzAQsflj9D20dcYOqctHgJU1JOxTl4V93
IX4fPF8zuSw6rCUc7L8ac8Kt+MFBWNey1WUwac1errMhnylJHm/XYJpFuCq+vzyH
ow5ray1zk8KbVLYWslXj/+Pgnel8r/wRh6Eqg6vqHGIwtQ/Rhuu2KJooHwXICjAE
zu3Q9vi7bMqscEryyIu4gd3cojCphVAQ19b0O2ROkDLTWa72WInJaclcGtjpzx2Y
sMS7ZRplPmDNFuWHKTLi5YW0huVFdXxNLTaTWWqoXC+iwmYthGK3OAiqwxFn2e6r
fML26xRDfNuR+IxMqmP+ZBk/+2NUjVEj5denV1wUrv2KxDPB0jiHbpMOY7RdMCPS
0cGtw/eli9Dk3V8qek9jc8noXXMsYEBljOBV39kcbgjgAQtAtyle052dXg2f5w/W
bOoqSr82fD/y+DjmtsQZFPgZEtVQe2F/7nZskEhsZMoB+qUuG8AM3BFveefLdJJG
bIjS3uPRApPCG0G1PHGJC2TJI0MFzdh6r7DF09G8v5QAnwgN2etBagi+bvubteA/
5znQWX+pTRHYPMXE/JaKNhCGyLsuaWZgcRoRCjoHCoz5IisTwEQqnxwN/KUqY0NI
g/NxkvAxtTM08S6pDIZG0mTcMFIZ+JYv2nsndr7tWVoRNZYMIuThYvHELZlutZHb
QVsr7oCQHClA05UOppSdrw1lyli75pRETx8a+vr81eSqYtok7GA+OJKXcqO+XjPb
cKFsdWpjlxsuPkhfZwe6YnkGbvXY5Ur4MslO0q+H2ovlNO5zvXdKclWmwv83sO2k
YlnOYtuCq1iUMcCNZ23IGNzhPv48zj2yScOy9jqGaSRzEKfc6Zt4PIBL2tidDMZ3
/yqFthS3sWV1zeboaOGNTElLSECHTM+zV7Qx7YPAvO4n8dly+MfixMThPtdHx4Gb
Z6OJQaOLEJpUQrShtMKBxOamCx3RSbzeHul9Cf3i76zuPPrPutL/urHcpQJceahH
K7kgG9FpXOASUmIUxqQNDi1sFW1prkNGyfutGDMwkf7mTr1wB6uLnZ7ZFJ2BxSLO
2Unp8CtJ0wvNPleamw7t6VWtXAFkYeqaOcis4lEHSGjV6ISjRqrZOInFNoHHAXDn
DT8F7jD0HHEtyp8fU5BcEc3ohCIPAtTQjSrkH5IQzBd1tLaEKWX98/jVffjFYEVt
qlCW4SkwaNVUCFZWyojx5mGQjhbbEiErEwMhXuRgFiKif1L1ayn3v+/CX+ZeRp75
bVXYf4cUm0g09DNjxW01iJmiX2U1iH1EBn/xPcN/+dca6dKPQJMQ46Hs7ODMh5ru
FW3ndpNHBTHVBOlfLtAzzUZfV7PknNGw9pazm3ynRmzegX/aqIDZiL1ELOyz0Ub0
yHl3awCeqaYnVZ9rGfdGPG7eQvMA7Vourprk1kyt4yujGj+tHXPFgLutLRfBGQDi
BPLIeIZJ/3fdCVsG3lNNX/Pe8dj+hB6Yy9tdm5w7LrHOfii9bGMXxVsLb1yQMZig
9foiybtEconI+XeQ/D6KgnJDC20dnnZKVabIw1CKZuW5YMr7dqV32KMMvtlqfuER
EdjGbr08R85PP+OIET6D0nH7dKKBk+iOgIv/iJzGNfeaqaid1SELl+d9G5sBN6XP
eWQRAWc9Mjm7167+f0/Kpepmyuob2pGSMmbpNt1LDIDNiBojJwAGk3jWsJs3FIMy
Rfewr0KRrg3OAgIPEvQzxv4Fk3yA/QMveAxNtG9/FkI0J0NTJMrG0071MUvtpUnS
FNXaIcwocsdmBF37VZZtlVubJjvQjQXp0DvzPHNvv7uiP8yOu72c+Au0WDVtJS2t
Z98MCLP1OS9bdFFLCWb2qXYD63jau+yIx0ppo2HJsKTq/JkynFRXA3drMqogabNA
zTV9MUR0T9An9PxXaWR7PixkDW6ZEQAyvY6VLLw2Lv0v1z6ZnbkNmqZaU0wa6GiK
TbF75fiTrPIRhO+kLPUYrGtti13msC1fp+A9lLZK5cbFNhFkHELU+Nx/RhtOEmwy
EKuts9kFgn6f+VtF8ih/e8vDxpKqZxed3qlOJnf5ma2Cxel6vDER558Jcj2rkhjc
i5l0005qk2Qlc5jC/arkB+q1CGVzN2eU2PokIpndPwvlgCA9Hhgo77gjc9LNTG6m
fXzu17qlxaTjysAM9rFocrpwhEWhvlL/GrUt5pYNLF4VRr+Si2UBX21qe1Q9icLt
FG8fd6xXx+8rVFpMwExWODHeaQizvTu7fMDirxlsB9kfFvYhSvwO2HoYWcdIRtBT
wFGKAvCPIte6L/cuLw4NhhF3l+ExKX55LylPDw/f3FhM/derbsxoUqee8sfc8pu9
bm7qf4lAHchF3Pp1n799AI5hdlUzxTCoDp762ezij7YHb90KwEgByNQw+GyQmAUP
IkJiq1Wy1fGBaXnt2QTy+SFBb553rxJ9B9uUFBNf38vL3E+WRrWqdVbTOZo+q9mX
0MJgxkk5GpobVW6fTvPGIONnNPp6DHN1uChLQvbAFL+25Ir+7nFdKZ0ZJy5KQgyh
rJOVr0t2yJaa02XQHCYXe0g0x8gPkbh2S0eUYDfRtYf1KgeOkn2Djn1bFMWK2fKZ
3vFeuEXhuClDxafGzHfXkyX840kfr6wqDCjC3m/KEgzt9uRQuvisvqNbmKGhmEAR
tWjIYlB21NilrT4cCz2QqZAw7NBOCySp5U0hcyWznbGgH2OS1k2/QBkfO/TJ6wuT
GxyZOrvNIZFQTOWMvbxQvOgAFcirQkGvKoWHcvO60PSmA09WhEMlHac8mQMFVC9V
Y6RxcLEV6N3okKIkfgcS3EGCRTB36paLgwFKfy7MlgECaC5ACGT39HZBm2WkqTDU
n1KFeVBBuPJYky4rVuT49sQGUZv6kQPzwC42H8EwVez0Y/Qb+aAhnhMVASFzes5y
1ZPDanmJ1ZUbXxyIzaq0Wa6ZbVESMveYqu6J09luoaYzoKZlpwruTmzaI2ZhB8DV
m1AFBU2KLnzO335kv+Z/0Fv58iQ+iCziKZUs1XkjQBXlqW4XOwNWaA2TE6vFBHrn
I22AeiSCitDOFRrF572UnkUOCf/D6FhiDU/vbyTxaFe0KMGlr9+1/aUYT36p0lIr
jjQBX3bHpwxkLlN91AWzcKXK2B5AtdZW472+sU+nA+hCDkLIvc/UnO6QLdJQPLzo
m8ln4GmjoSREUsre/AjJoORapFpp1iVJpHXKrrqaM9rXVLanGzZfFmkbIn0ps2I5
qyB8tYRxud4XBusy4W9TTPx6vEcenVqP0iw0kJcv9ppqWioZ/7aI/TqvmXPCk9AI
J7wn6UcYAgCteNrd9tI8BZvHqbR0JCedxykt0qqvF1LVksxmw6C60B2tlE3psO49
YvFly8HTZjlcEZv448ADKrezvR6zdcg7Y/Qws56xXxvPlECm6sxcBAeIXJcNuAT2
jEbneLZ/XaHySwKG21EbbLOl++zi1QACNWXuV6fVUlKXNpaegUs+zAl2768orgdm
4SEY+8zCbKvacRUxHasKLRvm0jGqOxDQC6Cz1zqn6jm1VRL/ucNuuLG8S6BIgnLI
LJWe3i03z17cnb7gptuzENn159tn8S6hoOVO+t18IeIM1lg476+nEIBIoiDmPiBu
xjUXMebtl5AXUy1UViloGgU+/h2gTwHK6bVCzno48BuSY3QMJ6PjySs+nQ4X3xoh
4TYVfI73qe1uTMI7fIHuGy6A86Pc+VOw45lwF/vWsOoF7scexuc2XOu4YFtujey6
U2ZTYqvNcL6VvEIMLLsHvYJcLKyizRYXHnMiHUwpCxU5ikj+HUEF6MkP959hHAoI
9zLWN0eZQbAW7ayh93wXtwCaTD/cSeZZsm3GegpX+uwgHaG+7D1vprCQ5Wi43gJo
7cOQAEmXaXD/fZUhPChRlmNm39XP9qmFX6gIMlGhrgsGteXbf7KEdkecJjbI8AG9
xk6rQIR2Xx4ZebpmjwybtBKe0cTm9o7gGEaaFk/c9bQju578E7l7L4vcy3CmZYQ8
f+BZztP0uRqeBh64ToMnAyMQHVJbA/9+Voju8mKLM+dawSzvFVlcGV6Cs6VsbK0x
qCm0A5hPiaHx0n9RbvghrrxvdTCa/CZ7/ojn20G2bwyRZYyedY1VLI4ETPLr+/fY
r0GyuPMVbdVNazkWPG8YZ2BKe+2fk25hqwEGOgNds8atCOnjnlvY/d+k0YKDXt5K
8AEqsPGwhZbXaM+/a6csxJC0QLcT80D4MPqkKlrZ2W8yDapuKijzEmbz0c/uN4kK
cvgum8zbpO7y461AGoOTDBotb0ydMr3lvRS0jvmQRPhfCOu/h7n9Smz12YBCOBVO
XUg9BmLJn/jvEXf8wlrj2mJECJbnco0O1DtgBRSe/lD3glXMXvS/UxdiwlXpHPt8
i6YKl54cc3/xDFlv00TdmK3AflcMOmoYNiGtKdMivK/7ZMF/0AGIZYbZj6KYKNaC
yAiTFYuApxQTeZJu5WjMtr0a4ef5YCh8CgRaN1lmluqrP9LhxhaSvZfWL6zx6EWt
icHuXKpPCRt3wcUGugdpgNAdTHpLeLBSFexYIxXCHgrrG+c7NEM1c99Ws1u6LeJl
Y1jH40mncnzm7Sy8ZvL14PAv+bjUArM67zsw+3IyLd9WGYr0ohnpaBSU8HWWoCrt
j+blOYirmEfvOTqqitEfiHyw/81ztRODTbK4PK0DstWr6lov3JDVK1gfpcT6eMSk
Gd6zH/XCtivH00Y97rpEPK+g02onNHHlYzhZlJApZSWJbOtXu9DRgXhXv073xwNX
9AUU6BbFx26hfaLR1za22Z88GvvO6tHt/kW2qaP8W/s7NP/F8s9ZlOvmEh9IC49i
mobhVkmT6xCNLBxtO+ng8SdKFHI8rLgULIdkDhQELhobuP7gGwYxfzY13yCHXLLG
C4b8mJd/tbpjyIPpb3ZDxaOS7UQNBe/Lb3UqbG1tV78/TmdWwrUJvkDnzxbslJfl
I22XgDYz9bPgemRxuSYTn+e5H5zegkdvJl7KEZBJSyl1m0GLofcMSlIa2/fDSgvM
PzVf4A/E1LxOisxQJoOAmIFouVAx2ThujF41gY0fd3r0n9RBeIJZzK64TgM4VyHd
xjmRd1e5fS0V6QUtMIR8smM4RfMLqxTEaa6B5C4FyAjSLgRED/Kd9GgX3N9ypCuI
XXxYdz+ODg0V7sLmAoneUvkiU8kNh9nASV96I65kAdxUU6uNlwYSdc/YwWoJmUqo
U2GTjOjYrsN3U2mobpvuG0r1vBQ185E/l6Y213lQioT0ZI4441s9E/BUa3BWGdkz
rXTW74XsIGhe+FGbpd9CmOjgu6tpa8ZYHZmdNzxBRbhMJf+WBIfugH47Zz1gN0Zx
3D12FHFwxbbAK7A1Y0hwT/PFaOCdNNjpHzvjddOGyXxoFRnQtRjZgvlLc4Ul5Idw
xSsEBEPfthMSTfjLxjSwHK/PT1wQPp67+xAIyQejVFAZPgaJ2eFjHuR/Q5z8yK4X
cX4Wyx6D01o0NRLyBsp9rQlGuf9WDoe/iBHm1icEMFY/0/kJUAoIYIFWwvVZHQVo
uGk+hIixOR6skUPjTl/czx1MFibrBoueayMLIMDHL6NAshPfiJ4Z9l8M0uByvtQW
60VjDoe45JvVwBmNbgGWyLJ73lOD3REZWQE5k42c7VYEiTRA0JGonO1GLEL0a6MT
R+c4EKO5qHKcQHRwGxXJC7TH9SsGBlbnC+zCX5bnLupihpCqI4CsXO4FyfIWWy3N
6YmnrQt3zgIDAN9T3HO8zNZQkxI5hNv2zA0MWujmP8QtSyt58xyF+3cYOAQws3/B
ORLQG4zccn3frx+2LUs8vREsIBP3YUCwZ8DQR4WWTJp6R3GALfeTwS1wWB55wnpB
DcfT26VNFLP8y7/jnzuBnoNML/vs6CpsGwRgw68EWb7CZRov2flesAtDNrGZkcts
X8G8e8a6G6mlB0QOTPbj9pmfY85XPRJ3/a53fvhKedb/0FJdG8sj9udHa6dzcLqm
Na9hjDL2eMBL/VJrTwqE9O1skPne+qbEaOMKq25Z7UVZsHmetNbMNbpELHP4QdDW
KkovtvR8qE2qLcT73UA+4p4IsuFCz/FH6zcJCC/KL0WSW+ctLmWNOsOyVAqfM7vL
SqSWKcgQZKg35lcXtl5BT5cengas3y7wQgvM8D6PruolD8la0123HVy4HBT775C8
GC+p0pj+X+7h8zvyoBI8MQFEfaSn7GTe97yWwno/hBs1xkkES/nv8m3JEzL4ZDp8
xCJUaCTMQjplddsptyHUSfK2MFY4QT7/YqBu5sFkFbeJ9XmLiv78fUx/GTKuvCpA
kYHL6rdJXo7Ds5qz397HZW6P2cjwZ7Z6AJnNzbRtZ8sFOObxESAnGDsx6rY3fK40
d9KiHjAUKbyGbtO1mU5QWJyP0JbnppIxp9XDExONJ0OuH/Ptj/oQ5Ihe2ZNeZ9Oh
oGJIV03C0C4XaCy1SwRiD0Ou6HLJB+VpqBZLZNgbAP28TAz+VWlveeC8oowgMKKK
jcRJIl7wD6cFio+Ecr96A5JOKGUbKOrj9XnUNfHWP7+gdDuEhZEbIxUqpNU+2T4i
e7ghWcSiYWe3HWPa/iFLD1Y74hZEbcupYQlQAS5dhrcwWRCVoiIUMhrt+HKd93CS
K2O7y4DB+qJPT8DKRwWwC0ooroMKwmQG2q4NlcmnIyY8BgJRIvObWhZ8X0ePx/BV
hpKdQwb70m5Lg5xkaGr6Ze1VCTiWCMRYUJCfr0ctpAle64AMVPHkzFLS1HKJM87z
MD5bgmwcjmNc29Y1QbLQlwMdGRcrBBAt9kjaiEBQqrUVZOeNlZV/sSiaLWXfmF24
0PsjcfnlhqMV3xhjtDW4nUi4cXdVVwNFs721Xd7lmBFMYNd1CHCBGwOHVxuVfgAQ
q0us1HBkVqiQoQtZ6Kol3SIVrD2UkZ7hIxUjFpwFdx8+X/5DIRr9qscRHxgaDZIS
DGsxMdRdZ3XndSpRLTiqsSGG2U/VESCmfp3Optt78R5/R9X3QvpwGuZUpOnOL4qu
1XEHkWXsDim615czbqwMn3fxHxqqLsDkxcEp5vkdAZyC6c+VhoB4X1cg8e7Hq7L5
srZZe23wffhJLtxT8CVvc8bl41MpFv72YnUwLTA1cd6Xq1/2vxvPz6lA9eh528Ya
Zxy19xV0/K5TN/EOYM58IAoXk+CuzrEI/HcYnnQG5bo/lOCFGRU/pa/D1UHo2VB9
hbLfUOhYKurxm3NT6pu8cK20/BDHxIl7h6RqpGzdP0JK/RtQnFgWldKHSkFIxW7P
skKDHSEcJqm44NNoSvXRitHuT/CNsUeXg88pgi4xn1GYAKlTsOTxgW9epc6jfOiO
q2BwS0O04sk1W3nk+sf7e5nY7w7EI05ecWzL3fXQZz14Pwyf5Xz8GiI+HRXeE/0q
tjQSfowimhcUTGvBQ5ekdw1K5usOBtygSjqUazi9pvXJ51IbPmH0vi62trwnko/f
95S022hlPb7B0e0pHbZqZkcPcNYceA9v1ZnqUEIeS7XqdfO4Yxpr+ixCvrVwxmzL
gzIS5SOcsJQCb5N8zO4owgemj5OT1kws9Umet/PPbU2eeetrH7lv37ZlIC6RaQLR
dkt1X1+nfj/jTgD1mfubSEPBJ0eBiOmiauPZn65m3i6MzPUY/lm5OLeIfGsCfbUF
/RzH90QE1KfG8aFDOfVLzqQTODVQp+Q1NhPyCEam4Iglu2bxN6yAse8VUaPAnqsd
SuuAuHE9vE+5mzkhgvVCVMPuB3rPyvQOI8VigfFP9zlzhCi42xEo/jw/n/4/92G2
DN06si1WWl4crEufZ5NcUXcOSgdjYNnhmX9fZDFqIMWv06z+TsyHdKwXxemkOtWq
qkToGe/0N82a3JMAtTa6eoOlMU+QtLOCaXZBRmF6pKZ+YrIniPJX/B9qNguHamAo
A+U1vePfIrwK8f/PTTgwVyfVeKOhqL9LiC2wvk0vdOsSV6TlIvsVPR45YRJMxVAb
2dCDR+Xr0XfFeb1uXAqw/aovf7h7Rr/wyD5fYqHa7SBygXYeLV9oRl7zIlFFddw3
nEnevj5ot8qguoIlbonKkTxofqk5b+yTnyf2kH420w/jY1fn2L0bPIBTzxoLiRDC
nwe8qUXk7yggJqjq/JpH6MyBZeqPnSpRjp2sFrbiBQE02ij4LJGCcH6dcIt1Ae4O
aVRFUhmjrowpzySbtMCU90QC7TJmtvHmrpV02SzJQVgaXZVAwgvBN/kF37XJ/vdV
tGOF8ZWcVp7KWxHT37lQA+jBXunRcqRLMm/+86Q76fhTtyboA/K9fzdN2PSrTzq6
r3Afxjw5B0cToeLUZgE/wtGzuTEoWUs3nfR4m7mPzIZOhhPMwnAnWwFzHMfRFxJo
0yCU11UmpJBE01KNkmdLQQQnumq0NwUd4KpwJ4/GhXAAgXl7yk/Vilpm9A+YzCCd
ICM3tsh406cBjTZwGkNt0+W2oXYN1cCVCXdHqSkwq5+GyN7N/wUPzducVL+wzOAp
BTjhdL9Q54YqqP0CxSxWbqkV+IPnZH9aa8SYguNJ/G5aTWD3Ja5ztDTLra044Yrn
yuXznsvNS1jj8xSjyAPxr5sAo8IubS1yMXNSZahqxStLYFFeMMFgPtXC9wYt6Qsd
/Spp4yTqpZrMbCcN4zOaU8hpsc2lVZ+xrTakgtSu9KshepUJmmO1Dd6Uatx2Df+O
MBojNybI+ayLdOvEY3uIiISNBr61a6kzkDYC1MhSO9Y4Y7bXYAylyas9nogTz1zO
zSeGqqDfEderM0ro5jH5BWmujNxN38a+9TEoUlkzYFmGIBXaNl0ACmvcRhbqTvmH
D8OEgImftNWSlk9w+i2KnGkGcmn3B3Eg+w9hRshGSMcZNvzmb4map6WYokvC715x
w5o7gKvqzkBvCwCV+d4qJjGL8OkxgluW8lawzvDmkG5USf566AKUl3ayNFISUOae
4zTUFSG2Nftdt6N5yGGP2YYzXTUYOXV2C6urhw4w3QfSa+jDPGJcWRnX6igBP4Dh
dUgw/tPe1eaUz/hP4QF5l8I6sHpWjw6F+ql6gRFjDEmhwNiHcciRkwf1TI06xK3/
Yu/BYooMs8WrFjJ0kpLmFc9sANAva+BlKWCien8SwY9CVkUw+kk5tsvoKIKzs6/n
C6YyINGVFawoikM4sgaN5cIv51A4De9VvoTQAnNJOH9V0a0dwazU74znsTI2QqPU
RFbIzHWBWnkq8P/eLuzG//XFjdQSj7k59IB/DXu2Ip69t/hXTLJ1Jc4ztj2eA5DQ
k7OhvLx9opj5PmdTCCgFfs4b3UWLAz4yNSwRLv697z4tf/LnnmkTzQk4HcV5ZJ2O
NTqgbTYGKsvbKwTRBE8Z/G+mvijpLF8pYAcG2maTZszvu8qSrbHESg3ER+2YnRy8
oGZcTg6l37pkK3q3BwwC3RSBJU1mW5HL5MAhxVr2f0vTgR6g9vagtIF4i/mVfcUy
fAn0mDGwhfUQuUxFrswJ7dynWwPT68iF6UXSysOZEkQgKetmUW5stPGUssmGtmwJ
ytZSspQyRqkYpKKt48ApM7HSAAVZCnlfG/KG+wR1v6dB+CLm1DmqO3TOysn+WR4E
ECRcdlKcMO0dsdkVfoNdIPtT1WZrhlC+5Z3m/6ON56PRM7UykC4QXYVt1oq8jKmC
oMbYZYfbIqupTeM3vCz2gzQ2E1BHV0aFwYEhi3jN3b4B7OvkHlNXlUqkW+TDiVgS
99RWTFCoSSzN+h7EiRu7ShqnDhu2hDEY5YV+oxd7xJ2NPQHjuiF5wsEynTFyzY2o
7wLIhOqv+FrqIcxYHKJ9/3+gTrM4jpf87WxLKbHKg/ZjSXwLE7N1lsq4fUnKGCfQ
1TxsF9zv4Xi0eoUCJ8LZz0eSGM9f0sZif0hlUpjTz67cDAee7UiDBEbmUQDbi0oy
qjxDxO6uINc2qy4RgpraQDHkYH6xcDPDwWoTzUwBVLC7okyXiSxdtgI1Ebts85Tw
rtdfbqEfLi/xqMh3APODZVBhH9NXExEcluTf0CiDljypuAgobcnmMc2oQ2DAecYV
dRQp96I2yIo2X13XbUa9UwurIFWyazohmYylQ2S3iloCd1S+mynweGWPNDZUDf4Z
qG2gRCgABLSM4O28L+yys1eqJfB2rSEifXfhNOQ1oKCQjjRyOzQGUZxMQnx4CT19
TgNgvNobSvJIge0Cw5yLmGwrjlI6JThjBAoPkrHXgMs5J8rugL+Sm/HlAg9l2ZOV
3Oo1fsLgTf/2n436JjtShb5ycKj9ael8w93qYmsdurIzD38buVXHQpJpN6qGIHLD
eptGpdieCSkjWnWdtmkJXHne5dwlmfsL1/fKwrquUktnVWgZYwv68JihuiaQn9Kj
MILTwo1rz19NS6WoMKCIF6zSX789QXzqraFzHxkfJjc+MIT3GwRoWZapzK5ZqM2+
/7jKhsIy63Y+HkIFsCI6EoiE3R0DO4LnAW+yjq7UZjS1vAl4F0A/F67eIUJODpxY
Xva/WGQLE/zdYSWNdaZGoZFT8bZRNUkyrxEPLTu1Y3guCFBk2YCdiPKHBushYMAP
ryipVBfcdYkWgvkbw5AEKZeLOlWX2Eiv2/aRfuMe/oHtxlNImvugMQZiSbDGCH2s
ngaJGTzqElGFyqWZUdiAs+/GBd5lo9VXX+zFj1LDbNcvCdaXeftE7W74ZhmISIxz
nysk/0N0oC2ugQsNLNhUZI7LtrXqAXxVcNqHNPMGJ/GIAbyQuEWkHPPl5x0BIwO4
LymE5cI2xt74Np4v3ru8qwp0GqYGqzvfUNrRCnYLHlSpxmEy+NCbVKrP2chPw26N
gNsezg9b/wVaCvjrbcwaXE8p3OYN/dAnBlixoHf/sSHxDY+KPQtScFF68XL8EwyC
c/ox7dE2Cxu4FCRGBsieZizzvNT3qcMZ1JvBklby6WUerujwVLE3rVJSuausyngm
i3UtqTz0wzi8tB+0J96CcW/x0I2ZE5AWHlWaws6pZd/c3DI1sAHzPwbCZ7f5kDv3
dipmxge0G9tqfEji9HFh3vtgMOupMnCycoUF7MdqSf5aUx+32p0V3hIPkAxB4ncJ
3/bexRWVhvRHD023Eeim9XMcDfaAHDHlddfEWRHd/svWtJt70QJV9Bw3fiupELA4
tpul0jUD/2GgDANRx0C8URh3M214Ji5hPxf5NdkrkT3PQ+2+SmrnK++FKg77YbMf
T05VBNuPtl4RWy+E/4kmEKU2vHjr+G0jPRnaMGSoS8A/9HOck/PboA7ejsbFrtKt
iER8at6QwPGPiPvfxZJm2s9/fnk3mNvel2AghehGnZwOw7o81diee+ROH14Vm0gG
xMy9X8KfDbPKa3a6hD6Kdzbd5s0JiRkiSpTCMnm0nMYhDGy4SgfdD3v5uANeB/c4
YPEIJc0R31rB+c9DGXpDE4cad9tWaYa+RwZorKFBrWkciJvn9drPHPOrZBzKTMnc
18FMNL8nxoXwRFic8zH3ZvRajk4lUgmRoL5dRUeNFfxFLkYqKUR7xU0OKv2PKK53
OxDTiUxaSDdj29t82vDjbe8h5DvBJ/IMNptwspi/CC6rd7wO0k4RFF7OXUG85Jaw
BXdzMBEBneUvCaOAYfUItExbCgmVQ7tIf99nBbNcB+Y4ssMcv+2vhyZE5aRLG/J3
1nKTmoPbuRnEG8X6xAbjPMJdkTSCKMTy7v+8tiOizaQsH6edl2j8DdwuApmJzcZD
g7C0qDDBK1Qqe/9vqEHMdppPoYCtN/3xWWTGeBRZnJeDAvbXossPDBjJ9muncOuL
qXMCcv5Wnx7yyea/+5BYiGy/Aa1G8Ds8EG6IubBaLZW9m9OGLOlCb88V8BTfwUn+
9lhRhpywScyGU4Z4ivPwN9NlWZ5iX+7xA/d5gmPtqRtHV5ZtwjAdorFQjGO8I3iF
cxuk7CFNdY2UnvgF6TkixcZrfvVLKNCKrW7JyxFuYHvjpRiHKcVcGh/rL+gT8mV7
b2GzN0fVhFVrQBWrA7t3q1oT9If20xq+GAOjpWZn28n1IhcUJWjFhwQ+2f+lTwTo
WrpynoPilP3BBKaIimFOC5eQMygf8xZ7tveFw9v5uLZ9VY4I2bXBaZ8Xh+69nuBv
grM0B/Wz1yz9mjei1dE4rJiHBqwjwsUcbn7k6XE6hDw875MbhLOowm9tKYR0H7E2
mWi468Vj025x+eRQXXxt9gaInwaYjQyAQ9TOgPJPQB7TylfwUYJ8ADHNXSXx+Lmm
j3oVBjhjGocuzO2D70BQkILJQBPb9IyHFudBWbij+IEO/F2aGQDHy4HM4iv5t5Nd
X37OwycUXQ5nMEvdDaxpHD9wJwZLNgP1Y03hfK2PeOJnhtVFXYZwS4PJOffKX1ol
Zxaq8EgV3FI6YW7cEvFOzcDlN/wEdq1bza7yERUY48nctDHMkhLsBg+9R8ASQubt
JneyjwXCACVLNBcNej3EiMeB3sT9AJN5AMzqevIw0t1/zKx3sxS4vdnRDFQx9TjH
BuNDxuwfB8s2R0uBjy794t7XccaYomyQmhh3fhxSicHiQu5hBwdflSViC6rEKI/n
LD4QOxzqH6DzeDJHnuscX+At2XX4oYyw76u9gHupHuUW7VCfyEm/GrDslKDtPFgA
OQ5cxfINm5NAwmMZX9LHx2qpqmgurX3OnhqNLdksHiBU2TxW74aNt8cs+S/QeOWj
M+lXsJ9wyQU+VMqBw/Kgi4WXyaJ6whzucqCGQ1kY0or02Ny8d2CWgA+xmlNn7AGr
1dBLb+LpQkd874taOA37uOtETUmhN06EXfInNAVtan1Fx1tawsapZZgj6STAdZKH
Uednez7+lvc1jZnMXEuQzCc5VI2rqA/43yrWwIVpOX8V+i+kTw1zUwF+gqenbpTf
SWW1yMPrhVoD3TOVwpwqmaZOJ/CqMddlPdhQ0tqDr6lBw1n0+5zyrL6hg5LsrDKZ
kmv8reo5UkA+6gcBj8FaN6cWH2DmqmF/ShVMwQZwT44wtjuoyExakFdhnvnVWIZ0
MEIvxYSqMj5wuVLzf3MaSsYCtVxwCrYQD6wJBXQrV+5wue3dS6euWXfPlEesIUKl
/tQbYVSuMux9olCpFl2uH7hRqQF2grpp07JjXe8QlmnFuE0Mne42Tz57jXGGL4oP
a1AWIa2LqeQ7R7LkpHlSpl5OlytvwDpj0WwNxhUO+JAr5qf8iz2zNm5Bofly+Zj0
DtXBfIK3WKxG6sHlJiG+Jtf0wocd7RAm5jPN4+2k+vtEjHMqW9n6KO2zjEjMTByJ
fzpOUSik6iC3jy9TTF2TtepbzTCOcvu/G89IV05Pbt/OZQBPsjnr6RP5Q721vjqs
QEtVJ1IDHkatar/uLKhLKYxFQgsN90Sz1hzaVeX+G2b52obz2m74py/vSTXs2p+M
xkHa7Z8SGDWM4pw1ov7bexfJioQLbgT8e+RNliEtwmmw3ssCwkbzZKWk4CXYfo4/
7HiiOV5s1LI/b2HXUUZWcrDblXkltJq1TSGOMTgcxKsaYyD/Mu6cgovhP/hauEbu
zAcxhyBtDBcEP04Hqpf4+iKnLLfV4sGfWvjGi/uoR2bwdY4/nBEDJ0Te79FtUUaL
OjrSUpApQvW6AdIGZ9cJwu+SxjBe3Io7Cg1TaIinmQMJPZAQrsPoD7h1GuIY4mJ4
DFddvi57QVDGDXz5PvMDm0oSREXFh4cN+03o/5xGhC0UbGJINJqmaiMKr5tG65+y
4EPn9RoLFqueJyGXOulSEkCa88gmfdlrlUayimf95sQWgN3sOxOyR6jOxpmXM66q
3Lpo1GwODlqrsCSVLpOJ8UVkFHAf4yUmM+0+r7AgzUFy8DbfKUnnU4jLR6k6IBWV
yc1hAwgnUhm2Qk/PFlasD17wFJcpzmMij6WcSSn7AkTwXUpBYszSeACejW1WqVHy
GnG82nk6vl3pcMPoeQcbdENTeTClwZvWrTUSSL7IrrLSm+1+X6gX2wJ1GYGs8C4f
jNLseMBfEZIC5U18d+Xh0cZq2p7fXlZTQKmeiPw8kqMJxD+Xlr3FKw2isQh9IPLJ
TMTuzy4Hu1Q3wjA9uk3goOuR0PIL+mfC/qBxQBhd1IF0SpzCXs0dlbRWlrvXPnSs
Bu+GspPfY9bhaDkI3CUQJA9QeVP1LY9TMmgwLXDsVOL/5alecK5ifq/0tMgLxW9b
qbhWXVBOlxWr4RlbYd04aZl0O30+/BjsLM8zB6kHerr128eORrr+wq8CKuhajRL0
6SawaF/YiVBbZYz6qeuhdR7ZFopOCHV5B7hb8RH7SdZAUW5BqyehsZVDMyord2KQ
uvKsPWsePkWQgwm7YzKWcbPzHIAElafheScWGyXQrwydHk/XiA3tlM2QfEeHOuKa
YWtLPjF4xmGYr0pv6gFBWl8AjPpyRgXFb4KQjLVxfBbYQmXkAmpk5VEjZ62v18PA
Hcz+F2cx4+bG4lXse4ZfFijvQdQhw/6Exx2mKYn6iw8H1Rq+2X0+/bGKJWaVZKha
DDNkmqApddZ9NwsfOBrjy5gwmkNGJNE1Uo2ECd5KfeqILxRmCgDcKjJPQ1sQNCyR
dqKixCOuNJnRmhmbhEqOeRzynezVWm07OuiqKHMdmdz7183ks8BuCn6SlfMAbVbt
ZGN7c+MuFh+jN52TAtyYwp0Ag1qNu0rllFSDocJULvLCxzcy6pV3XlCvvkn4xxXg
gKMj/OfdInxK23Llj2+NZIuQD4n1XHdV1KCDmKSFvzC9L0YBYOl8vbZZtRBGWpN4
D6MAiCHX/sZoh1dZ5bO7OfAs3OzzOS2xMOcKhHUpLiYKJyvTxGUL8Ka249+4/RLm
4jLd42hT6aLOqQgI4aCvi0Dx2TuO/ei+QGiua0DrVyykb0lfcDoV40mWo1xaYtNP
swIu4Qk5HxppTxENBuw9pz77mYkbMtfeRJWNqYW6xA2iRq7ZuLdb5ubwyPBJwAi+
xOTAKMpomijpEpxzsqy/tG+PjWwtmxcYoH0Svg0R1ygv5jWbQ4hyXE6mb9u6bHgd
8kd7YlhVSPG3mj/FBmxOCOJBJGbFRmB9U5CBPQg4QqxEZv1ixSo4aiMBRuTBPH+5
YsM2333L02+6M9KkE9mvFDT/O2vN3GJn6b0JMQ0MqnicfA/fUvoLHaaqD5dK/51q
FiHqbbi+422MFm40RQ/NEvLCeRMSKK/hm4+WxqbXPQ00BHPufqyUB7zT0u80yBw6
QdZIFAg4c+bFjI5EWnGpiNya/Gz+uQPk4d7Vhww3CLBvrPqPj42xrWhFpnEAd0Io
iwS/M15jZmbRppLavQ7j+U5WVFHqUNPq2MBQ/5f00spOTdLycyZ8ZNEGv5Of6HyW
PgQlq6bwy9xAHo2NDXdwSWw9RVRz56xlh7ErRhC7/Ebov7lSGasiOu/1hsimxNwX
CHUUK3SYd3xN4W2sKx2Red3mDsJGtcWZNQCX54paxj1x6aFVPdwkCv05CAgWaO63
RqnblZW8YshmiY0O7PIP6RLRey3BQrdRyPLeCVXjgDSQ887trkxm5TZ+Upr30Fj1
5WnPRcdB/pBl1H3jMf+gkN+VCkMngvYhOYkAteH1kFHQon1wnxhxh2UeNf7W9yN4
twwUdbQkS0aNvSp5jd1JZwkVX4jxgRYoXxAj15M4bN0/EuuGycyA2r1DaAz3pNxt
6aG5tJbm54KebYeIRRQd/ucW3llFZsaQMaWBR+FYAxX/AceWaf/qN0bg/hGTgBoq
Hb0nzRJOIO7/k11c7S8TWujviXOPQXiYcHkiwsBAvb3AhMeYmuJCh95k5sMbFDHT
a2YGHe2/L1VDK80QZN12S/AvmMiUdAT7K8dlSeUw5C2b/KiMhp6PAbpMyP3JzlyK
FQ99gbaYtPlbE+KT1DiJ9sduwZtUDEAxB/RygrdueSStU3yYASBGlr+e10OEnsWn
5wWSNMGrnjkniGYKZRRtb5D/trLP0Dqu+bbnTUKbZVkrLKnJQB55blulk+nfSg2h
rw8v/NwbKPy1WSPPy8Ez0PSAFjKBvln4zICQ1uVR5btvIQV1IRoKVuPf3Q79Q457
7mLr9FrGBbb4yeE79rChV84AAQ/dydWjLuhOKMWmRBt0RaiErCRPyuAtJELKFBKY
Cssn/pz/FNb9LlPBEhaQytjLwRcIhhTbgnvCKn/x+wIKfFmIoMJVoe2xwwvElqqi
cYaubhVZ6m+cieP31eBLSAS4aExyq9Toh0x3+zsovdZGUMC7VfmoZNZk3M3/qwi+
JKriJlblFnbR0ch1DoqszT/szOZpHLPxf1cwFNmyrLDKnJkywSJuck47NVA/xDUN
TRExa/Z27PJxqSyMP+dOnzyR4eXMcE+xNaxoHUq4sb1tRyI92NoCVj1Jbn3zOjyF
uMTS5f1nK7nc9zNRvKYJbDGDE6bzL3Y0PtxFCv34s2ZOFdm8FHt3UU6DrKsqSdso
RR92pjKbCpqGs/TpZMwZCLlN37EEkKWAW6DkoYAvIwnKfNX99JWF0izdlymKo3YN
AQMI1pwdw17BPZuFDnu3crMfrVDAHyz8AY7n/dLc9kt506J/u/IotuqaAFslYgyT
NwwSAIuFOYMuO0eBiTOEm7/wrRWHTgG9AdOkFlVgdUaiycgWzd8TqlAYzKUaDasg
E7QlELtvYUkUbdAaGv4MUAFow/FvL7pY6TUZjjo8n8n/8EE87rXvNMNIglSMhSFt
M7edyVOKDXMR5Nko3AamUyPnnp1jPS/lHiNO5KQ3FTI91VY74w96tnqXwpDq3RCU
Bdymlna4yEuUnROA9awZH0/bZKd5iPVSuIIpRsQ2v/YpoFdFK9BiQuOHoa0WtX1c
wc+TFNerTCQ03i0KJFq63jIzmZ88sBITrP6Ee5Vz3Z4rzEZ5C+hlwwJK1j2zafGe
cDhX0UfKPr7pwm6NOvoSfVxdd3aCKp5an+xjH8rzr8CH8+hsYleHZcHe/i/abpPD
GCbCNJSIeLOCJlWrk1/7vu2530w+u8qFn+55z17VZ17ZBTqcHOr2scO/Xmz5Wknu
J0xNdvMxRS/ZtmC4/IChB4+1oUK/BkjIkIDDznvUE/KZoflHFoVnao1Jz8WL+Ox1
juGX/2h7F7rzaiwWHDZEQM/3StbJBaxiKmi9B1Imdw4OHx44uo/G6CCTXcm0L36y
0Xhhvb6uK3xHYFf5yjew7tJ7UB0Ww+dyZOBVvPC9SbbEL3wdwIW1aeUY4KfY0c+P
C3UVs1meInrgz85R2c/xX8A/EsJhTZ9aWNh/Y+ivlnXdXTKK/dCJGNddwWihQjk6
5WGbniS8U6HciE7LJfCB1LH0dxBr1qprs7pC8AKGK/UWA7+nN60sV4kza28yG/Zq
dDqedFgP7e51l4OW32oYTmnT2+Cc2eGAdK26L0DVizfQ66PXcJxYD9cbcztxvFUB
Bb1biVCNY6FZtC1YnYMoukwcX8/QJUWV58zqHdQQaurpwkhLOP7MN2iX/lQXXpDn
eyThBdLqLOSU77qqVR9t0yycWm54yUyRCH+XHMLpf7Me0PDP+LAf1pJLeaL6CMR2
Gg0EUOQmZTxIxjVL+S7H9SzjXlQ71cczGdExbmXkXqGnvQQcVmccTvuC0uCVU3Zu
zUC4dLH8TqEDyoGP5ShxR/jSR6KK0hJkI370ocg5Ls0Xb6SWNKDA1THvNZN1Q7Ng
nWgI5bkb9Kk0b2LEgsfq21va9XCLDBSpzmEbll6BNwT4qQ+D6hRIqWGefWhyogcz
Hcef/7vGbq/fBIfBv3LbYOaDBZNfxke7KGdww8c9DGhjaSJ4WuJWaM3fLb6Jdg9+
NmzJrM4QIVWkKNYsZBhABpxXf7v0CTI+ov6rwnAZEJW1LRqC+nyC61o+0YpSY/lQ
K9DUteN1zWoujmkye6y7EaowSNma6jcCHnxg/hc49fW3DiyVdXnwbeHwBknyCThV
NWu/CQNN4ZEyk67dRbA0duguCggvblPePvu4qc8wkc1kFxIm+hxk4N7aWKCnsDo4
BWNeoHTRm7Z2C7wclOMjruFisRYuPfoHPzax62mPxHKsN7Bikz+2LCgVtH9kS2wu
HERR9ZTc5YKB6cODcmtnf3qLS8TPyRWFoahYJvCcEIdc6NEkD42tiG/5ic9/8Obb
Dl8agWbm1CreqFLUutl9dkMOKmVnwyZytmtxgWHzlSfilybXEjuHJ8O/qUuz1AIo
Vq0YwWcYYnKBiOi9pqLnurk7OKkWivNOEKDoOUiILs8svH8RgPtTanL9CDPxYi+3
PevoJi7gR+n+KHs9an+RltaNXFUUOEvRFrTc0DWe1R+S5PQuvj4Gies19hawJe0z
uEnEYOsRHI76vXzNl0r/TpJBaKuA/SX0DTt+OIF8D7DwlDIAFlr7ym0zAVw00iYr
7ibgu66wuXjmJEoL5sZz4QGsEYxgapFj1kKO+JJ13ezfOFUc91+I6x6aj9XKsnfX
o8TqrBjdRmKoXC/LF34lLECPqYWbq8/mwsoawAP21AES1TByZp6g7Vq9bK5cc0S6
AP2LubdsTPUuu0Z9VHq+la9QZxvCVtHyHrvTnJtFHVIqcL1cJUZfjIuPPXcS9f7t
bodj1helk1YkHHjtHdN2mE6q4YR1Ou43g2HW02nMxSAu+GdHyQpVFGxA+rNbTZej
jJqb9Xrt1IJ582AIvCouY9zPPqqCp34A+UpfKyzUBMzQ7tOC3Egao6KCWvsPf3BS
SedI0wC8vjAksKWk84x7RK70wLQ7e5x+5R+IryFcwtUaOwbKGEEhA0ECxN6k334V
/8qZhoc5Gft4AcuarvlOMLNA/ptoHV2zt/ne8HPI8o14g8Esw+tRZaYmkvEmx9xU
3qVX5oPcQGr+ST6LLsH+POYmyO3gRHLFcfEmh/OQzSZVHUtap/EbxPW2c/opWFiC
ictsTjZXyjRFH9dcqfFY64fcaiWwChWk9YY33QUiq+dD97W+sJVlqmT6zs9oOycV
tJTteOA5YtWvSYPLqBKAngw9hmsILE+NSJW6dWng8M1fdfY+sJqtoJ5X/P7mIuC/
SEsWkKQOX9OcDZLB/LAW6Q4PjeWCPY/DUKEuS39qi8HMIrwGLngNLHCVM8fh8pva
PM27d9ZXKRgZ+s1zOivg1d2jaIAZPzJsMw03f34uybrsbqQNyiVzgTq+SLtj7Ws3
5QudXsG+F99fMBIYeuzJLAQYlnGDHls3V8yORNkagx9vD26lmLdn6ZlzeZr/nFz4
+/zPwf7XF/Z8aUqaj0bve6+rQoncn0w4QtDr10WoApAVcZrQPWABpeqq/WzYcA2r
P66s+3vitZjAOxwh6I4T60amuLhs4lPbPhq6YX7Cr267Vv3e7qM4SNy36RxCXWtO
/bUy8rXVPYeZHdeY5hkGleqf1PWE5bZ7TN/2KPNLsT8gapzv5S6o6+kN7sYsg1CQ
H5iimPHHP7vv/YUcfSvDnkTltDYP5OexKEtZrWzfQtXyi37ha90olMBo1qmN6Z4/
FSYew2LyYsXsCdMBuXhkLjv1uSHt9FrPfwYhTAsddPD1LtFgveT7pycA38Ocq6lL
k1c82LtrblANygfdsAQbPaietJXViO0yZrQFM6gjLoGu1U09v9V0K05L0XQQlkB7
GA9Ikrk2K6CZMdqC44Cp9PbHc/Usf9VaBnDIr0b0Qby5A+9bbRvNy2iqcbm8TY0O
LRnxaO2HL6dXQbkhRus90fwSPrguw+bKrJWi5stI1bk3z3vl9CyNSk5xQd6vr5Tk
bZwXarf/wOMl3de9MdN1b4IduacVPC4zEUDWnIjoKaCujXkmQBtZD/ZkaxgfVGU4
Mswxmwl9uliF8eIplYY75JhCjPp45xr3JT9sC3k7LEejKAURIaed1imhtSHTIA40
RsdgSCDRMppqeFC5R5xNuy0n6KkhUJa3nmJkL2Wyn6kV32hlOMvNCaucvNbv5JvK
sINOFdWmuSRi1r32OCNU9iBFGowjfKvk7uyLSHavDw/SmvuO3gM/VXCjBhRj0UTi
OAHgfeQ+MPZGFIQpFAVxvMwJGm0QhfvXq1FEmmUw2mbih2fjktDm9THHjFWk85PU
BIq7EsfuL+JiNzeFhsuVnGt6HvJLQhPvRgUVIwIQr+Sf/wQuHwTCNO7e4XBdvkqo
g1Wb0h1MuvGr8/gRQqNm/hN52mvcKN5sNJJvegqe8ZbOUlaXrMMuySDcbqEb1QwR
Z1ntMjkfzVSjC+TbQDdO3FNHi5TXKY9bMK4x7RpuJ3luyTb0NdCK7RSjsbtk5L4r
yQf2mnYCQTDw5ag43+AZXpa85joVO1eJIH3OzsothEsxAT/+wcWwUHG3sU/sEFtu
sm+Bb9epNCAXT1cCn5K1ET9h9U5/XApGknJ5yfBhW7j5hUmAEIlo1uO0TyeyyVbG
qkC+Fr6DBpFQXgn9Khxa1pPMYIh9xJFLs0WnHv1FBTPIYBiRtxxeeQ/MYnCQ8rzH
99RkAjnJzijvI+cpxTLJ8GJwU1/RNVGAitrADisFca7pWT1wKbGkSPK1LhttO8/N
yUoOjkv8aTiUAYRCjt8Ui5VmhL4NItc2UCQ06XAilbMVXkGaX8kfFovPAmVVhlu8
cv628a/Ah2OVrWI/9OJTXJpHMcz7vNMq2hCT1qTkXqbhe58gneLAKEHqe4OCQj7v
rKc27LT4Ii/2q3vBRTBXS2W4q2SikvfTss/vhGTW3F5ifc+NnHVQLqqxYoKwnQQ0
tfLitO8/qSMSpyhQU5czM2GiE5Nfn+LD6V3t/hntLu44t2uJeKbQB1TXPnY9hm/Q
iW8iRAJuvtOJaZkuMNVnkEpXCksUsdwuiLJRVINmSeUOq88xztQ8Fe8JSTBrtOha
W1k/8GgrXHUL5Jx6ATlfBZjaL3+pRLdYwfbKAO9xZG38wb9j7tIKzMhtBntEpSM1
H3zzqJI9eVqLn0sYx4WruCL95Tqbh2+JXSjukBmJEKSHzTi8htEGTc6GF0ePryOB
SxJ670/viqHd7mzY2pB8KiU3YXBZuhmAyMF+2nBlA4iM4RmPtrUmT8IBEVVkmb4O
qABUFf5gNQHoDuOLZ64ELefiXjiXPhgGc841XC6WOuvy/7ovLSZCMjqE1yasw+V3
11qK0cRFmk/VeER75xZONjByAoTklhEdimUuCJNnX5IfuHOHfLIEPVsijdDxYk59
MJaF1WqTkyyLZiVee2s0ZD/D0G65GPmwPwmGPSbZeY4Zq4R+Z+rnitlSvHgRnGY2
PNPUqvESCCe+QkbltujQeDYAXD9sZ8UqNjDoea+Y1nG0lwv+tP8NFk4E5uP6kTAo
04d0wLqvM482Da5FBGE+wXuumCclHQPO4BjAkhBha2HA51xjqFquBPhSzIKAb4nn
9a7rJu2MyiebC8KO+WMcwWOL1d7zLTOaP+GtSKA87w4GgAYEuXuyHe6dDjH32diQ
+sc4TW+8z8KC1iBDuLx2AoxzUF77QjyzZiJNPVbBOureCBS7FcXFAD1xkEY5So2R
FCYj/AxGZ6kDMZvbjfEOGJlVja3sx9vNw+H7/DmQ8SW0+rICsyDlUY0QsCApbMZ1
LsSbXzFxYyE+p1zuqs9AO4+ZYWSnAFB4apjamIIsPMaIxt5NA3v20LkO/0PbYKqK
yywir67wWLoYWGxX6FoHzzzX5qqtrXfcbHBmqgQ274ctKUK9wmmICeS+3uBYsAFu
o8SSOSFFLQQRJhhccynnSCzm1aBpdejhbGFXWnSCOlvFvOuKzbJn/QVORdkBtR5l
8Jxy1zsruvk5qmaSIlg04FBu1GCR4QxI/YwzlX/1kLVTfyHkJqRBQ0HT2J+Nne37
f1iI6hEaqe3JqtstPuxJqmw+QEfmXDxunDCX/OE8TDLbxohMknVSsIx2M9rGx3E8
LbXD6/Xs14GEUHHoj1hPUmI/9C5KLyQjj+AK2R80MyjIVQKiXxVZZHjIKHyJ/5xc
9UVQoY7rK3jI27kex+YNuwsJEC/iM3REb+rNQ/PLdZpBZdd+S5/tqbSlKXGAXTVx
eNF4nPZxlsuHnqmbfR+6o8zmV7Cw9cDrvYRx6JDJBpxX+XNjLjp0v/tt9TMFTqbN
vTnmHVLhim08VyBSu0mwc1j+/ecW6bN/tSzkB8wUaVqDmEg+Z5LYyglbgxOCBAfV
gp/7UDgtLh7G2d9gBo6zDmx+k35ndUaEZOZdyGplVjvTxDUYJNHYGQbkjB9YIHlx
o83Pn+RNobs63uyap0/Vz/ZNdoC51EXnpF8joSV3+7Sf9rLg56GPBvywOBYaCtaK
IiA8hlxuUbyQG4Gekg/2nr/8GN+iX7Lxym4qM3P8Y6JKn8n5gOzrgedWinIRdn5P
QHv9J0yrwLlqT8PnYmwx9c+rcr4GjM1e5AX6mGE9ZksvCDBXb/gSgwaco9lPoM+u
Fik8t9hpUuqs2TuJsJWrHQOVz1Ljq0R2is686CkP3lm0RhhoNjLooS4mi25/c7e4
/3gnjReiCgfcCc+8aLSnT6GG6++Q59c9rusfFiiOrbOqhsEhV9j9i714kotPKWe5
PHvhBDfIHE8XxjgqkGCx+uT0nRvyAwlhDzmxuzB2iyJnGqeZHhIu0VVsqhAjsgMR
53rJ/kDq4XpKGuMueRptrpbkjb+m69Td85CtMEBe0zTiO0i23W9to3SiZp4wYJQY
qJ3ftMA69vn18XlIK1alqi7K6JR7FdV32xQBnDXaEid9tnD7pRzHc7NptUYQivSO
+8wgHcwYK/y9jiYxSbKXgKd5yU/DF9YeM/THuVMiPW+086olzVaMH6JYzXBaI9Ng
tOhI97FA6CoVLTEh9Lk5l38adXBPtlPU9BIjcMxP8uoWLOipfqyMnFOQ1U3NuceB
eVUxQGFcBxxUqjEGdKcYKEydmJozS7Vos2xPbpUMHm8msLENmVWZExFYrjVh5Ffl
C6ozWc4njLxKrxwQMSXlSGSxGSOsaXI7dVWvssanYLoZ099tmAELGFgbd9tm8Ls3
kqxr+67ZVdOnXmBnEXAkcfDN1gVFl4okFZJwf1dv/t/Tt8yRhQf5heQEjfjx6FrT
xD5fZJxAbp6yyMeQSlGNjzh5qianK0uIuyYs04QIiDVaMbiKCkNk9hqXBTBhNEVG
ZnmtxB+1xggF3q9GC/HvAS5/T9Flvw9N4MVZNh4gjKQWa4edxH6v36vjlnAuyLg5
wzZVxibUgWXUm5CnJ9fldEKmJdxzlamdIn4An7CgPc4QuDMIdB3+YSvZyokVm298
/ZCe5o68kX9VTOlxgfq43y/4cEplZ3VvxMT9OVNPpyCPye77SUe2zm6OkdrrXouf
hvi4oy4JsgLaT614pW+fypFC0aEgmdmYSL+qqMglrnf3s9v/IIUQd8qsI4LMAN9B
w64qVkuBdDgxh545a3eb1W/oAOza5whHFDXk09rpqPwkzjIfevbnd6nO2uc0bvob
Yx+L+OmURNWTLxV6H8b3UFi38gxg4Vmabxbw1xgb6mrO8HbaJYvCqih1E2Hx5cW/
Q9U2Wha9CHwPLah40UOwzsqssLOOKL92hcOIE7cN84mUQUi0TCXGPyOpZk9fKljC
6q1zJNGL2Pr49rduBrCcvtb1NM1mFTFx+ugmSbuLsUNYcqczZ/kZyrsHgC52F1EX
XIvDUnZq0AvTHyPQIyLh2yZpna8b57k6iBoC0XBNJpvkPt1/bb3c50u+Yaa6YCwu
BZBEtISfcYuAjTWW0AV//zH1ser13k5irAk3Y3Junimv1wdcU1guTfZwbVIFTRBg
34KgQEOZ/7kJCDu2xr8I829RpHhMQY8iWCrdW8NsDJjwJMVXJOA19b3xGdRQk/mk
UbXyF01k6AHKPUZxNGDnJB3e5Jf0Wovwzz6kIX4tRdaTLhwOhHHT/fnq0xmfo69+
yZXJyO1BI64o4cC072zHaOZLdNkQP49j/dfP9Llgasudq5GXj5isx1PUirnl1nBs
JtwwUE1xooOzZa/hzb2006aLv8BIW7/O05zsk0KZQUi7y9ZIw5iXLL5DxAOEg30D
a7TRc9AzGcpvlg6m16TNugoSmqDjVyMjFhLWuSzXD9CarEmx1PyjeRQ/OxdDl8fM
abcAsFV88Au7O3xN37CbuSK+syj2rYSwJ5DFID2l8ZXocBHuc8jUR26Vbn+BI51s
GYT6iRoTH+vxPFTrjBSXyfhpOjQDXL+oUkNZ8UyGTy9ihBIVQnZPwWGMVcavFEN+
/tFk/q0JPW9VgS/NnkWPsHTIh0F6xzKrbQW0d6E2iiOOOINFprc1X1mQmNmHtn0H
GhCUMC0GibnPRLj4SJVpK1SCUqjslYeVjOvz+NAevql+SGhqm8TlKeSMIIN+X+8H
T5b95nmdEnMrZScHFt7216WxUOtMwvhcaufcoCYdqfR/qtbIyGe9DzcAVWqulYjF
/6P/JYpnZr4BDapEfucLLxKxsqyaQ3+vdHYYAH97Aq/twve9zhsYctxzgp8hDDI9
KDwdeAmYaT9dUA2Klo1jzT5MjOVmCh+JWHHIJ4KJbolMlTln/VNf1kky6ZKS+aLU
wIsxm3SRGWIKb2Q97f1mD3ToWea3db8lftx/M6rV+D6MATlTWCTfm63WFU3h79k4
4Lmgx7cJPQz8w6fsYsGjj33dDqDavh4/yf1ABAwVJONTcZmwUdzoNQ1SxwcCnios
fsotJ40GpF2T7j3UnrUQtTvk4sBbZV6pTtne6u33sqvFLv/Weza6PZRgPCw36xC3
7Ynwy3i8sjuPmSfDk5/D+9KZJy0n0s73n+iVDDjToQ7GGVsfmNDOmdwpmWydAvir
me9/gFfV+z1MyLbdChKM7OKep6wy2KZXlajxlRL80vYt9NMI+7eQXFH4pshSY+jB
EEnbWsGRca9BtIs7mevivG9wm2wvgZR9d7Gipb3FxqycVl7i9D/s57gOlbNhLsiI
ZR1LHVPGaef6Oi0EKtrXwiwtGogSFpnGofGjxncp8AAHebaCXL1nucPdGlBDy9Ya
bLIyuSBl0iKBXTqQVj9yFiO6afCpPeZEDL9bzA+nAPkeK+yAjaJ/Tj0t94LobVLY
yIG4cD/Do8m1tt3+l61rVL2NWbJ5q4mSr5MQBCyPUEvUNZZ4THOBPPi0UbvyszOg
UW57/1rNM+3GMu30Hl/wP5h4hdt/8bt/IuhZ2sputyBzTp8e/Kry2HOdzaZus85p
V8On5v2RuvzSI+MgFBh2oM2RFEmYT04F/DrP+QnsGlRKsp1PrQXDAznsDWCQ3zMO
TmBHFTdfs1GWQW0JfWBj9TbfLWMAcsgBgSgcVi4Ry4rZtwrjCPEeKxgfCuAB8Ndz
DEAjoWvKRxzxtepwl56Se28oHi7wLZRfzy0FbdhyK6rjIYgI5c8pWZ+40A4Y3TEi
1dElXOmiJcONMOisAsQmtoyW53ZTrCaW52oinR+MimqDWtLg+B9YehNBVqYFbNyY
TUwEPl5Yn6TF8l6PjBTyVLax38sp3m8LWJArEouPwYRHNxtnGp7I3mxQSKT3K8dT
BnSHLu+T7x8YVk06HWJu3NXMWJRCeUA1aBaF2zADzdkakNeNRcL0f10U8oJpCuz1
qJ2TIrUKoeEuNkxqHsCQ30XV4UOp4ZLkcKsUMhWIcSBQMz9Mg6YiUmLIMNDb0Fex
F9erGvfh/WorhvGtXh7EIXOFhJwVSPMIJ2JlxFaKYVVwBu6DcOtGRvtR3qdA1izA
gSzRLXyVSIJDFYpIb6TeAGzFvIt7l5fB/8CFN1WFzyDlCUwYB7h4AD+wFrHET4JR
XYjVplNzN6+vdYPjkBu05e9ex4DiGLZgmyY5dYaBXxn7xd7dWisvpZYpRmkHY+KV
LDM+cV8G12QkvRHBBqKnrQgUHT2RnoLt5H9uyji0M2iZAmOvYkeOG8z4rlYed1do
YKGUvnliFfJd0vErSGYTREf3WtDpU5M36HTWFpc85CZtLsgIyBwaBF0rFznm2xhm
xra5IWHbW5RtJpDbr3tEMG8ZtvSqzJ3cpki3JZbe1wd7OxWr0gvse5UIvXB6r8Vb
YflFlpL226xiSj3I8N0ZUacmmUU5j2wEIvYh1ez98kOiO9CdFMI6FIrnPSZifJbi
pScgkruOpKhjoXXowr2hgbrIBpgIXGrgtjXQVGah4jgsLWcEGHviYR8xj6Kv45NE
DJ1A684ewzJi8UHwG8v1GaioH8t3avgEp+PCGD/iol4wkGz5CrmM+n48fX7Ku1rw
9sXsIUAM94UBzRLsNxzFjSxo9r7ilg1V/ruHRRFNB0MXu6n/oRqtv8HvshnFzL+W
9yNYjs8//SASguzoQ1xuaMbHQc/huxe5IcBI+sH1BWCkMb7LqKFxVH4a9TqkAUtY
/mfGfaeBWevOR+W7RE295ALq8b3uRd8HZUfnZEbKR28OPbh0origTE7BgildhyP2
K5wnxw23Abo+OVI3fXjMTjfUD9vuR0SobjhcLiVi4yHeTPsUJsS7fsmFWLD/XEFw
dw6wSVuIuMsZanZgPnYGabiHIjxzXbYSqSzHxnAQegV8RcqLfVDzpZOcaKIQyHJV
TOBQBhQuqeiYXLHQZusddDR1G4T5jUoItVbMplIztCp2gTFWb5yGAryowLPQU5GM
rvHIzt7DFTGiz4N92KP4r64UjNNQiurmLhEEhJl3995/jX/8D5pK+F35Zt2icnj8
6kLzqm7Tbhi22lWrJYGULExIx4YXF5SgpJGvENS4JLq4VQomdwo94krOMteNPh2y
wwDpCChwhd3B1b0kLez+n/qrnyI6HpsVQfV6TLgBrHXysdQmKR6WPfHdaqZNRWJx
BSi46gB8lZeYRH6eEoHI1X6Kwbg1Fca+chzRsNR6h0pk1NDs1AGDcRqPODjf6Tks
sCi3Thrxk47XNZ82Qt5JjD4lC7NhtkIYr7QdQVACxxH/6PW+uhjBR7bUrMejSlt7
3QQOsgxen+GNg/anOIT7M1SURkLi0F4iF2xBL6yZ/dwaF4V1ygD1QILrTuPHGF/a
qpdu2rrXTVcvvtQp/Grr9YebMFU6zKARYE0//H24AkFjKl+3exUc3L451KMhq9ON
tbnMTKoGYuGLE9l0Dg72k3KHGTzAEiXx1/Bp+lxxUh52MGSMzvU/L/FDn017+eCP
5vwJeCev1iBl/vzohsTxI7t6MbOBtAuOTR2//ZmnYp+MDk0lUxAH6DVu+K1/CeG1
nZ2GB9EB/Axt8gfTjm8946vR1ahw4rCZKpcvPgQoWlzqN5IZ7bfKzNMgMniIMy1j
QXDayn4voZoCwKO4j1rZRI0VijhnsZ7FluzGgomA81Svg3lOO5OvKBtW9hVB3A4w
xVVKXwwonm0gX9Fs1gnAoH9oERyAhXhYmU4NKt6Ngvw/5+umz1R8q2wzGsJFktJa
++dIJyZDtfxqhTb5xA/qv0K6qOvapOj0yRW/ZqDhW+VNloZUVfDrwHX6gwK1opuf
Sscmrd6o3oFFa4XD/jSqVIExLQobX0q6wnuRCHvt0YXa8ufPssqsKS/A9oMbpiJn
Twavtoes2PfDktSCCM+EfYDgJbVo9ZgNRDAnq0pFHoBqQuqHy9S4xpTa9y7VJIuF
9N8BYZDp4a32Oh3NkDdBrRkP92l/oDQAPOYAnNkCZhwOiOBKUfIZHWt8nkh9jzvp
5lIrDxXU7596+7w6FUqdHONZWyWiStxPiB2K9vp6PzMgiZ88XInIpvYa16fE0VQi
3rob3XsAiBrSNLuncdTB7zL/8p9lLslHSjMMpv2DVkexDltXHCQf/pZ2yxHE1xY8
bnQ1Xl/bV5z24XWzJp4AUI1TT8R6LnLQN7c+/g1cVT1Wm+HQxGHRGNNnOCVTRN4T
ON1aK821icmIMPY8mqZ+Jj0UM+8ocsOJPW692ikclX6IpwOHVeEFcKQfMuTXzcdh
RHTcSMCWIKrSZdBx0tpUeojX56CGcVdjWyJe+e6aWhCXEzKQ3ti+b9qX1+hajlHk
EE8qCLy/KlDeaOlVhTPzhR84aIdJGhLEB4dJuOqmHUtkIUzh06sV+lbMlZ4Xmmnh
QeIasCrV5iNcMEI/6Mjo8sBQ9fq+wycG8HAwWWSN11amQ2qVwSssIVK6IfAdJwRM
vr5jx3f2BZuStTh0vV28b91+M4dJNS3CtN1qITSoHqnThpxngIKbpIxM9wyWFKpX
n+uWS3Cl/MLQw1GW+Rdw0i0wx73oleqwAqM4+doIykAMgLAIclxvq/ahbkn00Ku2
XxlwPIw87Fd5+5FxvH7S5m2TiBvvuaW/M7g3J2cV7BF4VIkD8Cs1jWrb+ydOOsZD
SG0vgux8u3yInUj4//Pncpkr73u08/JT24YLKXscP7SDMkBm/byVzPmTjWvH5yan
uvb6BKDoB3mEIeBPYEXb3mbkutuPAKHehg2S3O+pruTUv4465zgWn0EPbrruJtsm
DogBCuuFrSKlUdbFu5NvRXILluILnbkaD7WLm1T+b37N9TWzPwN8MxEDyL+VhocE
g1ajrJ4OkEErWjMuoE1T53k1NSvtH6fMgz+3z4NzXiRz8cdg4J2cjx5TFGVR5Ftu
faBNakN8xS9JJSM+1TG92/+3V7YWVvYfE6p4gDOkGvym0XL6/wpKZYtN/6EzMoCq
1pHT/l2alcod84v8XWtVM9iQAnt/+cqLggpfIy+AixkSfskNpiXm/kedMlIC6u1A
57NVEHQstc6PTh+WeU0pviGbkJ82NoaHaSPxZAlGFnNl7PLLOeDocQ79Zl9oLq9R
wuLDb9R7hv4tcgFHjxOP5x9oyuUaYGH4XrJZf3KprNvHxLBMaSDWTU1jkCtxN7yR
FgkV+3JFydmdkaB5demC3PJzUc2p9Q+I2aK7LfPe2fDa0CwI6SWXtLyDIKbYr9HB
WnZNOnKtckvEePrR2b6yCbooYEBiCsbsX33bCrHXyIxM7HGpJQsHa2Xsh1U19FeO
CJdcGXhYYFF7ay3e8um4zma2DeV8NM01zs5svv9EgQe8jO0brjZICIRdcItZOfpV
UnAwnSklAzkNVozWN/ZN49eXnxZN9rzQPomb6x0170p4QJlkA3VaPTBxtQL4xeBi
O1CA1c3ajCH78bV9PlgpesP+VHL3m9L8M6hqmwQvkecaFpDa4F0wofqz559Pot8i
5DwJsEOD/X/wv0jONr0VbWp7sVTtAJw4bsl6CV+OOxv7S9NNxbpLtzDlH/FB5a4x
nM9KvSdja/Xw5IDnIDBQDwf1/+j1hhP022+wIDJcKYKz2JqJXGlxutaz2A/zElWX
A6NiVzswLGMaxLMBBT2tLok4FLN1Mf7PMCf4M1jb/D++MD2QLdwhS8v1RWMp00hx
CO9H9Xm2W5qwAmviW8sXn4WEzOabL/xiI7/Zg6cKJ++EQi7laWP8BDH/wjzThCet
d/u4k2+stzaAsVPZ4VukrlQtKBPHhvH0MP09op7Y/91WzjlqguQFZ7atixNWxOry
/pMUKNKoin5scLnDnY6yWpEdz0SmpM4S//ymBiTS/75pc6RwZZjz4+oBOKGwecAK
QTM/SK68yznbmd76O8q6cvebNwMSBXjLHTb5PTFb+YhdfZgABAwmhjoM0E2hxgnW
r2nyH8cmRG1IRxCMOL7gMUYjN9vJk98GRD/upVGSwM8lP+dvtrBJBk2ViENIY+js
J5bALAR0Q2BboVIczdy6FBD1b1I+9JQ8hL8xtWO0BFMdv8Ly3+p3sPT+DrqllHo2
cD+rRGRbTQ1figTBa1mAt89p8XjRBeXUFI5gOAlPicS7iJ3Ay3YAVoNhgEA0ICp4
E/r79IINagrLfc4QDRUK+J79DVaGXGbPMuZfLOUx8GLMnGrGI7Pr2Ep5ypOvbgui
CJR7zsLwEesA7T1/dXzN9Ueej11WHQuBlSPYJubEWOzrjqpRVz3QM486ukfHfqsw
7Zd0yKFKu1kFrPvU0Tfy8QiH8dTp/8AnISFv3SsUeLgknZNgfUwCZKY17FhejhhT
U5KODg8LYRc9vAwFBYd2TW7D8Zn0lfU5pV4JUT0eZTt46UNbxStsiBFEiWZym79H
cCJd2ypasFJGeqvAlqZ6m7XMXjIRK2jhS8LsApG9ipOJrPIdmbYv15U+dqVRtnMD
AP/USVbaqQg1lJ7efjPD9uzPpj1sUhIus5Vb9P2zur2BKfmCvRDtz8mwQsLYR1bd
pXzhUJkav8ltGDYtsAzuCz4fX6u/tmgKa6fnqzTESZV0X+Xr0l+nnSVSTz9svl7f
j2Iq8YIFGainE/PlWiIDgd3e8CIqKNbq34ZusLrO3ivePMAtrj72e5t+88JRW900
OqDSTfT0PvTT0T03nvaGclcwI9r6QN5bAWoim+m4qINZguKoNqki3YbSeItq0vjJ
wIfClVoWuClCSNo5gacCNAkdbKJPkH4FKI0TQLzaSX42DpzPYCLYYNGkhiUi4QCk
w36otLq2I1La4tDRM3vUk1WsZKzqiVsINtu8kVydBoGCeDQVBtH49WswG9e1T3jY
qKAl+oQGFtMErR4n6FaK4nfgiktjUIQfrgCKhiUmQedHGAqEuiY2xjtOAxPdnLyi
NUA9XTq0+rmgJbujb+XsKyw8nKAWCAt3Q2w5cEOiwD6bcvo750DUMbYsKgIT2NyT
NYM/Xl4Pi1bAjFydTr4YVYiSeiXQLwbzxIkih0xi4Ex+E+YwSL+VJhzv8mVa7CQ+
4MwIZxSpmouMPHLSZu6oHaPwFP505OZ2oRIInyfTweHxXlxlrc2+UdmQVytu3zdR
pVMICRMz0bL6TinY82QYEFzC00ENBhEmfNS5N+mjjcHsXF7CvyrTRSouMMwK2pjP
qCqQUY3Gn9WhHwjQj7VXEu7vjw3OxIXZsJqanbdDlfxXEA/HeF7w7xsGrCFmgKZW
fAoiVZPU/mw6YognplrxWeT8c7al4Z+lE7nOxWa9aIX8xAgyS6lRWnzFn6hYS5Fq
ZjjETYmPXKTXI4FSQCjbczD8RXJUB+j5ZnbNU56MZ1Raarets5fZ1hA3AjE/2uwa
5mpknmO+kvYuyiTGlhaiSWH5VnvX7SpjSwxQLQoffBuf9NNjjQuzxbIfA/yS9Azu
WontoqFcaFuVyxSOY0lIgi8xhHba7XhfmshafdnhRfTseA/FNezvhIdRjtXRJg78
yzptE+f1kl4npqnbRmg/s6oSh8uWO+vW+jz7O9d0+WDm4G6zUqRKVTgrAQpQQ1FM
jKwcqv5C9+yfH0XO6vz01ZJdCaPM1IkpH2SF46Z/XMlQ/xSSDSq4aVQIqrF1aQeC
vbwPhxtRI4h4QUx8ybArTtaHseo+OiRFovNYMJGjaMQDUMsbKjC2Uk6hwjQ8mCub
BeCW5rBRnhmsEjNGp0wR65PkTx+VsfluufZQXv3sByt1Tz1dftoyT5jOmRnjNG2G
j+EeIocmUAgAqhYykRCPq/beiZX2wywHwX13sjwFibT1nWqOGFkUhYwT73m+kKVG
kjkrWpcZTBRncWa+xYHZHzWUQNNwUcCVlLySSg69GOZoot3rScAyaOTivr0tzj2A
DB43J4J4e65wWH0uj0OVP0Vu4NQdSHT/4OkIHwnsXSMfc29m4haW82Tchrbq49LU
0GKphECGFhbNR9TKBPR6AWmPYXGszGTv5rYupKKJPug5aggWXTfFE9RkKU8eDSWn
HPOoktMBfaHdTpj6CEpIOp81n2vfJlO51+7zzlmYBzUGmpHJ71AoOp5w4con6WUL
Fka6hd+6Iwezc0LAoLrFMXVuPI708TmI3sKQSp0WhWc5QP4wOpsf+5Wt797FcR69
C+DTUbOWwBnLw9dUJNDaefsiaQUGEVZlZta4XC5BATee3Xj1fqdIzeKdsueqYeZO
57MZqEhm99FPkC2StdLYw2ZI/NXj2PWZnNwbUECWV54+g601L5gf+0q6xzHxZ5i8
B++FNvMFrmQSIijK8rdpaBV/NXD0HodO4vLJ1eVu/pZVsrNW32lgPyZY4JZWBtph
rR906FNa16oxIhLVia2zzsJogKyLzGdXWj4/zubg0TrqwqHze2X7wRjmJmEYqYkB
F+JepWyTSOEtXUqiW4Ocr9gjJeEExIu2iYMGYcZhuLR0/98BpmC13UFEQ57jAdKz
yh+312IGH4/uuwUAp0M3ux+radkkbWhKxm2kuLi0UV4x3XIoomXohM2L+G1tHBNV
aTwE5013AHpBsGucTFb9GV3ynRt2cdbEUFN7CMD6c4KEyn6PJmHIOKnnmB38yShf
+hCnGBkNkrOLWKy/5WOeaqcerG0fRkQjXG13q7E1xP1Z3mq2xc0c/i1lrCPsUhop
3tV746ZXMmiSV4g+7qyMT9k41jm4dGOV8d3ymaeNqONBH/ZBuMAVknWc4zNcGhED
BTwKXoyuISP7Dow7NQytWgZPGL05nb3YeNcq+g0UCq47BN7v/UxHDctv5/xM/K3v
CsHfNmZygT77ESsrHdF+O3vLV9zLw8GpKiHj5uzUzPM4R+57SYn19iFWIuKamfvJ
jzu+1fnDh1vF/ZGM0uYPUyEsGi+K6mjoZdGeCIoVV8rCu9RXt9x7u0bWDudFLR6k
8kXmPHRfJvr+MhHZbweZOxk1se7CoPdfYb4p6RhRYij0rUCaq4wWCMZcsOhxdS6l
6mpAnqja1DuD2TvVR5S8GgB9L/gkjmAtm2NGkbTol9HrkjEh5k6QEZtvJb50GEMV
UbH8JVU5wXmRqc9TATqby2WFJXTq+k+8KC/5fhuzX+yuNlueNm4hivxvY69k8zye
kxBvBcHVT1nr1dHI9aaCWRtvCmm6YwhVk2y1XyUzR+2bxdfzzLB36+9bGWYJNF1Z
YaWWan0ElVzAFW+vTA9fWoqxMnm811EWJbqb5Q0m9E5eGpcr6lRhQn79NtGG2vAo
bzumXJ3hexPQQB1G/mvCkHV2IOi8NgUkSCC+3x/omn8HMsE2vrhg+NUTJb0w/TA1
76YJnDDInQo+WZ4p57VNbLYERh4LVn43F3hyQZJPERJueWfm0OX9dxNMlOvct6UW
cQqhuht/puI8xSfs8i5vPD39N61ZBw17nwnv/mi4gW4JR4qYACfDZrhTVmJbUgNR
gXlQoF0pihSKm3ezxC/oyL4xStleT9vhn1X/89iYDtatEemaF7x3IWuueD5tkZIX
CDVdY0yZFlY3Y+kjetjwqORpOEQZjFArLFwnBdpeTSs+yR9fvK7lvD96fP/cAfh/
t8Ktpqa97dsqjyeVyZNY+d8+g6FA1m0qO+wMGw9uWyKxuTzXpuYA5ghhKu1J/6c2
3vujnm34YpSWVG6jYIfE9xBG0cmMTmakptY6G0Znp+VMfkbxTHxZroPYcW9mbkkz
/o5tOA6o8jXPyBu/+Zzv9YJVQgUe7wYPuILtQsitu9lvMb0/HHbzmN+tD/48mP+n
Dt3cC2Sc8R0ztkZuKaPWHpHM9wbrjS83pGw348cZbMt2j2Jl6q5jmT9iNfJVudMQ
bsVlkucugnr1KaPihGXZXQjV50oIH1Omb0dix8fgiHP0z7969OWdWTFf2DFIScb2
WoGjaWvGOQOe3MRIhSe6qLBsvq3bXgtBOvYXhQ6PVGxszRhMNSHptudJw8i30WSW
NdZ0+XWGj90jsisekKa9Q0YmPls4Xi5zUSfVK6MjDtpqU9yForNVDGl8GUtQ24sM
keozdMpcneXx+G2N4Uh+z/M8t6mmKbd3Zc4GicOjg1rRVDEms2b+m/mkxJXeiv9Y
cK/qnjXy426pp6twPQlJz2tEpcClkhiTqzuJq3wrtu8iGm5fO2ZeV2O+OECRTq5L
fGoMesQYSiGEacgTzS4SH+Svfs6TeDVPfN9bMj+1BUHIE8ZPGYsSOxAuNbKOrBdZ
skwQYX8sriVxfT+Ln/Qkd+Ev//i97mGVbovyK3oWNZuFtFTVP0OI9xCMfxLkhpUC
FqJnKbKhe4Afhva0f0DYAo50ZLVFHuz8TKMFqKEb+a/8z48oh+07KywwjomNgqHQ
h4ATijJVb5qW9/rZ6DgSn6gAoMGOq7mLH2+BwVfsqgFbsqgoV5/L/EW7EkP8nqVh
FxvOawYADED+wt2rbOtOW25C8wOLxos5ElWZ90ckZXYQVj+LWhYry3ywROwa1HIa
GyHr0XVi4ZPL8GcyzNh6Ldr1sEL36OiHH9MjP2SRG6ig2zRwelpdX38pZzJSAprX
cfVDta9QwztoyH6KrI/upiK2v93GqdghsBa+3Auq5IvpInvaCQFZ+45GGvdqBMed
AAxsVIHymYON3mT2xUHSYpfYOArI46iEx9RXAnWV6snlcaX7BW3Qi67vM+kVMxUp
JGnFB85ACGvrBcc4lIFNKT4X5j6NcndtQmMPgvGOfnzye+F5P2iJ9moFKQ9yCn1Z
v9maTvm9aJJiGXru+yKH9zU80Bs5cDmaa+xaFPZroDrUiGsFIwdwLRfcJe+s/+C3
JsAWYZwA3G8zQgT16Sv/ryoI5grQj0ZrOySbwN9ZQc5g9g+CexmDNULosuXicIF2
nJDxZKMMg4bcoZ/92ltvJUouAPKj0pZa6wajhSoOSvFTzlEYavl/f9Z6NnIsbAeX
Dug07NBsUQbwDqE7cXs6JBkyCS0W+L3SaFRr8bxG6P6r84DUwDaGheLPdpoH3ty9
cJvpGLjFCDCZ61anKhw4xFg810FblAmsQXKANUmxGQrsxV5/UediqygjHbSG8uwu
wHzkxeaRqWruLzkk/5CkuM/m6a9URXYmcr/KdQZ96dTxmoyvo5Yw1IyJofOuqw8b
18NZd98/ps2UvAm0iNAW/ZkgI1BaT55biHkZakB8NuzzeDWyDR7XjdHhbJe2knTK
mO/kpvznhrwUI4LJ+YKQWQB44AhEs9uUINbgd3i2nS77Ri59ggXkcirBPtZ9uVJ8
yvumN1ifkmT8NkLaorW38UtBS+jOcRA7GPKqwf7qkWxhsSZQXgv90wWduRjCrop4
qvMkmVs3HkZw4UxikhqzNT/3AaPeY7qVDuKw0Jhw75n5jF7qs8ROuOAo+yDA5nPj
f7LUfWf7KGr2ACc0nwcYhXsSNmW5a3so0FKZdDIZ1ziykudDUSJ/EavHHlBLwSbw
DsaPJC0iB6gvakIvvFPdc2FN7kU+PcZomnHWrYbBYjn/nAIybPEyCPhwp6PSYLQ5
PgiOBuucPMLx6XCuaPRHjCCYH+TfqPaA7mEk0woMIpIft6vfTlXyJv7LjNaYVW9Y
Re4DvE1a8an+n3CjNIHWigH5zi40dWleT+DlUZLJDPApJF6sljtw/MT+Bg91h9lN
8ObwfxU6e1O63jrUhuYLpleLa7wBgcXKfPgOyYpTmI91Zc0nRQJjHvyw6a8TJ7BV
WaNKoQkMOcft6M9D2EGP58ZY5jjYqWu0eS1CH5p7FgPhSmV5ESCkYwwWtQYdxsS7
nW/FYu3mOO2FuU+9HYp9FIqYODVm+QP9IOQzBRpmBVHwE68XnDnXjsdVG/Cyncz3
B0xkDdXS/zC6mjSUVnSwDEgSp3d2dubdGv+NN+MhnrvVuc3GsWgeQNGi8C7O5uUH
J3OKsNDWaliXiIrLpm40Cr79WuwrjoAFD3bS5RHieLKpPz+OZ0GUR8YwldaVYoiM
A68CFQ7LpDI7/a9pCGHQhVl/wNnG+XZ28WivoxkbMas5KbTHAf3DWUpTRFbFbKD9
ww3PxTzJXdvaxk6cUjcGbse/F8dnpigsOv9+QyxkWEpiDvaSSsPQmGVB9BW/8PEf
Mgk4QWnApGHBZSUaBkLI2HGnZ9zzb+bWS9qmmGsRIOtn5TtFBHc6zLH/V9U8ggsJ
ici9OXfgnZ9W05B16BOVi3rQgqnr35uC3qGkzKw+4vjEv98raNTWiIPMbiyeV2/0
LzNLCiW1Q41M7EVd9sKFGfRKOkO2xOUDNiVJ2l23vouy7o/9Oo/cBYU8rsDTgL4r
n1wgLF1l7UWHDlLpxjuqL6CJkheYnzQxGb/aDaz0EKglyUuvGb3ed/zsHy0+tQ/5
hriO0yDKt8WBcIPzDAJmY1nYadYsFsbCBKlNKhpZ665Y2BI0bCz8+NYiZZxajbCY
DitC4TS82XC8wN5AJy4Dm0gjsD67DhdJUvSV8e/af+2+VBN6Ujw87Q7dnOvTy6pl
IOMlRu63zivZNjkPR8k9C6q909foL30N35Wo1qdZXvw3rV55Ca5BxMRzAaFHKQhD
qhx8v96eHeniSlVYPULnfHqxS9s5BqwJKaCmNelHF3HAo2bYHNIE1RRb7Jagmz9r
DbdAAPRSxLH81U6PBMCoVKwp5AWz9Ige/Iz8VVmDrymMbs6VoXUhGn0mmX7dJVuF
IZNOiBM2E3OxpUUfmIG9K1bj2/TFsv6djh828pxBhcgjUr5hJCkm0nRuaZ8m2q0E
5pXkbLfTTLzudNfLqHhedU0xVQ+OPsqTY+mvDEN8d9vkGw1K/G7uMt2Qk/0OtLIo
A62wJqwukOlxd5P7A6oMDu4kQYF8bWhV58cso05yhdzD7Z4nQAMcITr79WmPRqQ2
18DStxBg3SoTdYucly6y478Vlg0hMqlh7IyIVgt2w7zgJasqDrYYjfyqewkTAAQJ
DZ2RbBydzLX8ekENt9jbGjRiEtRbqhqQQLh/tDCCxVWiA08ZKydW7O+YeAROdKLo
DyAE1Ll7aUV5jFF35Uc7hIRaSgZbrJBk6GpkX/FrcFbD2IUMmvlb1QvsJzU47ZMe
paQuvRpJGu/3Q7MluFIcuntZmhliZRxs2gC516G5SNDe9rAH6GZfDbA0tocES4Dr
dYy72uMSWlCy72DtYRyKV/dLGIa3e4ALuH0eDSBoU20tImL7NRTLkR2lQXqvg9EK
vWdT2+TKOOmKiLnUikTUpHl3e74a4n6n5oxHmLH64qXwb2Ad9bsdaq68u6mwM00n
mS5gIpOWzA9llFzn3F2iqEku8AIo7StmlKbb9XWAaiR7eCxTQKEj34tesBQHK0MM
u3m4V4qgh6Um8TrEchdoPP2FQH6t9mHWtgDBwqaVw7OvIHmkhCg2pbGnIBh73zyv
PkRkEXhIZoRS15r8UDialFUjOCUULRPvA+qPkiARX81GAQQzflMjA7Vw626BUu7i
GjPmsaQmZwvL1pdX9twwHTX7oasrGb9tbOT1bjGjv+2ImIThZfJhSkeoksW6el1y
A/J/gKnRCNIuRmpus0h845aZYW2JdstHAy8rp9pW5xq7armPIMm57c5aVySyGWua
DFmN7wJbOpmzGPt3u+dqSAnMNJh7YVP1kS1FcjYBWaGsqlI2QkBWVsGC80o2PieV
/XhKcTTifW084bjREclwOl9rfSxGZVqG6Gg8533u0SPgTdbowaq2bT7hldEvgLCB
PYQoAZiljHsgjW1/7LYi0VgdfnCdfM45fplsPO80ruSXoTEra0godUD2qBsVI+pM
IIWjAK9l7pB1Frz2egdCz83b1V9XUSpRIndbv0u1qGSgJwPm0e2AhssJ84/S4eUm
+twvgxx+exNIyrUCwN/ChR49zmHk5UqpmG/lEHvSls5XQyl1ubZjnE7hKwlkIxsu
6XXhvNtX5UlFwG/jKl7imANsYbaXoyMjjoFoJNfgs5ZQJy4NQVLUn0K3Y0ZD7rYt
008GfAfAgvJyYSp5MyfIiYsd6Ejm7Be4VVMfFJ+CYt4qZjrwRZ2tYE6Th/COZxhI
biKCyX6K8yFir1VwQB9GmcEaI0N3BuZdBylLaTwQPlmczoM5gZ5KiS+Th4wtpz4D
MGKTyh+t1ILpIE6mh34ml+jikmvc/t6kgYVkiFgwRbQZuU5WNFrNfvBrZSxQrTD8
M+3pTYQA6AdTs3uifkF61VNXPEwNlTqk7l/rf4Ynq7Z3CmOXDlYU5NKz6ehqUmF8
yKVeomSUgqdZOfa0L5b4f+KuJmKSWz/UZjC9okyopFPlKLhoCNStps4UsOJEHyCN
/8x0cJtzq3m4PTGSb92mXkG4OG6Vj7KvAo3aqP5zhdIL0tmGWpXhnH1jdmHFHqec
4DwCC/77cftmaLbj//V5f+g8UqSXGAHCMqn3S0MEECJRHB+SVCLwKOyuNJv8cxPr
m72d75IV6UBDNG6zLyEKaZRWsYNPZvN/lzEQvzZcVdVGduUWYN5I4JxSrmSR1/LL
w1AAz6RvlRTQVFX+vtHkKUhIXv7x3AIrTCnxOCLZIW8B+qhaMQEehvwJbE/LamNt
4yVd0bQdI3MhMsEBZpFG6gsDXlmUIsVHG+KfUVbEJFb3RRx0EjQSbmR2ctht5TrT
oAnq4IeWa6dkSUa/99fm7OAUB3xwOYR7vpY9h8LYrAZKweWjj5njKtPGdFlPUVSf
NzyHt90QKqiApi6cyPTFp9DQKFezC9ZdWvvLFQYvoxgtVO0BuHBd1WGNe9sf0udr
/3d/ThKhKPq9tB27/SCYyS6u/xcDn00GGKMB8dE1vGBxUcZQtwGZceOmpd4e9Fbw
s0bjCKgaPv7xz+oqRwbnb0A/FKWmNdOjFm8U1zYKcd8KgQIYgOPSdpcInUGUuxWV
tagxs53aqsz9J6PvudNI52EmnqhO4KtzoE9pOOlmLU590dLMcnX/RQXIsRFJJ0yb
nmWkOKqJJLiyYdNsCtaBweOvUwfxycm9gjPqmcGkSze8PQYFz/FrhlPA7nergnJh
u6RTNgOVHF/zBMvA+6/VyRUBo9zWXkEDEWhI4Ip8K/vp+CRH7Z8qfyx7qjFPat6l
tForOVsglN1jXnmSzA/7zPjuALHwlqzaBK4yTVVAHfsbm0Cr/41RGp2oi/yewwnm
LvkA2ZLUCdurOCi9q9x3/EAl3YO16gWDFiNayz2iDD209FYU8S/FQp5dQmK940W8
Qvs7oJwq58WLGLvDWeKwbwXIJYCp3+viytp6WioEj0Nwzb5Kp0tfU6Ow5iHY1xSb
c8n6W4XaACbdqTgpY8XMBMm0Sgq/lobjvidRTelJRqPASOSJZ0/Z9fJt9rZlecR/
7rxgShTcNnZLvPcekmuYqfpI5YlVkreaxhTUcIcb9PyQOrYsyZnHrC7TzDDVqBt9
vSSO4nacDsumF6Ekpy/C6QrqN6QxixbVbMUWwZCc4UfOVvydMW1WrdR7XQcm3JxC
5X0CfzK7jDJyTerleUK+1hm0NsnqO9s5ApWzSA9ceXO3qvgl7G1V+hp/LcQ0O/UK
2Ave/P4njGMWzoaMxUMNCDGSonRl1QeBvAn7Qk7UakjW4P4h/CPn5C3Nq1kt8DWY
dJ06S+IRSsoA5RZeLU1CvQ+T9kS3it0DcqSTghkmyO9pYv6IKyexfguZOO+JTlEX
S8YgxzsFymZsWFtQuvNXkGpZ+jYu3f6NdviWyYXhR7sVYv65BERjtvsQ1V5v4i1Y
YVmX4w/Ej8nO4vOalALUSO0/mjT425MvvGWQpjOhBaqMlRkUVk4MlW+RISutCdBG
Dbpg/0tUsSrSP+j4vKdm2MMHUsV8HwU28C8J+cjzjA/xgO9MNmJXbictU7coL0Ay
R3HvZ2DpiE/TONQOUd5Kk/sblQjMHdQZgNe1WWPfcZIFy7++ed5eUGsWtjjgrbzR
GkMgu1YTbBIpR6hnWZGr/AAfPyML1KM8smI3f0RL0AR5JIFmSEF+YPSd/LSlqZAe
/l0Zt/I6HnHb/qy15WzekAMDLuoB94BYkFdsRl30MaahBhLVHIZj+jP9SiSzOl+e
RyPtnbjmJ5j89eZb0QXSQhabRfR5vQ0lx2L78DGmKtPplucTQ652yKDAr2TP2wOa
3PWc0vUiC8kHa4oWjtCsOW4fQ3QpYafqrHt7zSy/g8ufRu4FeySApWMaMk6n4d6y
AlcMa1ekq1G6xeEkbkR0TYDNo/bmAwQ3SatkEoCj9PvNTr1tOiQv9kh4xfqvCkHC
Klgj4KDXI2rdvNtPBp/3xYHCMUVERMhcoXUAxmuBM/4jsIm/ki+GGGAAStJ654XW
HRThCTVydQVV4HJXTmsZJ80PM6VfFQhxuv5gIcgw8uj02dPtbCyY5AH2sME8kDmT
I+Oc+4enuWqnj83ZZPxEFxLKl3OeH8PhYyuwAVhxbJK3O7nHegU1sPrLXtt+iR3m
4jR6HKUrPHRqeTGBT7O2IxMyGgRtcIZXwjb4X2qCySugocNEaU4HWsECZMKRQuaG
z1HWXPpLBXfHrsz6uF2Vxt12dWvM7jQJCcIoE7IRahEh2VXQMkuTVASe+FMQg0Td
vQ0tSHPkEqKA/fr0ihweNbMa1UdogUBGaMtIyfzn1AKojvfaUJrGFjNiAZIASVIW
ay5e1b6R1O8fSK7vsGrANlGyLfh+HhL6/4VO1AAl23ReqnpsysU+7HSqB90lyaVl
569J2QV3AT1ESpSmvjErWo0lq6llhOK9BlyQcwaL3AE/uE/A5UQfHX2CsVVocBVb
tDNQS+Ut78gAqNT9MMolypPnU+XblYSCpCrbKn8l1wzEruHqj716wFg37SnrecAc
Dcz6dGoCCFsmS5wA4TMHt5F1ApTQ1DPAczZAe1hAlA67YV4+P5wTCKEcbbsisbVh
UYXuKCXsujjGnkNAkQ369HgY+SNU0f/3FHkA4Vwi0YdIz54qR787ogUwXRJN1/Pt
D2V/23wB8CORUkSiUyWcpXoXuRXO2Dz8hd0aAOMj7a75yKeI9QDkor/sXtsEVZ4t
FuNeANG0i2DKw1AAuSMTiKnG2olDC9dOd3XeUXnfXRQOjlx1yg/KenhMj1bu/ldF
L/KjaZ1oCPmheHYIp+HM77Pncsu2AIK4xfSX+8tcR1XNN0GtOWncBIMdFfk42Ksg
sf9ADm0IeHTfMiso4krJEunss/i6ei35GP85Dl2VrLI6pxQVlGT8QMDqW0H2BEvU
1/k77f2nuMNGOjaug0xGvR1dZY6U1r9+ExGcc39DAAujtbUq9zNQ12B71Fds3nSK
9eZl6VuE5BTVU9CfT1wNl6AW3Ms69u/+w3xf2ll+WnY5jL5kme2Yvs1pgjVAWzK3
zRbZIaddpaSX3tXsUq+8CKwQxIaoYLexPuEedmmfS2z05fSzgVklm7z+AgeiEOwp
ED5XsrRL32aROcJhjqv8+EVVWGgcHZnU5YpaBFpeiZ4PE/GWzPx2Q+pr4CNTEFh1
Y4au5+ivlwt8J8eAjvWWoj0UPxjDy2OHtIrmwgCrPFtpG0XjRYKzl8Dcvn1kfKLQ
PLvKCDt692+Kg53UnOjyVtJ8w5JmvN/4kxlJR7zDNQHhHm+rNmGBNociJgobB9A2
hYxsCRthZR2XXwkbv0cCEuAl03KhMaA3JjFlSA3I9xOmiQvaCxyttT+QUeJO030y
6P/szO2/uRLt5NX1FaqGompxKueUi10fDyvGOop3NYtHooDGiHAHN4vMVe9J3F0E
VXobfHGM/H5qpqZxbvJqoPrTFSq2v2f8H943VIkvNg5xRGvqG7wLE9Kp1tNUlAO1
fv4pzbDdh7Y5iWG5xaizWzVlAiuiLWXRphqqHWE2VXOsycl5AGd4W5PB15mIYc7S
1/UllDJauXB0RRHT3HoWPnkCfD6EJ2OskQAoDf5XZHOHRF4NQVPLL+RcRGujY+1I
fbaCuPwevJlIyqjn7uCUKsaA63uzWxDnjIEzFIqVKgAGDfEl+sc0f1g9sbLyYukw
weGy67Exx7xVU1J1PYQFd6a9cCdSM+cKq/kXNRwxu/OkPc7F2VjbbYq4D8s6k8sP
pnTXhHWfu41gAzu+vflETcrBJWyji9wsdD3NFbSRA0ej78tlhkffYepD5B7SVWgy
/odubST0chjfp63DW01T2t4sfslVuyP6DPKsCP+5BfGB2rPRgUbeEM7XA4CA4goY
omDCDaFILPnj3X4mt8aR4hzEOzUqr8edZRmCte7/nHd/vulA0wrz26HKl5k5RjBD
QIOabvF1NLsYup8hK6wca2RPcwHtGOjJaAfK4TJcMgVgsXZ96UnV9C17kgRuVWXn
rcezQQiHsVcjZJ94ss5K2QCUSjLcFKFw+ZXp8iMsgj7ZhfN15K+2JfHUfYycsRw/
1EsJ1v8yR3hAuOu86YJQZ7kL72A7YCwEsLDZdHZf5rZChcSc2tbgrMAYYoll74Pb
0E+y68kN2zdRqdlH+SANVdt9VmqQIQCBKCO88i9fNiBwVLtYNVM5Wdo0P7ceEz5w
ZrV15ng37PxEfG+E8IYVnX335PZeLZEq3n22s774LlFqvwkHzSkjq4fpYKOXy8Ma
kVTYH8DeEv7SxpT1PkcZNhOjv2b6Zwbtb3SDeyidOv7JWhGVj1nIuZPvV8q5oezM
Nup59TmwXbYM4q90LWYrqZBlXPqCOVSfCKVuT688u0WjpUurrgJbT1DSJ1Ii+vLf
WdU3La4EnpA/neC5FzXxmS441oL3pF7WVJ4sABOHQNHa8/iw9AslXS+3u0ukhWzz
IC1CppYfT9Z3ytglBoQ8Hd8LUrtYJLRCWDr6L/OZOj9XlGl2cPWIcl6k/g9sSxAy
YRxJsMm9oMhOVmCy5DxQjXqKS+YYqYBCMRkh9T1K9hH+ZZpTYqSgSkCgPhiX3Phm
71mzdWZGlxZrn52UoUJXvRWRM4/0BP5TRpDGCaPdU2wdGW8VvixppyG5+F14AeLd
6Y72dL4Y+eEDvrYB4Nl1qQQt5WpoiRWewONYgoVFqFbkOXfq6e/OKeLChXkTSA9R
yt9HeTatQpyDKXJihgm0Nh7eFvypbs9TiaDe+meAhepxDhS4P2/uGvCju/keFtWn
PE6GGn3JwA4T6pBXzb+GXvD3fvXNw6DykMzH33dwhJ8bwW5XtWsLsmLL56w0MMTr
r2yM+63LchhZ2zn3589JWQJ6E4JGTqEPOQ7R572XUP5dyNv/QwagfulMDJzsI81h
RtkwP827VOrxrUh4nvXpGscGiAuWe0CRGRRRX/phVj8eXvmXI/cX1gCpBP7HdLkj
v5iGZ6ed2rrSkL3h01psB4+auPWtuIpoyWzOAcxALBdMxbFKrEsb55uKvJoc5sUT
vN5NgBAXaifhOlXMPYM8dBX1L3cOqaLVv5HrF81/gL1u0bLmBUsROyI1T6FPJYWu
knrrZCud4WNY88/qx+upuUbxVHNmAJGUiJiJTqrV6qeNrbskrP8jeINR3w+/68dZ
aryOvYTUAYZAdw07zLjkYoBkrdqia9Nr/mx6rfrHR2aV4R98g0oiZ5s6he5hT7an
5yfZ/i1qTi96DF1uPggdZTAy5ApBzOYqvLjUOudaItOvvlfiYB+CHFz5td0Z+lZd
l/1TPeOcJvJfq4XDdnA3gjYUJaS6SASs1fsAVvpMDdTkXCWd6JeSHhPwRgvYMH6h
Xxp1ZiByc3EZoC0lBcbnEkC+zhlBUi1tvu8sCWt7BmpLuWMGxmtPDogZyb0DSlhs
3rwEAOp5ZuaLDCD23eM48V/IDj36MNRUmW8kamvkmxnp8A+6wTHxnEYy5saZEhyO
5TG67smv4ANzvTqLxAk+OmeXoUfc2TuRgGgfCujGO4edWiudfJ6hveGecjqQhMUt
9sKcm/KHwgc3/j9O6/fDgr3nUJDlm1kiyzPcIZD6jI2ZegUEO9Xk4MT2T3kmqZge
X3dYdtng7/S1//cnbLNtQ5l0IHUkNZPHXIKzJUE4/UhDJq4GM7trDb7aT7U87HWf
tUatW2jaRxfc2tx/TCecsDNn9FMAfJ8Fvr+7t126dRcBCWCB1LpOc5kWNht+eO45
CBE3dnMwKysDWQh3CpODvSObgvTfr+ntaDFTfXemoBEAhQ0QN62n2Qcn51Wx/5G3
P5ByR+gqCa9gutjOFoq+qQJyB4vwa+qvwZQEu6OO51ECIfz8DNtmo9pfO6w+D6CZ
Gt/PG2w5lAmwLizTmYRA5qrRXb9NEw+pTsQRP+vvyb5MZslXo+V2nNFiMH9cGxxi
gpFaOyHbiSCtVeqwpMzxlB3ARLjP1eqkOrFGjb327jbKrG0raw8mvJtNC/N4DnDG
1oK0TxE8Dja9NDw+f9NWEXy2WAGdhFwVx2S0mBsXsimlDRv31+8PNZpnsjlNRRl1
+wx+eSdql9z4OlN9AP5vQOJeJCNa62jv1FdkoCRz4IZ06iy4xda/fEz5LYunglHH
idtlWJDE7d+EjPiuqH0tPtEFjE+KPsrnutf3hM+PPjAYRO34mVgqMc/U2C2lfM9z
fBMGzGtDtCGcv0SgjVG/KuX+EczcqU+f3h9ziTuhizM6pFQylHzIzzqt+C9QdBKS
7ZlsHti6NTA6JOdVbLX5rRkA9/bZ3zgGwvvLlip/LVpecHGFYvLR2NzuuCT93tDH
oZWz7pJJ9kdJTAlGDX5F+ndHqV3qT7SKI+QRKA4IqfbhP0BUMftAKk5XT1gpp0lF
Hxrq3qlUTXl1w8FzCGEr0clGdqCiHkeIndR3ZSgQTBUv1vDg239nbZUDnW3ECdWM
h+tJVKzPuh0b9szVnQ584a5gDpEoYPoil/JyuKNMVbuZDk8FwJ3r79z5JXXB4oJb
I7BFIR7yKJN2jeYcIqTa9QVeB2yzjaAQXzhJL8j3kNlXKdgYh2KF1zFaXUkvLS6N
mYIKRb2w6Y4rPJcqJtMY2Hg47354I6/jARnvptqHwtJGpaBs5ZG1UlWBcMxCfFR7
bem/3/SSHk+cBIMZzuqffCOK4nkS9l4IoO2hiqKYc7KBoa73pUKAK1Ulvy4t5+FY
yF6R5B3ZLCgsJ6GOQ6xZxOPirSTzjUyZS36kF5MfzfC9kUATrbuVvw+hGc3LyaSk
3Z4kzLxHw+n9S4SkfoUbg2AihHGIT6iY4/Eh2iiE7f7POzXCh+bh8pTKZ0pbs572
20QHw7/yctnF+dX9czwEMV+izIvW+L6MJAj1px796ZWCy7imGuCVduW10SuADPZa
R++2M0jREIcYSS1KgzGAhwPJ6ouDva8hOmpcaH/uQ/aS2IRtAyZSJaEbcxIMLYwz
kIT3A0KPbbI0UeQ4NzyKf62nuFY3XR9vxAGtbO8qrbk+GN6gBF1hnCW61SlUwjcs
dcRoA9NU/ccTksvyu13NHNq8huDnoyzpVTcqGpbM7aurGzgWakO/UCUdf+psQGgM
8RnojjV+PI0Zzzmgw2r4NeNsx8GZFVur8HLug6sZpJwRtTKyYBMHmOOkTCHENSFn
XlkElPC88h0tzty37DiF163/ieMwiyF/TNecMDtpYwZ4QlXV5WtZCqvMAyWt32p+
ytAufMaY1FJBxjO8eqkOdZtg/PIiyvw6pZorCcroV6i9ZM9iJOW9J1cgU9GGl/Fx
EOytG0U8r7j5J5bi8+OxyW6DDunl3jG2/Uo6bWj1fMjyvPHBjj/b3IqfIFWUYQyi
7XZg2cohu9+aI1wpb6u9+QO/Gc7Ym3+gAr177VSaCmWfmKFKv8j967TPcBZm7k8N
ZGzhR7F84hjxdnM92EmZ2OBHpIOEFBRuXKe7WkRx6OFe8KSbr/g4OJhTXeusROJG
9l/PH6kbUeji3ZOaM9/93vY00MnHdfVn1VB/aAcuJMxabTYmgmXI9jCQue/twPmJ
L/CXVorX+Uga6DHHQR7DyqaxJ9gFBxuhtkl5ICDzJacASsBHSxuaKmtZU6eZZHYP
EICRidRCq899Mr8Th/tx4ofWSBFI/GTKuKwb2/c/YVdLjU53eEsmUvT3oLRrlMiT
3OYcu+OsFOo6DGnX62HVqOXdUq32MLGSvqqMLJZPn67A0HeqY1P6Du/nIydY2mul
g+XZdsmqU0F9Aq6/Ucfyw/+ju9vF1wZ+xp0WEeBr3ugoH45F8uWn9YnLB5fDDZqN
8qO69Nr66N//Mu/bf6pXCLekLIXFGAIGvYEBkAo7IDe5yMRWwUkUzhy6sfi2PqGH
VIFLocaXJf+3OHqDA9G+J+dLNhjmxKhaibMeLdut63L7VRsZUxpSmzyJp6mz8Shf
vl7dWzrvFCju3O89NgrsXx7sxgu5SSBlD+v6RexNW04Ao55zV9yZblI2LmFuu6oO
K1B3lyRIfhLxCE0aSVplu57H2QG80pU+8ebV0fG/ZIgsOcBqb9D7RFzoAvYIx2bK
D2STqTzgdWR0XAMao+qRmZeG8cLQXntewWHZqgBYl5b3U24qexUBRx1XBZ36aiwH
ka/uz6q/N07jtTZ69PotBeJLJ8gGdxb6aly6LwAyAbFM8v5NZ0lifZHCyA0tVLnB
GZ61qtOvtO9/ALOm2swI0jMlbAsZNo+xPEUUry8wVItjCYBdNObHe9QeZids+rZ7
xV+TWZI3WIfFvMrP4GsaHBkOnZsfiw6ImO//7WPx7sg27SkuOvUhRWNevSktq17a
J53t4bA5cnJjw9j8PnfZDpaORzEb5BmCQBB960768k1+cv6hJ3zgayqv1iykyBi7
rcFFORCgIzPRFsBpkzLlxXzSfaFNMEJjc/YG85nakk4aDsdrbm9TBxy6rYWUQVEY
pvjRNbHDzWTaBuAp67bsxXxXThEg6Fv9yxwlLUHsl4WRJWNOzHMY+Z65UD/ThTrf
Vk28pd/i7mqj+yGLzlrbkskD2gTqkusF6gvZXx5GfLAu14PKV2nfdkJjTrKCHFfH
h2MVac1FeQo5odICjkCGU8BiA/zFS5G7RwlgyHnLp3vQYGEhdGuj77dDmWSc91NV
XMytKO+oPjKAKtFPeW7cbth/L88LfU0GAt9Cx+lY6XNaOLtk0KLpWsCQloJaejLf
+p3KZMX81jUMCR8lzrEkPK5saAa/vcBDDbpEHF0qSlKKQl5rpMjunJm886jCOXlS
w3WWBLEV9F9ua2t8n2CYbYOl4k+JjJqHmIwxej2VxLhophXJHkp68MeAb+I7YMfZ
Ly8JoiumjYjpfwCXSn8oqKwXE+WmKGPh1OT+fJxYPp2Xdd5CC1EuBuHQfCCuU+62
y/tWWrTZ0VLADsXRaXMy9vIDj7WZ3hOroFQzTFQiz25uTuBMH9FFfG0QcqMOsm0u
Y/IRxAoeEqjL2IwYakQuHJYj5n+nR15nOqEVQUhWjfhyJv4t7Q7y3IshhyxGo4SZ
T+AhPayV4BMi53tWXEa1iYKua1361VbF4a7Mo6ke0HJKqTuAvbdjCys1tAGqPLiz
TFz4u6CMhbBqV4F/vmMVasqtA8mtT13q6kNS833Ucvv6vUryMk7+bn0+o1JXK8I9
6L0UdAV8xkvYzHhWEojhdTlSVXLX+vJxUDi6cOXuK1WBesKqx/J/8uz8KVUK+0KZ
wtHePEzIspRsYlycvlWwLgPY3c0lOwEkHe5bE5XVuKj3zvUurY5WwIuN92qKmBUm
5mgJO2QGmcN+fL+MwpNLWjgmZfAntH+92eg6ZoJuspSQXUKKFRSKy6h9R3VwtXjg
iJuSWBYwn15E3xi7idVqSHVaL9JseR9ji2YzVejw417RzzL5wBSAvTsAtR+v5zIn
ZdqGQfs5oPutyNUnON/J+489nJYOI/coiyNwEKP9Wt+Ntph7hW4Db6GUhQ69C1eV
H3+D18+MQ0a5zEJmh/WQ6MdxDacTh41sSzF4Iq3XPhC2cYay9N9uv+qVmUr9UcU5
ffWDIRlTZTD1Y9orjD3ZRDqmG2mTq6z7AJH2CMmCCTSbGvuwPTmB2kOoBe2T+Yui
Qyhw5eT0eN71X0qrmN/nwXA8w8hSL7O9RPUCa+v2IB1FuFBuH0dYbJFjq0zetq4R
0OoUakwSvLqGVdPYVzAMl7ZdJ2jMwMA8FNS7gXSST8kq/t3KlktYR1yzqlfKfpcV
du+EwWvLtRTLK9Fr8qmJ3rzraRT4oNW0w07tPQmsNrfbbFw9MZOapefC59nrWl3o
1ISC4mfpLMuGmzAB8kM41Qi04BTPZCDeqj+QzGSEBxc1HRkj/8mwb4XjvLVlT3Pd
QHc4h4NsCMjU/zxbHwhBmGOfakvy2ivjyNq/q0Nku62I+KOIfbTQYSztd+kf1rCa
kb148iZmgQz1T1IZLa1uhH+KVsYa1AkL979lEceP4MpYCuBgCeytDBaYv08KmFnD
XJ41qfmkUxCUkxSz/XOMXnSIXv4fuylJdfBnddRIxQuX4EIE9JjDYOEqiK5VG9mz
1e7qBDBwrptoyCS5rEewpX+6fvH1f15aflVeGtDVJojHZWs5jN4PhrZAZkT8AKFr
AkHy2vL8V1Q621KaYncPzMOIddXoAcEfOFF3PouMbEqUzUl1BgQrQmhsYDDp2aA1
X05sRnOL7nT9DNScCllpD3tXgBJ9UIUTh8EJ65hb2yePfn6DRucBbJGI9LNnN3Ox
Oi0Os7Gw6LTc1TRu4sW6cU9Mu4ACxHXB9lhKohO3DCj61T0c2rjyF/YPzpoky1/a
ycdfK0CNNS0Q7q58I5CLLNdFayRVQUpQY4R0H960BqPYHPnqu4J0DDrFoIqcferQ
V1bcOVpvDdNXfZp1nlyMPaQlTgxLEwwzBtcpzN75RkVOHA3DA3ul9dpll5f5minD
W7T5wLDQP8DgUwftRTzQ3maTkkgxuFC1GmlA9zBEENF/uadcm/DvB/rLi0+3DkM3
UQu39f1kNVctQv3SbnWE5an9ixWvuoDKBKwl6gGBazn4qX0fgJ3nLRlnj5bPpZAI
UpXi9BJyHbXhFZ4aXMZLzAxNTZRg5QQtu0XU+dxVpv3+xYn8Z+QIEuuZkpLGyIDF
eQRg9nKUID1/k9rc53AJkiFPizeaW1iy8y8Cz0h0ehxxEQy7czSamXHTZ7wRNeES
AVmruv1iLc+LdVak49T3Hz8uBP8KFATB4u824vOC/tsDSHbuoxu01IawSO4I0/jk
q8JXrajc4hIz6+l4bfIO0hgHwB9jgIDb79F+FBecyNAu5uN1E2cVCEnlBCtJQcYP
IVsTDSnquNA7jwP3pQOb7NU9P6x2254l01g8XBgdhYjAOzJjRVzcwDnyJ0QgQSPt
HPQ92aheQQlZjq2w0RRb/s7f18yZN4ZcrJ4tC/5a9d0bLJkSp455uUZD1A1AAkTb
qPn8tOW6YSUzy2glTyiLVa/nZ6g4I3kgjawJXDQfgKNbgJALuqIOui7VMCa0FypS
/sEjuxvKzUHywAZJivD7mx2Jcwl3xbdI0F1hHNYM4IYKA0HVjH/A+x0lqUyrrFbB
eCZcsZbxUrDkcl5pPQNp75jZmXx5Yq/gSz2rL98jJQbJFthurddj7D+MEySYS7+j
4xL5+3f3A0nL9G2G3DRVaf2iLBxQ7i5HA6vPcGunh+06YQIiSNCrAC621SUV3TIP
3VhsCiloStQEsKxxjDmqO02cWYF674jmduXG5lYwdCfyyH2wlYjFJE6lhTDGGLPk
SjTnfgsVqlMjETGCvcbpvLCi1WoMKTXBvRc7QGts6IRKpETG+agXWrX86C3TpMhI
xxQmBS1+YjkhKMLOsbziEjoBvoEmrA/qww0nT4n7QCUUV9mbanEDue02OLLizepz
bzUYey1VesavRbDxizext5hGtJOeJKdWL5/MHeSjT1wax0DG7LCHk9OFQbkPNgIh
rff8srWmORatwfoZUj7Q9P5ex5UiS9X3HY4YQPNeJ3SKPvHRoGM3BqxICA4ktV1B
EnX+nxgjMfrA1n6bfc2kzz9aO+qMR48y4KrbKZomx8dN4dPuMwwhIqJc/Ly4YjkY
E41g4ZPSQqhgOrtG83y8CKVQTGtLKkxuvlEZQYVTUK+0q2p+BjZCjjQOWZaOVeGn
Prw4wcmKo4FAVxGf2szXIbkDQtMFIAuRuasa2jBS2LmCUb+z1VG3FfAqkTaJryVZ
Sxbxgk68FTg/8beHPdc/T/OFehYtaxWDs2aV5pNPgSdWhDht8EEcm2CNYZ7C1tJt
reHrFg8T+ZYL/aVMy3WCHXn6qPLAgR1NC8Fg1taw4xTmIR/v1mBkE4e2pRZ3eHvA
P5sR4NxW4sAZFNxFGDU3O69U1S7TxETtOZccI1MOgJHynqmjmQ/DBMd4z0wLzzD0
5ZrHPAZ+acNgDR7DCGi72UtEne0yKmTJxPjhjxwYxceG1XV2RCU0EQdb9RzbFOsg
yZqaxr9HYdpgz1rRh1hvfnse+AhbxPnJq+3j6CnMN42hSNbDSJI63XEFg4Cs08/W
EGlN0pdTLFwLZzcYYBNDYIB4K+sbaKgf2ysFMDud01yGJKD9A8nZd0xmEn3uP1Es
0UKyEYCJjk7ydspvpo41x9qZt/xBKiSzyrRt7BXLyoB+ib/Y2R8r+mfl/rZm22Dn
nl+CWGxyFRjGmztDtqU57FOl3tSZCbJHVlaJ6Q8B2JApjzMP6v2oNSbnEsgixaNd
Oy4v+GMoSJs32Ufexj1jzrQEgnAu09v7p1X1I83YQDag8xWqFEZu6Fl34ZMGTCUL
z55GOztDM7l78GdsuKDsEEnrHXgMBKjOmcAZKGSzPUZVnOqBVjCQ9jrRGh47x3tk
HUwaQHHS2lSy5LrIK1LhZNc7KpOSdBJyim7bVRnKnSBd/QRHHswXzRGvah/8QfAm
wnnabCeDnNw7z8MvcwtTnr9gKF7U3NDdquO39b7Xte2SxHYBQ+obMqVsb92/+hdj
QMT+fUPKE3czihU6f0oQXQhU5pTUO70ovCr62S+M9cHG7JyswN4iD1Sswqse1jiv
r5IBeR9LVtKsDkUiZWiKqiHFkKACQmkZz45Bbjl+76REzxTq2uAoKbTcFUlCI8rh
zR2p/858UXh/SteZNZXoO9oCSkFCtOsqQ2+RHrRwT3cTp4jprtWOYfNgL4y1ugU0
zM+Fja6lWVsyZ8FAcCREt6/BjVmic+9aqje9JP+hn3C4pDNmECZVp1IExfflD/ZH
iapqyMFRUCP0p6t5OXE2QkwuVixTZPqQuXEQam7FyzyeUK2XePMEOUaqpCzmCfLc
4uba9/LnAslmm5kCO7sGA3Tj6B3VUvBxzJ6bTY77hs60lbq4Yzh5eLOCXvpRjleR
P70KKaxnzjawynxqB0fy1MmlBAFbwChvgWMr90F1M9a64q42s1qR0o2gBvl3GJos
Kf2aNfrYeojH9L0LeDACSzKisAiFOw6SG71Pfa6pETeQjKHYXOEHNxlSdHUKZLQT
fxVpOiPfLZBEPNo4wYa5Ngvot1Kp/oCjOc8qzG840ImgfXrmT0y6MA47s2u7wuZ1
R3JvOVa0zXVF8ej3auJ9wdysQHqX2MjpDiIVn79ap0pedRAtZbajuSAI+AkXlwIF
HtiPzlZ2DyjeEE9eBExcMvF4YwIqFTA/SMRRc3cVETUP4NOwr/M9qpWHUMN5j02v
odroM7PMCcn/jALMqothmL0QmzeE3y8rKnaSrqZtsMtdzGu456tO0lE0+2cWs4w6
hV5yGzY/DG6M9tC/ycX+S68l9tCsKevkNi4JkhShasQn3fY+yv/kpwRuJc4ti+0z
r5f/iTCsX6ZJXE27CauHtf5hZa4cqVbQIe3VmTSE8tfx6RdYu4D/osVDSfzyJ9wv
5daxeDTVjBHUlM57WqijVXwkllMyghtgmWHK6bAv6Yyf850QWB3/j17aGVEf8C0K
4r+pRgXcKJY7R2BCRj5Ok5RKZt5Hh4B0Jl9UW8ZX09sBSNzDvNTawIAVwSCEOWbO
o2GKYEEDDfqPNmzFGtIxKsnbDyxuBXjOEnq4T+mOC9+gC+O12AEQ8UlqkwQ3fLDu
ut9SsdhXujBEhi/KYZ8+lviqg1mcMGqLqpk5KNHk1cuXMUZUS+2qKnwWzvU2Z513
JAbo0Eb+loD2C7f8BKcnJWb5OBai5S3CRWD73g5YvEYytr99dXw46BYcSgT3Z70q
40naYM0gzGsTFwPwTN5gqpxxP9Di3hLhbCKr+iFpzEKyBdd1emA/+owGD0JGGJky
f0BBVM0yLfxUSoabYLg68AKUIXMWNwy3Lh/TAjcQp9flJpGqU/Qompkvi+/uiRYx
5n8+lFR2PW1bd+k+nKkkk8woGKovRti3SMhGnahukUknTGQ20TKEc9GbTPVXFxCK
SbJGcdPmqkIEx5E/SiyzUt+OAHf2wS0dn6KtIPGWKBoioTBkRlOUVHlBeVQa95cD
W/2B411r8CiLQnVWH7N27lKR1fd6Ud//BEkaR/h/vLJgAtxmeq5Pax+u0CQ7yqv/
L5iHxytVScsAlAxf75EJfVFeM9WBVWAFN0izcpoNInPpz9wGD8NbnbGXBNKk56s8
nbAmeuRWSLqNtIw/ZAywgBG1VIOLIElzIMSMivzTQtMMaCTqukqiRsSObHTgRxJ7
nZkgmpwv9IAtJzYYm1lEuPr0DTeMYoIk47VOeQjCQSlYmRxlNTD2NRC1Vtt0rht9
dFsLt8n+TyhuZQsuPdvU8OsQ+v7xjp4Sq03R++TWQt0zwC2NpOSh6Rp5bTw2uQFY
hCzacd7XfOWZf4/2LrHuIWo85f+cHGPG2FvAmaC75NHFqEIdUv5knxaWHbnC1XS7
LSaxkQ9ZAmNleWC5sNDfc4fkAd8KhpNKY6eXA3+C5kKsgo1lV+Q/A7rEzepSLB+b
+a8V3PMvHaTk9xxGjwOXNYAeDYTZtkhrgHaAikgTnzRWIvSLEsvDA1nIlzvDPM3I
gUnOmofEiSjRdHbcPqxggjdY1hkwHH4jX+78r2dmVdG9kLIBA8X4RvSG19Wp6OR+
3TJH01EB8lU9Q7oaljWrEQUJb7cuCPrLyXCwyghFZQflWwG7T77Rwp4+3LV150R0
tYec1QOXZu59jveuj/BVayJ11eWvbXOUtg+nsg4uBBL0Zqc4MztRBWFdVa8+3YHe
N2LibVY2cOVqpLf1rV0UNnyQspgIbRB/WYfY7CyEIg626ZyoXK7tsZu1bUKR48Kb
rZi0sBIeFWBMK+hjsWr493NV+q5DHgXZkT8hQlKxd/H70jOjYwFWtxSd7z1daKYl
WUDZ+OpXl1mLKDgmhEiYTRc7gNgj4ltFVE44NiIdo+uUJ7Hwk8DYJakXCUTB0OGa
GRkn8yK/BVteOnwpnUWtJvrjxIzjml/9O5LYL/jm3o7XDLqjgPeu97GXVUo3q1Pe
Wbk1dwAtP3i7GUKMi7OW/d54GsE9q724raYlh9BYlIG0Dz/9nTiQeKDLIOVq9OXg
CiU/SlJmhWImkLVGUOV7Ibb5JpHm+CjhypLYxUZq+g4LaXNMpojvhZKGzxu/8aWd
9MeaWf/jeRvxIHGaNtEoHCfJ27Tg6bYNz9oE0dc6OAAl+uHaRRRAFWESVvIW9wn5
k7Qq0t5/z5i0lwct9jMR8U4IKqFJEeJsi4KlX8rynlWIg/YFyHq/ykut/JJ6r+0/
MWS2XMxNvQ2SAjWRPYN6r34D45ma5NTnO88e+IiE05s+X+AhfQAI8X7ymu1BH7b2
ALfNkk3L4EyNRuC6FhJmIzU+RtpCJC2G5Tpc1MNhcZnFJTUp/4jYjmsgWfIk0B+y
hBvTBDcBjwBDKKUafcz6KxtorjjEYQ3vVtR6s0+XsVHdP7T/vipy03CD6T+/rdjv
0u83KQ8AokE+zMv5ksWJUrHWlRB3gKcSltkvS3gsixJifw/fa75Zn4I9Gq+zgdOz
LXjI3TXFQIyAzzPC0yb2dhwUjYBPSu9kBPPx3/iPKJ0I5o3imK34iSaMKEZx/EvX
AKIzbYHCS/B+ESBJDU+gxmQxTAimO1e4PIDr4SbnKDHNAvRch6zEMhH9OBnxHLx3
1jB9rT0NMEEnI8aVkUgvDYT34TVWxoqNrUPUhiWpXHs1+/dhyHrwD1lUohbiHIPC
Kpak01ktQ2Yo7jA8f7aMDLtJjGHJ2bPRqz8qeMtw5DxKCZUzBYPE8nBmAJ6ck28u
7DBcDD79S//iRel6UrTNiyFjhEfCPWuIaiWnlHe34jztIxlVg+MwSLobwOzevbM8
DQ2eLJtVV1A75kin3oZcJJNHQ0WcVTCJY5dvYrR0JFJxQavKlc/MV9WcjZA4VH9s
G35n8+Sx9gReIQ9JDvyLvCs7lGcM+aYYsnlO8eoubA4bmAZIuURITU1k7RZ21EdF
exvTnvUG9putFUmWM11ASokKGKdXS1duiDrtiGy20taPa8AZSTwgX0yyCr2eAkwl
I2rxXvLd48LCMWjD6+0iJYHnu9NSsIb0FAY3+4NbA6Cg5oYNqULCoiDiY/Rndn2h
vDJKI8APt6cheI1fjwy08JrQXZU7JEZUMzkz5Cwg8WNuge1smW25BAAozlcDRY/r
XM/hC/dY/u+RRI1n+FgtIFdNCwQ+Bzmjd9Po4C8J/nWulkdGxe+kenS5nlo82MP/
Vn5em0pENarLLnVlPUbbjHMNPYidH1S6CBjTtm4lYV4ROawnOXPkUAi2O2zKTFEx
ccjit68lQvsbYVNkoWI7vY7ANSyaBxics45e2ZzPidO22IZ3hfzsJh2iUMDZricH
m+BKKgJPp95cRqUCNyP8PePiA21N27Dkl/n70Dbcv+oOKLODyTgjkJPomJo1vHJL
VIpE4uFbXBOofpWKtHmPHdv+pQtj/+r5sk6/DQGCFY2bKSHAL8chcBEU/W1aK847
FR33xRkHOzXEuax/ia4YWZQj48df9SbKGPxxFLTIE1keY9ipY/fKDOhUL18iJYkk
wsZeTcBGz8X5Mdjk9yyFB/wOPa9RXApebbOVp/RO6LiIC1pldYAAltG/B6bR4KCv
vK/yFLrhQvCSCEa2RkQOCc8pNM+tkUPSgskepjbtCwxTlGO9RrH2tIBcbPSXbv+8
hpYf1SPMY0j97BTWUDMfqd9tmto/ZSmcK7EiI7ZCmMr3VBZvCesx4P1uVCKkWLu6
qRHFAIIBTylLZ/hAR+WLfbUA3cfpF4v5mibszBTa7Eq+OO8CT0ZOoz/Dz+4hbU1l
o9BxcGlff7Wbvjx91+1q1BtwHPVkJ44/0SOwSlRoaaAvXhflLNm71pNXG2I244FJ
jmJ+VfMhXMm2j4olt/JF1Yoq9Dg+6mZBXVK0XXH9vkJwAQmoaEChst3YR1yRehlh
N/joewULdCg6gi9EWu16SYCTewpypuXMdBjYq8M09LH6UM7VhohuCluUJ6QSKNSd
DBN0XqkUIqqv/W1r8aVZwrb7dBSicJigsLHItGXGwdEQwKam0Mj+lNu6l8ZUOdBB
sn6KKE4Lb/W81lrRpqyCGMDVPf4B2+u7zgmhJKK+qoo8X461uxukCSYgnBdAwySG
Qcv9nuyfC7wkSN3ClRojNThUvVlzvRRTwR6/M9RNa/NVzV2bvlVJJPYCdPTNkMn/
WWeGF7Wtmj9s5aFbUlGjwQRXJVZtQ4r2qyxJd6ttKCE23ylY7aN4j0hoc3lln2LD
c3w43WGW99XCCAkECAAljXt/96QLVcLZG9Pm5Oy4PmQpMCorehV7WXd2R7MW32Q1
A/9giLm/+8PJRaN5vc6pQpzOrrQXJW71aUZyAvm4wDMVPQRixyMWDZwDOoq05g5z
Kf0AWI4DENExGEbwOrwDCddqtzzL9TmdSaEn2hd5XKIZcQ8U0vHNp7An6tGUbD+m
54bLKvOWaik+9O0Vo9PgfwmcObEKmHRbHQSKGwM6QrMefmRr8hD3KpBdXzmH/NyK
lsHPPTT0IG5pfpQlHHxkxv5IHjAaXUsEN8zBWS9Ub8rneC7z2o8gdcg7IhrbOmBL
nJGSbQk5+UXLZVu5zHw1iJCB3lFd/Q7GmxAlOnQqa9FArpqFjZLKGrbkJ6zXBvy9
oZ0BO/t81EvCMtxFe1bwFSEpgOBZq528ZRihkPOeLKRjFdzeCd3nibSMmCEiZPUT
mA8c8Oq7YrO3Uut/X3blREefxLoygfoETNRld+6QzeFDstJg5CLomVxXgZB4Kx0a
9BYnWe7AYsmROwLTSi/mjKIUte4DBCGw3uiae5uDKWxvhPheGEYII+Zkcp/Tp38L
xMCJMFN4zKHQgVC1R7yx7I9eKJMd3NrMQyxbbVTepnbVgy9KGYwzgCQSb+BS8OCT
QXOLSpwA9YXqJ9qeZp2oPbDgTzOiV6607bicjQt3jOrhulLLZwd+FvzzJMYaGMPr
hFxuqYlI6gC8b4LNMPj7tgMjPDP41I7d9Ee4/ed57FJJXqrDishPiQ3StYix5aOG
oNI6rc+zpQbaIIPcLGqGv03gBT2k5+B0psNqx+2m9xN7WzdHgmBNIyxL6QKUKyuo
yE1LDQwDROYoPRuZmUl+10DvS+XBwAVqO7aqWApOyo0X7V0odQKn/e4x12sp2QIy
UUOgf3k5yO+L1gvRc1o7WuhrMNsDaL0xUrC5NMGOAniZuo1+t+bdQoErymMsQZhY
6DDaEi+EXN6aq8rAVmKE0LWGZXZWAIIUPs6c++lWPG0Zss5wI0XocYFcaOJ/UOfN
WpR8Zb7z4abi8FKePktbdQLEYw6kNxfkZ6JQS8zLbrX8JTRujo5gWt6f7BEOtRU3
N1nrQvoYLgECHj5mWDCRl5+yk96fhPYU46U85rkBY0D4y+vbylOybHgSCLvCQ49U
Rnz8JssHs1nPE1dcTmpCtBsl9Xmm5uqfbkhL9wSU3iVLuvU+I59nscy9MX+uhkZ7
mmv+3rU7hSxaTF2Kr7EoQNNdVbBMZgmpRoGX8sGoaTPkA5iQILo5cZtPorn3KU/k
WkJvWG37h5DmkmgDJXNEEAP9GFQXWXQc9AeFWO8lu4O8z7tuYIF8YOHEeo3WAjR2
KiniXVZ2weh7GNxpsFHliJqcef4UN3rZMgRIUwoeFWmFXJxK5sORJQDewxWjcGAs
iO55bw9zxZZaadAhwEJrLeaqU7lLSCVXr2irrfqf6f1D5sX90eb1jc/R3l1Vd3J7
lBSwXc/4wHtst6apORQw9IQ90HYe1G0I/D4q62T54IvfajHbDenIzF87vY+Fe72N
T6rroOQQARk3tjgyTjH1RyVYmySNBnjOcVMWcpGERzk4Fg+rjhWTgrZx3N/OS31n
4k+PRwGoeij6hLEpGzvd69Wy9mCvDELC/77H4biPfVaMH+6v7xLXtfKYrSIWVRih
XSrdCaMEawU1A+c7y16ziJ+djd7TH0uqABtuzhIY3j+OMij4jTcYDw3MclUhvog3
YnuLi51qDH3EVDOTHgEqY9qVN/mQaXaiiogon/VJFcFdcYEUid1zMxVtJ0hgtLwd
FHr3sAlnmSmspTR6OaKikKfbs04hLztdPJaMUXZDPmZzoNmA/ubWC2z0sFnSwm1K
YDFue3q/pVPER5k52kNbBSlU7/cnEk96IZjWURLnvvS2u0pMO0yIFDwj8L8cJ9Wb
Wpcd5QHjPFzvCtfUXMSh2UxDzLPhj905g6ieGrsQrNqUL4TLL0uPWjA2BXDXrU6s
4xKfQn1YA1YyeBAbU29/L2b0EDcVEwiHageYTOjfKDcgFUl+iLFp+MMd9zus4wKf
Sh/fZyY6dkK4ZzR1WsNUgMCqWixfA7gokKtpQ/20y15+JRumomTRrtI3C/xl5nl7
WAuBHj7UG9/uQKnW2eSsr4LMESWssmeW0EVVWkDbrI96Dy4EggJXiGmPJPM7Yh9/
LJqV/cuf93H7M2sqWsY9hb7OGEa5mrugk9O39YU/QRXHLb3tpDA9I4iCmCovar08
uZPMOYqrj+BtrvKa5G26kR5SunvV+EeE/SlL0dSGZEL0AuHQcFtsnDqkAJSGU30D
BvX037ImnuMrbcJnuvg0JbfPyEtv0ir0U801SGBgSk/+0PULODoV7eWGsGDQkG5B
gF9oW5uNt5woor8Kcg6yPiRyiaAul2blSgYUiwPxPSg7uWQNzdcwiQfnxqjEfERB
TKX4vJediJpnfPaaZZvoH81oYbgWrMFNzDR35tC2wL+zRKqGVs38NcXyNAI/69xK
WFbMJ3vNyGmx4NXfQfkL4hWtrNcavQw8Y4+OPwUPqcHqn0c6eqFHUoL2oL4vogMJ
CLddzqu9R+I94gzWjVZYOrQexldtj6wVoAQtiPCJXGUsw9rClLE+rtVcs+FlN3Zz
qCDAxYj0xs8XWc/rGFJl4zyXuCHNnXly5LZhfcvaCfuaDAsNz3Q78SBJLAN8FnZZ
agtTG3ahboTfoFuyv4rKTZiNt72XYJ+sGYP6y5yiahWfhxOM+NbzOTagndS+czX8
H/5Phx0E0o+0jVMpSXU4sG/dmSBgcpx3PO8ryIGkW1ibIbEKTnCTVNuQqImIYhfk
4hI0OHZLFsoeiIueoMGkKNNVYiFNiSWTkwZ48StqxDS4Fnc8izHzguCIF59JYOIN
iylyyDxyJcuajkLnTmlDAzqu0Mq7B6TLzUHdN/kfsijr2qAlyXbtHbjLNI+B2sTe
s9gKWRHFo2ANDJ6mkdnKV9w0Zrtu7yi2UGDgDh1G3gXUOJlRiTYJq0c4YLnrpLdh
JcJ5Rwg7u59Nwz+TkzkCq9aV+YXXyvL5ItbbHw9cW4fDNwIzv6qW7NStMSKgEw5X
Gh8bzarjeGJ/hAgGhUSBgz5DrjilmzC1anGpeT26hQV6cjRgaeX1P92dDwo4HbXR
c7Yu9hvAZjl9VXPe1jgt4mjgtG4iss1ki23RizbhbsGLnOqAGmRgakc3TDEAwvW1
Zb3IkZevR5ptQKZAlURrwPvLhvaRtDmeRIKIq8Y1sjBBUkVYpqLw+s8Sp/9uLwKM
Edc8QxeZQN1pHJqO4nuX20XtHBnIQEcNbLT6QDbmJwgdddKFAKS/EK1yti19Qo5L
+uP66GBnQcHVJ3PDnlbPehnTUsj5njvOpdEMqBogde2FUZql6IRl4Qq8g0oIvEk2
vmjXE+rcq4aRG6UHLF5U/FoGxWtPHdUKfiP75pkbyJfZBxxGnr7fFUw2knKFN3ZB
TVdk8SEPrMAOPtHFHkmwEOTajB9fJkPqFWBHR6ag1Cs2NtYfQpyZYbXy/88OSwpe
/2kQu1R1gbryaznD7099jRR57mFYv8Lbi2xy4Ez+FTaFnlZWzLm5p6aiVikbwIqF
pThNhdWpmhBGhq8491j8A7Fpp4DcFzjgf2eIPzkGtQEtt6NdGFYDliiTiZmQLxVA
t4CNFvx7fNgBpxZf+5OwkRW5IH+2KumtxkK8EXt1ln/FtHWshxGOO/KGCJbvgqEo
nrTvu3jm3TrJvUyDuyp3X/jrYPcIHmF3TWskchisOwY5bswEPmBbL1iIHlchLja1
5sKNMrOKe0JUaYPABwfct5Lq2zi3bOiFkI31ay19enAmFbuJvvfTZfQq5Kl6SlVr
Y51yyISXU+CdNdto92xJzC8tkFcHQpDo92Ng4O4dQ04GkUFnYStBbrakz+F+BKWi
WdvqJOF4NMw4tZ10v8mCdFIDDODnQEZhTZTU9PRQ7bibz0eC4YVeZkZvykbbt7sJ
JIPrfYJMHSTSgz3W8vnkCO8t8+KCFLSznRUo1oNf/Vmtj9kBIdHCdWCqLsYGnZa+
2Ulxv8rp/uC2XpD3v4yCtrfTODoR42TtiwTtJuC90mQ02kp6hDqw1lO0cL8J1gLA
VBlivSIVQtAob51RT0lfDM0EnuB8FJliebqjFI3Qnz9QLEGmk8IiQZyp4N4+w6Bg
QS9NsPCgVZKgesg+4y4BbqwL+8pdYJkosEDNvyYuEyAxfuP0X8VNxBIsYKc76atP
4sNGUyyvC03+8zjbeUhnGZZu5ww/Ku7n/T/HKqv7O6DXP7k87JxPZplmeHE2OxBZ
rPD3Dyb8DWfw+Pdk0iCNNCJTUL9gH4thpJXMlc3iA1ysRsymcfgTzEOygnmHBdIe
h7QVjWx8v+kYFQ0qt9FSsgmV+ef7jE9Y4bUw7YKR2PY1fGGDBpxxyAihd1ztMFbg
K/w2LULIEA2tvlBa+2c0uykpr7yB6ENdOFzDhrImeylQGD8OLl87iHsZQwJdNHti
6b0G0slqOgxSM0uW1lxDHqwKyqEv3T4depN356MNukjef1tgEJaNY/jHvPgEMFfy
sjSVzxn08rlgb5MjF+uVf17jGRY/9ZHTGuKBtVc4ZP7AEl3vuLxVGikbXb0Og/rM
mOajtUhsZwxgyXF7Io83DaMm1lMHa6kH1nA1djfterTzs76v1P3xZIOoRHTlaxwa
whzc6Mv+VO08z43Py4eVNzAS0brQMntkjh3VzqiavxnPedMF2F0VXs3/Qw52CZ2R
mfesDpFoEAp4V5GoswamMFjowiARQiuTqNQmXUa0Et9Cvhs5b7gKAlF+mWlRnVje
UOoKn6YXPv+tz72QBlyxrziD0v0pSFq/7zpj2uaksW4+tAlfqZdcaO9OINv6pTv8
8GNt24bb+mdxvGwQuSyfv8N+fAfCFXXxzBn7G8p2EoUr1hHS8ej+7x3GzZUo8g5n
jRlzZk+Ps+H6fM/LVDgyPQ9HBC5T0uOuauRz77AGiPzjmSqeJvhh/orJ6O7z43ww
XFUh1fojrEirRa8VlD9F5iku6y1I4ldO2K4p81shF4HTTVzIWC/rCGwyw2tqtsYc
qGZS+WfcASnExOqpDnASTsdmHR5MI9KL6eGLQ5Wcm9GRFSisBuauXPVHkmbhWcYw
XXBpr9TOXUCLXOncmUIo7WC4Cd+PePa7kh2ofv98JBj3+SMoHTc6KrqHMj0t6Qtc
PFJQFjXLiNGN4Cd4E97rZCseB/p23NsnZQi1VGpmkyUkqMmTrj6TcpX2x0xj/nVh
tKhnXkBai0g1sQQiolCLbHErrm034yMZDUwKGuUjm0r0e565q/Ihr6L/cW8ZNmJx
3VbMaAd909Y/eNF1oBkwlvGf2S01UltJSdQY7iVB264Q+6W4tDjQzZif3whxGET6
fxA8JLiTOMHiYJIBPanevCTJExd+AielJf0sLF5BpOtTm21IU6OX7efyd9ObpXgv
SNz2WsZ7nHbHYUCwUOCQw5YxPCnv7VjCWVQBMxAAS/Fo96Qg7ScbDajhJGW77Gx7
4j8IGuyaK/iWHj4b4Zodh9HvmUuWBsVUhA7iLmanYmSpIU93sHX6RTNRi00fDSKA
tEnNC7A6d3A+y6lX24FzAbOpg6xq+A48ZjvqjtEE9H/XvDuYaNXCO3y6qaQY11oZ
LUAMy4AeXwEJhw++5g+aRRPZYryaSNWVMabZ64SxSyBA6DWdp3dpQOozA8Y3HJuq
5Hqc9C5fD6Svm5+Y+wDC2f7m+G+9kbzVzQBBWeqQWZKE/Fwy8uWmzk/t+q8i2vEu
VGFcyEuDZhvUxZKV++OLU7aSOtMu0qYyB/1Tgo+oYuwZu2ztV39K6kvLyQv83eI/
40N5KzOVRZVB9zvDEyfNIDtUxtLf9bIhcWljYohXGHzhqhyOqHnzDWI6ZVGfdF7g
dYWkJLV8C59N67NjpWwRFkCPu5GKxucaQOlqCd+kMnyh1e0YVajk1Mqo+3cRZimx
fFpBWdrsp4f2y6JZI/nusyD2oF0tD4YLvO2G2Yb/Aculo1Ky0IaEofmseo3A0GXh
2YQWaino6wJSfhaTPG3ki1ut9nCCvg+yidqWE9YpTOtLhfDDzd1TzpnCi/lBhSBr
9JTV0g6atzOKEtA9HboO+gaasg3ISRbVRhqW0Fl8nDVfjNTIvf/+YDjx3WHkg+Ec
acpfgGrA+1lpq4hQEmzLTFJzaxrpsMxthtK107eQXZ4wX3RJ0pE2Qb23vEGY1QT0
UPM4q22xMGh/0wO3szqKWUeiwwHLgrM0XkN32qOhni/M31olvgGB2PvoqS2pUfDf
yqgc66mtVAEDSHNxEcRKkoa+ZMtLJehlDRdGylN4tbBRNOkpDWY8Ze2Q1vA8b5Wu
/1kUJD5U1o26USLu401UCEAsYvBCYnnhMX0ST9DOBm5w0HkPs+M9Jnd4oOcwJcow
V9rg2lN993rlIN0OvWjAN2rYMaw7IY34OgHufkAmUan7yH6YXiwCRhT+K+0YvnZ9
5zBZj5ZcKt55c9J0H4d5cUcdH2dHNBCPKMqEJ3vJ3imUcl56iS1GmlD/1/d56T4R
sFsI82AdaNl9YJhKECjVy3yFE2teHlpOq1yV08tHF5MbRcqKf5T2SmojcowAxAoF
+W6BwUb3ZxMdTS82pXaxAsjyUXYud0n3i/UxERcgV3yGPIRdKl0DA4Mno8fdYfqe
rN5h2L3+z0CFwbi+UdNUqrhnzUQUqoPwlub1AhMh6YYLTNytEl8+E1nlEUxMSx3t
GKc8cCdc9bWJx+BeOTM47thc7jIl0WIlWAAcdVKDXQexM/4Q9Dh5i06Rkxx67yy1
dPw0oxWcudDEQmZxrL9jjSu4sZsAzDSL6flWY33q51SHdCuElal9ePNWmFmN7K5z
QvMjrwwaKC+Ag1ChBATQ5vEYwN4FC0pmvlSq3hyXU8dW/6BF50CKc/AoNDXwQQiT
PtG0zNkHvZszi5HSrDZ+tZg3QnyMiTndOGinB4TkVoY6vFzAWaMROOYQhPOvkYic
IDT6OCbdA5+A7XNQxlcAqGbVNPQSZa/AIecdQvlsqAzpMp2SvNsvL12T6cPXFVKN
S9on92R0BijIKHt8p/c8M/5tjDsvBV9+wjmTFloJclSM/7Zg9S1J9FcppXbZXI/N
y5cx++f3ZcN2PkjgMvf4LRNt1dR1YAIr746ONLrovqZaRtGMCVRZB7TlSVXQB1yH
cf12G+8gp+vJndR/YQ8EW4gcNQzFUS86FAp03vCpMXDwzls9dm6f6uTDtQxG7dIS
VncK2Xsm5oL5XC1454avo4ZbiHvNSaZ1sXN4rfUzW3j78aafdt3OWmmKg7UTqgLO
U+J/tKWibeZpXWXSPk4q/g4W4Cjf3MbQey3kREMXWQYEdTswMdpTZBHF55kX7WZi
4ro4Xir7z245GSxsrTzutIBpxkAjEZb1RWYDunkbVswxphPNoBqoMJ4DgR18Lrma
ipT26MGJ0pf8uO79qgBECTBC0jlI3drb1f/uOcB/Ru11soI7mkcX+lseZz8pHz0I
5rblqYcNU7oY4YsENyE0rKLTe9cixS5QUidZaHaMsFrXt4VFNOkw2/IBbMZkltxk
XV1gXCoxi8Hs2DxgqWvNP6BC7zA53Khkwc3QcrP55Xqccy2eeKc0HigNa7ieS2Ct
0rdItL9n/ZArm4QHosWotPKMKT4kZrzYihkI+QY0EQNcR90yQ0Qhh72NAIdRSlHd
iFDu4wzioq8QjQsZyC0hDFBG+x2sHxlaxgWU+zRpAaNt8bk13dM5Q8Tl8vA/XZkn
QOJZbc7mNK+WL3D88jeqgS3X/AyRtXpuvXPQJkV8LjVSXNiVQcw8LR2sv85UcmTI
A6iDWgZo8CWll/H4i/Y2cSN5rSKDIRe/zuGHTEKM58RDlQfzZgC+jjJnkmvziHfc
J2lxidfn+cYHHDPrvO5wMkEMRUgewv6wmRpbh4uPoyxwMdwXP+wDcVYKXxemdMP8
cHnwigQQQlBWDnvbJEyu5S4NhqRxtcgQNj5uOyQBdovBE80TkNDX087cXqTirIfw
+u3XHxiSC6PJIR1KBmoKjDlREXgScUQqWi+0V0feveVKMxPSkGX5qA/GUWtbaM/K
xbUaTY6KywwRJbeUboE6hMVYebM6tX7rQRs+awEC3j7DdhPSXvg15srOXZXHzyCv
Ivl8nV2s5lzVneqSNg9tvqCQNQ5m/bh4vPUU98BaniWx47jBH6hGrvYqSuooK2HF
3g5rTuEPMkG1NWFk/TcG+xsd6Rl1iEP4JeWxN6HeiMcyyFBa09m5G7tqLkqBH2qm
tAuTDB8Nngng9Ed5oL8JJnevzUjqCpDy/dzAnyllE+Q3lVxGTvok0RfMTvacnYDV
4+R7v+JCYoe9VyUuePqkHz3GryG6OueLW+x+GvkmNaM4GwZP3wgbu4oOJ2YewdDw
x5UvatVHuoo0qPAKwaBarZEpTEiAXQi6wfHA/ObdiK1GwGRk6w/DfVBTzfH6Aklj
vMeKPz7R4BpxiU0psr4J0KFISyQXcQmu7LqAAnoAFqCHY3IBV3FvRtAC2FFGzeHt
FucE4QUyELdWkMZjT8tNWPcyKVfAO9FcKm+tn5/VxHqbOYd0l9VpJ78dVnPIeMry
4/JSkh9hyupWc+y2Nn5xuD7WeXaD1lo/M7Ji2n9ywrXYeGIqoPCvsyWX0MV+9N0q
4K84RDtVbN4KxfiaGpYt4nLGNBnMKsgvXql53VYpaU3Fpk/hujP5E4jBCgFZ4rr4
2zEAIiXfYEhZucxcX5K5h3unjyTDYuYdPTNIWnHGT94/4dkGabqLDsy8yI56ZFOo
Zyakr44QsuN55rSC5shbRMrrUa2vFr/4ubLIO/O6AhuH0i+iY8OHGJG2WqvUWXDm
kIIdUjwjtUYQA1PdLdQ//WAXvv+i3dnMhEYsYTONLuuovZbIa1vHSWdWUGerUjen
KQMTZK2DlmfVvf6EJXDNxAwghuGVvQynXjPkdkCDqf6S4a3ebBvJGKuyeArJfQWs
RiM7zQpq/+dvp69p10eOvDGDcm2UvRnzGkyqAUors01tBHt4Y2C43arCrVQVYO7u
DeFxdVQYEfVaARO6frv7Pncw4qYep019nGxtCdyo+5tMxst4Bvk09OFQplh3Uovb
0y99Je/bdHuT2kGBoeebKeJSe45wD+r+4uYUczBuWa/7urhiBeZf87nxTQxqCetY
O+BIB5Qwm2wqcdDElg0aUf9uji83asK4ir4awplza6El11uUffhu0HW3CFDJUeVA
onkqKCFV7Z4rK1DPJgsUyvg1l0k8/rDEhNCW7QCqsYCxOUmRz/6yRrQuBJKE8ck2
0n+dr6Uiff8K2CNEDolGF5nWJ+29eD5rVGBvJvhUFmwx/ka+dYei722XGAOZBCh1
g3VWu1tYc7tuoNJmQjVFl11drUY8cBRZq6fhZ49VmjMmFscTVX9PpPw6OweN9wfr
8sRJz59wCArVqKzdC4MVz/bjBR0rJYSEZvdwnv66H5NqecBTr9SzhJSbyDD/wnRL
anTDBYp4rdSluUuBqDsxKUv0H/T5FCLz0FjWxwtm7awE8VdJPCbjuPEYnVVhf4RF
EdgxRMk0UxQwmLZjUXvQy9dOtMXpbBy0ZehIGQ3AqRaHh1yi8NTC2aQ9IpJvPHv/
6MLxzmgbJqEc8D5BMVOhvsnbrBCBEMkxz3Q/m6f+EVg0mw9btxR7ej1gZDQ5wIJN
g4B71FxNBoKWOQ6lZlcPuTX+3IPsLa094OrbaOi0BGw7g1+5y6PZMQ031W/X7gMs
KmU/qjHCTyuJQk14cZyoaECf3fZnLliaYepW2nJgnmFO854L20IhQa07Dawbdzqd
WLn6uNE0jNlvw6VcwH8cURig2D9UxNwa9bFN+JmP2MFCxIUa0I4XzL8oVQyeT2VN
RV+K7q7CpksY18aDi3iOwLiVSv6RGqhoTL8erQPPZAKl51yd0aJndy/s3KUmpFA6
wPk1HLmOYCmPIqOSbNGoLKltMEWFMdPIBnbAhLNCynnaIqFfbm6IXo1BTWIkb8/E
cLLbLgdzP957jG4OMIu97h4uGpuZSifKYJnKI6n0ASAWrx9BPs3c2AhVFCJPHdBV
VcdPZ375YPwdotYYB7RJ4DyHVRZtIz1N2pjvZfM0Zo2diGG9hsP511N0N4hWDASc
MoR9mDaS3GIzuby6gR5NW/mYwtPlv3Xz4PWvHj4QFRlIJJol+GonkASZ/k/Suc58
+CW6/Nqp/iy8nWch4LhrwQHLBMv0K/SPFxpzCXDi6QCW/4JgGXloW8FU8VW26pad
gInj0PcIDpD8fb4VairlExJz4Q3dKfvvQgNHx2zLvyb9oBaWLLDFQVBEYWAodwus
hXnvOWy80kJ0+qFSFvDYQZ1NgIwOkj88ai2I+0aISIJx0WWwb1K0DGXhZuS4KIAx
oBKNRL7iTjQXsUJTiG5zvdY132qmdL2KSqGu/q8wbKaKlfJv/vL2NpGFp4xDWnHW
cuhQO8XxnC+ZFTcnRB8R8offAT9NlwfEpWUItXOAytVH/sxZdMBIOIqGExDooWXp
C7s0Wto+1qNLj73lg+RMnzWuRheprhYv66P95flEE/QQFY7dEMisi5eXJok95QiY
4JT3kMd/wJADpnGVoJdactqGd/HtPnWQjgHnZiNEvL4sxoPSRTf7gpqY3JPF1hI1
zgV2Nrm0fNIXbH0PcgFWDbf2rxlGzpRO3aMTDrHmNKbIB5x9F7Zyf15nGHli7UdD
kws9mgE/+YRa1NTMR1eqtcCviYufHOv/rNLO9XKJP1iclgdH67u8duEpapMCIlNh
gIFWT/xUiDOMTMKfnL55vSylzQBbYqcGZAm9Kfl1ozjvWNm7jNY9XMwhmYW7nehX
pwym6+bbSSun/CdbcR45uywA2SyxFh0I6i5FJZl8o0V+kxR1pklz1rAO1bcoWSxF
wW4BXqkP0StxlOeQ9+215qtPJAu7RwCGp1HsYwXlRd13t68Fs9VVwp0eQeRo/sab
VcCWJbHseIfWuNb9shn1f5P9kLFm9UP04d54lUM6LFD7wJycJpomZm9BWJcnBLyo
WKXqD4KYT0UAAeAX5tFS6XQZiwgs56P0Fvoj7uuEFIJqdNQcC0RnH9mNflMdqIji
NVfMxAPg/IvmrY8SVbQ3SfF2sfaIv7Ca+7cb/50K95ekVD/kmhIpEAzCDrNDZMjT
SvTezaFA9ZYOWnF75c4K6QLyFD8LRJcrvToZQ6NseiFPZyASyl+PVVmmoO+2LHGR
RldkHbxLEY6P9Er5AUjUxvfCsJWpA1X39O9zbfVxvAO0GFocmf7dipINf/FMp2FS
6GGekIDItUquwYgqEf1Q3oWr6hlAMDz3U/4hlCza560013zvEuRbBk/0y3oS2oEM
2FLmZoSJSFD9+dZOgu1Eru5kETDT6foDfO96M8+QbkMX0Vdr8QrWCLRG82QVWElD
0P5pCxVBIaroCMFpsz+EmB4uDIYXfZBxArSqh3CDBb7jyzbcpLtvtMYVEybyXOLT
n0ZbH8AXDspTlXjPiK5n7qIiQ7Ux2JFCXQcO8KM7RqatN4CnP6N8tNRpREvNZgoq
VoU2GXXi0qoUL3xWnfslGL96Ax8yAbjnuWbuZVetNvOIWV6kqJMQ7aRZALRxN9d0
XgwkdnT+R0ZC6cTZ31JSB8p13R9fFAHdtFbw87VqjAZKoiXBR7BCXSmZt2HsJcb2
X7IEvK/Mv1YiqsgtBiaH8y15fbhhaJubbCyrDCIaYI+dcesMOfKtcTtIAeqkU2nF
HW1BtAkwIqryQHPt15SX6PYtYbc2yg07+AP4oHnP9TXoWC6OVvp0QukIIMZ1j9En
vKIlMypX+lVxnxVxnA0/atdMaqOSBbdK7Xtg1LP1LS6Ol8a9x/G4D7Q4BeLoiVlQ
5yDALcYJhDEhUKt+Mb1JTco8700QTNBPC1t927/l10aQOGktWxrJFIeTlFyWp08F
AEktZ1lGRaYj3M3CZGXOdxz12Xu8z7iTgwY69ei5iRzbBNSJdrM3+2JA1V9LYxPY
89EFJ0kcOZCiOVhCu5RNiF3g0vrOItTHnLHbk5S1puMEwyXimzvLymbriT06mCYr
qVyPpKoez+pcdKw16Fmed0xzCvenm/cACOZ6UgkPv75rk+IEMNwRM6sa+6EBAXVA
ecQuiU2QxHNIprpI5j9OtiMz4dWohETsVkS2moStdRvV8Jd8b+5qNaxGpsPRgIvt
Fcsn679wWSF2+8JHnBOfo6OgX33oZ5gkOoxUOPX2oPUDVHywBr2/bZ76X2avhPqT
QjxKu5qqca2sszUWR0xoOtM4wURegTBex7t83mR58VGHSPDlYKVjuDdtve/1ClCc
9cjfjsAaj5aGY3TXWVZJqDz3q21NMUnH1RvrMz3COJYmZ57oMvvqrlvRWbGVJhdB
PUQK4EoAlxKyn9OsKwFkMm3sysF6VV4q6dDLhWR2TxKF3I77IpJYhFZIstDtD63r
f6VHM12DrCSulDlHyTd4+RN/Syo7DddFmClN0RUURfr9yQ9uch1bcEHJ4ENhsoMy
7pw/It31qpp4wWXMLW93FvPYF7xFC9n7IWNvRa64CKwV7i1+gbExF6XIuNw0nYbC
KIXAu6A9s9GsKiGO12q2Xhx/TaW+i+gaeceSpDcJkpx/2Tx6CQX4lbHIs9V9KmV2
/9x6oh0jEUnpz2fj81HBDRHyNcHOs53Rmf+gj0COLh7zopDIyrRF6RfAqkNSjIYR
JdjksgB0nsh2WWmAY0Cmy1Pi8Q92xBXRRFJKlMz+ECleMlkTxwJ9oSKLZ8jzXOwJ
oHyzbA7PqBpJ+bwPQWcKYKn/A2lw4i6woD3ZG62uEXaHEZCzJo2eqyAe8nH/gnrK
RSHLZu9ps3jCGrfLOJKr2Ar0hlEKnMe0BnNI4yD0FfKi7LD+YczgIHPprvrW6tSW
3/XHnSp5ex3eakXlE8nOjgi4pi+YGAP9cdXw7MGLxLGULY8lgJp/xFXxpzaE4ecB
c5vcKSQ9Dm4LLocgfuxhUAdj3yhQrQ9tsHaaq91OkbezB0uOh3CP1ixboJanDpDl
8nXo478twjNrBPsKfGfHda8rnbQd9mkOIlZm4b5hGb3jxqoBu7f/boLmvGczCUBq
htukO7wrrXExBejUHRbrBoKEkBs6EGfDXsCyBhwtBmjjmEkFN4ypU/nri147f/9T
76bMz7U3NDcamoZYoMxG/0BHVloJ8md3B49pbSxAsRrPNyjA1qoOmAEINwwBz0gO
P8NDR15dz35I2ICivBywrOMknN1zPmlktQrD1oMBTHlir+PyUbsj0JhiQINwf7sO
vSbIA5HytGITYjEL/4EvpGdvM28F7QL7kRlHQfW33V59lZWn0aGylXciQ0jkaBiY
yTeBRkgWcQT+ZyNQ6onkaAr+ei51/Pb1AF3JSJJMgLjn80bXzvLpIsZUva+ebadM
fa72/IW7V6rPuPJlynxN76MAUVIEngKMeOI8KMOKPYG+92STPFJTQfE8exNNSnIH
XCw4v7pEGMsyh9DI3OrSJX0Y07zTBLHn9EWhVzS29CRP/0bpyHrCmFbfoSVKhlTO
XRynRX3zsMFMjPmHf80lVIYUFi6Px0Qe8X2oxyNwPTVAmxo9dBblilCy/4glg+4U
ky2Piy+QJswdmFV90Ityfv796Vc1No5U59DwrmPTvi0RN+U0NdI+htEtiUJ+ld0Q
m+QayeBToZZLBdQzCTcY/LYZH3Bim/EyA7cIEgzCTkkSKLQpd7CokN+Lth/L/HqM
FtC2s0HRA+C/n6ksevgjtZgm0JH4o1uNA6y99u91mFo27zaxuJYZwLX7lrxN1h32
eVfDBEfkvx+BmM/gL/VBAWKKOKqzhlwTIpEv8asgVu1y6xySrLv3JtXQba/3l/Ct
QX67yMVe6tnSscN2DOtLVsvLCRRsqU+fwte0Z+e9cBCulrzzNznAc1RM8JhTlr4C
uSJeejJVuTE8oRhDRJwtyGBnewOrhz6ABlWaej9rdJdF0ICWQes0WV1W23Ct+xXp
LOonXOloEalbTLKivJmzCiura2Y6uiQfg3MwaEFHNCr68mfmyORVb5MCbbrv13RL
AxtbGnTSHp9SvrLoUHBGlxowHgkOuV6k1t1vP8GHI19avBd7Ya+8++//9zKQxXWR
XiI+C3ueN8QW+V1TKzSFw6S07wYcOLqfAHzSPvQ6lZ02UOKiKZWbbqreSUoTfP9u
xSkYg6hfSaIWHXmLTxUdeZoZ1g0M5BeH5v2/6X2HYVoyb5OQ90QBCuRhuP+1N7vl
b5AmnjlS6HEImIBQlv5SN+KTMBEM+oTfuj/3LCwg+16eqnwEQA8n3H53a83GG+VV
i2rRmPal1/6MjNp1N53ZrvbDw9JYOHgX0ngdCS89GV337Ejgr7o/X+AbDkPpOR8G
/nnAt6nuW/SCXCO/Ao2HwyF/IU9n13WIdeChWjaoGUgZHF+HWdelkAQw8/wLg42c
sRq5ePr215x0eT3oBZNQowADRERuKp1UUJ3NBmVryALO7y5+MsdM3OAWtCmEkMtK
ttzqlQbZhM1ItOUqj0yEgglz6lpPydbmfHNmDwP7Rx9SUkx4FUYA52dXSRTkbnfn
BW8xhc+RBzFTrH4So+6seulxidaxV+6jHLHqBPcYFMOEh8L0mz9PeHT1W0Cby9ST
MvMmZZ2UcbAKmMN+PiC0iVj9I4AJRg31ubacLm9Kz7RzMN0SEozV9esWHJ7ezrcw
IA/AvyCwLrJItPtSAKpD924XKePJBRPzo+Y3dLXc/V2P+b0M5FpU3gMLCFAP+I2J
qKpRfu1eugEWXmJzMwUTxVVZbX7UJJgCJS0E4A2fCEM2Up8UIYSpBt4w9x8hqBpl
Vh9vhITMsgR1IueXpuHvJsdfQXRE3q7wY/6QVkpziNUtlVZdyXs0Gay4X33AR/1u
MDDzOsCOScAlLKxFdiErCvr0E+cZ6r+sA+nIjx88vFPPfmbMxzXf18PsFf6kuRqq
MK3Gjqrr2P8htfa2vRPxad8iGxb7IgZS7WsGOZFBw7Om3nRff007vz0Ls3+2b4ZO
gGznaEbWBklj2fDmXxIHQZ+WfpEb5pFnyZRS8I3u4dsiqYmZffiP/I43EGdDrEaV
5M4J0bLE7t9i/1i1PbKlL8iEvlbGPIEFXU7OYI524iQmqq1TH1zbKauquOQT9Oer
oaMWMcxOp+6Lvg3ij7lLqeu8AMLpovBY/XEwPOtYgODq05QyjzZ2yAjEVUHmOy99
Ws6bFned8kEuUNlx9w9M5aIQArnK4mkqxmqOAqDcRurr+5eTzyqL0hp6C0oFmFTw
TpbnbIbOMptseSgoDAspKu/FZy7AB8BY2nkx/XkIaxw22fO6bhLlc3oPo6sqqg2U
TaZE2m8VfQhlIq/dr8VR83Pky9duWDZZGh+eUCeF7fWT/TqWgp/167BL4b8HY8oh
siwJR/5PJdLbiumXX9VSJVO1LzTD+YFqUkQjOdNPxXAfygk4ixwZexfLSxlXjMQK
f/fx4A0hOIFoZ1p+wcAq5bHCuSfbLEINpTMK6cYQ/Goqn+MblUhtcQTQlCFYddQr
6jXZ8fI3gT2yhpZWAes9fOFZpe3i6ISVHXKNRR3eaMZQCgsvIeOp0eb3axxqc5hq
+mRQLPeei4am4kMUh7DhH3YEtCfr1damSLel3P1OJ2wSPCmg9ui2gn5xBh7LMVMZ
9mzCjLlFHJloK2xdsphV21rl1KupbvbPfbUCpcyRseSohCQwlM7evL165uXbpcXh
/YzZ3FLFZxY7yRPCGLXnPnTHCxWDEbUv+YXH6kTI6ycm2yNZDC0TV4s7E2AgTLCK
Qmj61XpZp7kRM9uBkeBIO6G4UUWOm+ZgPGYPiYFifw0uiTmmkxIuJuqUgNZD6Vpa
WF01XVk6PXXRZShewpfJpr1kK0CuRmxBqREoyD/gZ1hAE8FMfK0C5K7EqVssJKe7
wFdHKwe/R0zXz0YskFxLjpZ+ecPX767VnoxPtpbvnXZoU1oc2g7LNDN2Kd6rI3Dy
KW0sbtf2HbPhReINtCBPmGQoj9aKzk0lGHQ2InlNHd82vHc+FnwcExW0yrFWd1Za
iK/YqGXtajHM3Zf5v0wmc0sQ+DzfFoilC7JGfxmdxKulxSYBCsk1R1r9pEDie5VW
IShhtup0w+MCloL4iJ7picXEPzMT5c71zLaFE/Hpcw9pUB6rJ4HlKKSSBnJTjiCo
TajM35mKL/l0gpbsVNmyJGcGoaqEH9odXKtAGCfRKZ85CyrSxVEyMKwTviGuocuI
3XvpWil1KuQtWSyMRIrXD73HFiKlQj55j0DRPUomtfspaxQGbkHlg3Ti7szcsl0l
o2o7A4ZhcayQL8sxwDBh11YnvnQGoVBoHjZ3GvDQkLUd1vbFIIUHHAyB//aCwBYa
HieS4oEDZQdKy7knWhOAc1W1lEFWSrcCF+bMTdNM/yPe8cMRQK1MW012k6ZJqE2L
pidm8yR85tecFKk1OZ/RgC8IYOSXFo9GPLJd1oiuvo4Gk+KHCrUKdUw5lLkaG6HO
G6vPFUiffXeFE/SPG85fg9lpGDpjOw1I5TslUGHh4l6+iMwcww/R43tJCWDnp4iL
QOLooOg/ijZzsYx3yZXraWS++cvTAVeRXzTOOOuWwAHSxLqVQX5bsoOh7ZSIO74J
OXqKmHWJt8Dvq9NL8tchCTUzcqBJgULfsiYnFzZmE1wLWXrKxc9AqET7kqRAs7rT
pC0i+sQ0O5g/tmBQEdnIlPl6NcIfIa+hxkbepilRlUg02nsgUh03th5QqIgphTRr
wVRq3HZuoENEoLLrsbkXpxlWx8NK8Ow7lw/WHUnTBb9v0jPeVXHE3FLKBCtWEgOM
d86IykzHspdKGZIYya0q5AWYjDLIOx2gJCjwh6a2hxomtNsJwIyLfH3h3Z+E9nO2
YEvkWTJqMNAiMddwYyeB5AK3Ok6tSIN+QLorR1uXT7NiIBpnPkuz6EnG3NUKWGQq
YLeDvEWp8IlmvnSRb4O/EErfM9BXONvAZB03wRBqzOiOm3Jjn9KT3qntOX5zeWcT
t3ga8ARUDSyXbEC+xa1fWADvF/B85vpN/KROxxhaKp8TrrAsmBQs8CxBLMgHH372
4XVW3aBAIIetLG6SK5Usb+yMuA4nEqojfc6qyjmdVOYcwTC3PqMym1JU7xovDE+j
czvJJa19INSH0DHFqzXDuQSQPb6OK/cLtZGUtKy6E43I0TWoQczksOe4H0b2Jk8g
EXrsxp66F8tGOQJffUeRl+9M9CKfi50M71v4x3LzzvQdJkBMRE59VQay2oe+5MRS
h8kQDPocqZtW46tVk3h7RzL3Qz/s9FzaH+8DPHpbXcd1VpZVp5cPuigzfepW83jj
aDf+1wfHV1VvZFOrJIXf5IpEC3gl965V+5EoytJErQ9aonml3VuopZMwDMLrVPhZ
IzTR1DAIjHm632r6jcC4iiX7gpb1GhKkUIwILTChX7v0+Wswnwa2b/lZCpAvtnCw
3sTunHzURQMzdnNevTu+6cjykWA7tRYyjAODLqaB309x7JJxidnIrP+n3tF/HGuF
tKLGQGJ3Ia1mzVUIdqtZDJPc+ymMKEMd6+l3RZR5gMGTR0YvlAW3P47n1m+59tAC
tMcvqQV09732SL7Ri3OABJCm3+ZMpJyNbtNCIkxNFHlV3UvikylUppHFTBfKN9ot
TMogkyAUc/XFkm8SeHkp7z+LO7Lng6PkHL8UaaK3sFB56RG4n2gIrff/N78QtebZ
RbEmoMN3BrCrXmwVUCvdxlfRVCR9itDTkA673JOBn9g7JCxqtUNCONq5ZGFjKI1j
1zmRl2OoZLmS2tWzC3hFnoAk7PcsM+aSihPgsZEaq7r1WKnHrmIj6pePSzcTuwqB
cy2t2oz5gXaoQeFzpIE2FMa12jvlC4IAO8aXbmcDe2EmXsDnusIkpipxU7biNqN5
PIA8x1x64d3CVfJcYLWdwpVr8io0LU9LVCXHt5dH9XqmGVD2qnmGbL/nIQ8aCC6g
18lRQ714PwvMdMsIfMayihBl0OlLYfEtRp0LCxVBDCzS/xlHenuNTeC0Sn3frJrh
/EsWQX7g3VwTzTWf9BMEM/9LXLK0xxPadwMTMpmWlvjjlBKhWLxZDTYZYHT93arY
QyrTOiEg2mJ3mjlBa7Mwer5kgWjQa9bblHnbGYVmnYTpWQ4/rKxooW5adDuRTTrJ
J0aFBu7UHS/fjsFUSy6Zd9jXpIY6PTmWZGKwc7R4/FUQEGLoMrJa4ly4jzyCvTjY
FvKa/Kjkm23M7FDB66IeQopUtUea8UP0cfX3JM9KYDmCwFfLLtF9U4vYXeu/O29u
FhN1AmEz1whGbBgRegjawwHZSc1uHZGgNmY2Ff+zjuDPD6QGYYi56lzJwj1+X9/L
GiQ7cF5dMc6Jcp4qG65XunBM8DBHL0SOF4c9BPqBXzhB87k/btFtRgnkvKfwjnyk
5oRVWUKD05RSpf3rSfwBg0kQ6ek3BxrtPpbWVKimESW/CVRAVfd1nbKzbn5bhxQH
XfhNy914P13z9GAb/MOFg9FAu5uZj8G/t14NIhOBej96Ud6+UtJnuiHuABuF2XhG
wY7OrwHnVx2ySm6EMiTP9aM2B7LvMl4YzTV/AX9jFVBcLBKT8DWoicahk+XK6IWA
+NzdmhD7qtyzye106P0w1EBjLc7wI/gIF5r3b3w+E2DayMiw2DAp69Jom3uUQ6Fc
GfM7Fdla/KiVl5BjnSlAa11/iEuf9Ycdmwhcyh0DhOpwEkG3sMIIz9F0RbVessLD
fQ0SdxQ/u82iIN4xetNVB15iWPRSewBNtp1bGJStWiY934LYpL9GdnTJuGjs4SNA
Rd7WyAIEeFUHdRjoKmOomPuuzjpZqMKa3az0OFQ5RDN/aTW9m3AFJ+cRMcpSj8Ng
lwSN60WXtZrwO+JFrQMmyGwBquFzuDtIiGDsAnB9iKJpDm/NaGL5YPOIQmwTZ7ek
lmvaQ3izpc0Y6/LCSjwrnFwUkHdEBCYMBCTz437GBV2o5/7tzLdiHmQ0Q1iXrPnV
12Hr6MOL4VOU//9IE8FHFrs0EluPa9fS4GY6svhBgK8dqtHkLXOk8syMOkT4cuhP
h/XSLqEhCsh/QziHz5v0rl1rkc59uyMsxXG6UnD8C6IYdm3lZBfiBuqOND8QsO/N
yOoUQ/bH3QKX/BbsrKRufMKZh9AThIR7+NstRgknGehmZjpNIKpXa7jA5acjOz8B
nd3m4cROdKdEcXBztT/X4c7zFcznlI1ot9kjggVEDZZuFpoIMSKrktifwFPhhvlx
lBwChsjgbZ4kuZgeGov/bnm4CcAYizEAGXuvB5FE1EILsrfCCm+9RYot8tNOyBmP
vFhOQDa/fQX3/Fw4iEIRJLmjPsrYBzoZKv99yRV1bKhcvzh4tahGP5qpe8i0yD/L
eAergGwG/8jzHu7mc6cfXx54hRbkZ3bwH7crjXdJ+l8hiN3ZO/YhUihMjYHkkFh/
lBX37zz1md7HdaQGoLNdyYOlmNUNVqPoheIjKihOxynqIuQ5hUTQFXvVUdQnMzsu
RmH1mCKtCC8y9gVU+CmLpE5aTkGL7hnha4ShCEVu+i9gVFeEDhHIftE/ujNHsQRy
Fw4ArhIMEEwypytwmujGlMNeqdItZqhDrQr8m1bGv7f4EL9O1ur0pkGRSqoy3Vsl
l9eCh2xFNx5S7b9S1GVDvWmZyWADbIeg+xmV32vt3GcQKBemnTe5Tv7szJb4/m4p
vbU6ZPucrLpTLD8R546XmvTJazSeaIsDoIDlBtUO/In9OB9TKWpTwRUmNEzqtIYV
pipPIm9Myqx8PxTruwotIQ6KNdHAhDOeppv2hIQrq28TTiD21oVEyNvS3lt5k5C8
K5JaC5d42DgKHHt/ZQfHQamJtPXnLZeymMDPlHSwQIj0xx6GkuLZK/v5ANvSU8wP
1QLHdGwzM5BxfHckvHXx8F2aC4LvJ9grfraOx+s6sIwC/ZwpflVMtY9HyKAnscks
zZsmfJfTaq4vzKMgZJptCUpt4BvqNox5R/3ZzqL++4/f+WYFj1OR/rAMavF4wdEX
+YKolBaFUh/A2CcugwqG4xMHB+ymmNdxb6UA2AtoS/waQuBcYtirWFcpdKokgA2m
YK0Dl2Eg+toWeX9+sbirmDlJJh18L91rztCk3nT1U3oGAF5KdWmqhoWyxrEatmJk
6lWCZuew2wdF3YlhQP3HFHIxSgHiGYHEc9YyTAqDVh+REWrskyx6O04emPGwEsnc
WmS81BqAfD6zW+/EI2kgN8TtnxO9dxweUsevwmCN410VA2DP+2tMaitLJ6HBLXOf
p/Pm3o/MA/qTH5/1s+c9Hdmkwq7QvoVYGMtuiMpcH+KcIYb+tL4ncjsA9+HHlLRQ
N2z6Zd30kH5H0Op6ISkfx3/8vqdZpwGMrlwoFZrS2RdznsqcWPzo2bbpuUTBfqyu
R/tW9mQJkAmDFMz2sngQc8FkM046Sf+cu6umqSjQfzapYetd1Kb0zCjI/1aDuihH
8NR4lLVKu1GMJUFG9e7JRhtzWU+OdDBd43ffJGY9b/L2pdADhLiCbOgpsziRPi8S
m42FFLDkF0ntb9fGrHIlcq6tUcn5ELwsBHd4HZydWpMc8Gs07zegWqK1cR7TkaGj
XNfaeJnAS/QXf7kLuU9wDkls3nnCVRxl4IeKyjHjBo1xQOvYGoobZHtE9a9ZUyVh
aDLOoz9n8O98iP6FFIyZx3aBIRAE2DkI+YhIH+TZPD6vPKiIqdOaKpieXnq+86wP
eEB95xAGJ+HuOTbegdN8O9RI/FwG1HAHPmxXww7lxyqlopftc9h3xvKZFYztFt7k
nL/9uHxTuLvlsn1oUdW4Gawg+8SIk8sRgph2emq+lADfpy5KTJFhpRg0T3EBABP0
oDqiKSqMVaGGjIfW1CXxCFgtu0khBRq5AE/neF8urA15y+nU39OxEi1OtCyIHayk
vJ8nfEwwj5I2VXGICCChoOGoKs9Egpqt0g7qe4Irm2c6cEysAAePpeMH4CUvkOyi
/GvCJCfOw+yHKx/Q9Vl5x34Rmbaa5KrY87/7+jMWbQDff0OksAPMFR1ftJcMM1gY
kIIaB0o8BfBORewrRR8M0uYULBywezMj5an54OBaiFCcJvDniCQ+PDn5PUydvOGV
GF0/I1uCSbwy4qgE69p6W78ggDIBudgYU42rFzbt9gEXReL4pKrNYVgIk3xnf6jH
szN+WRcDtES08zfLCtseSVJR1MXCgg1mmhhv1qHiikrFDOZ7xge++uXxlKyoiRLw
j3G5RrUaYnphwArk2tcBnQRaC94RChL077k8qFFUt5Ua0Z4RPFp3pmjF0IBhNMLy
c6iqEJiz9lq5PKkxWGu8xRP7zIkVYxkhxUdK8M4J/wwdZISR8+y0dtjOvUcM1AM1
9dvQ13vxJwC4KkRqKoydR+Gn1v7WoS18ov4kR5I28wOIBGHZ4ZmUAzXidcavDYX8
9ZPD5YGRP3uO+2cTLhOaTb68mu5XWY9dyZCzrYkhC/HODsKDsImS6cV+sFeH6DW2
oQ3Xtn7aa4gXMWnY9uLYHiUv2BAtlkOarTEHgNrt0fLVoI/oBf8sRkonUS/MNn6d
6VyzGD3/y6jdtIuJGgQ4JVWyQui3FTtHe5tBeBtKuFhqiaP9I/HuhaC4cidgCc9i
Ibg9Q38OtH8hangfq2tDPvx7UqCkpoK7ZTO5+IA/xNgqqcZLw9+ftQreTCen6/UC
ItsUtQutgL78LWeNDk/vxJTTaYOwqPY6ppkevsfeXWH9pywDArcFVwQWGqdrs2gF
22+Z6VhKD1VfCUXLa1gxhXVj290q585K5RWu4o3LCL5Iw7P44XQLHuVAtmf7/uUf
WtpzsqOdp19PVH1hXdqBWRpO4B6VgiyJ2enTRSTj+5SVdxduxcNYTzLbLKGlCrp8
RtTnaiQdD9tDweuIVj6xbSHr8N5tT8rJjdjCQmeEilq1yimWtRfOh6xllilo3xY6
dsbB4M3A38vdbk8ops8OKTX4Uc0n/hMJrcmDIrkJZV2XeWMHeOrJu9HNAg5NXxWz
81/acIgs44RXmnMqjol0K+0KU3sumcKz+rv735ARHMD0akLl9Nxszc056JgtU6TR
K5NjgB5fWvIACxLkm8qwA/WEDEmYrGeCb+dtEJuv7l/2Uf1cMSyqcEqexJ5X8pfJ
OTVSkhP7+Md6qh00R1exdlsb3dktNK9++gDwVbDuH9827QKrmV7AEyCecRU9A0b9
5NXQqPDv/gtM1BZ5CNvVcf59ucnUDBsTr4UBAtM9yJekemCZzqsRjawqxPqFxH3C
fDXClqUVaw208Ai+WmjB8zUtlel7jxvuipPK6flom5yS52H65jm4w97fclQnP0j8
U9wHVCv4bXh8ZUVZSwXPyjwEHoG/J5OBWVQQvwvDRRCc096aSWSwR7N7JH72C6Xp
oH9xH2bfq/W7bEMcAz45LSoEsGgx2nTOHPsYTO3DvPGfYIvIRViyd4IoYoJA2NfJ
l9SzOO5KXxILngtG3qbcf/5XzAcPnVP2QcaE0nDiEeaqX7LQ/VfNRiLiY8U6DdJE
KmlfWSa2QyTvC+4uPbAaAcArP1iwt1A5pqSQFvjKt89oYlMhOdm59xt0HBJOhf3j
0w7jQd7I7EWYETpKnApxqCIuCRsUqX01y+rzbINB5f0cqVKujbV6g8KCQeMzwWBj
klVyUXYDz9k30qS+NQfmO4zGonwAGX0afsCEyY3zBcMcz4EimietjwtgKc8/GfUY
4gR1ziLTR/7gdroeSyPRxUfBF09aLAPCmRq0C8o01t06SC3XQ/HzYG69SjV7l/vK
m+a4jOmhcoK987XxYiBePmoai54q48VGjZptnFvISbObs3/vHkcYqqgs3swdFvlu
k5YVMua11Sswve18Q09lRqZhHsEjyp7P3COxN0F1EcqTgOAdwxCs03TQy0LAKmr7
rhw4PCpcExvXoSOLZUApN7cTRt71ZkuCbd/5b7l/1tCoUB4pswN6Dh4yzN8+mVav
aiz58pzGos1WpX6H/JCENhicKs4b97SNZsAnhCR2apSwbGuhfiuyHyeJ3PIeOlGj
Nypr2ofWP40qYXYN+aAtla9HAwYIoJNsaLDpcFoMcNWLI62g1igE9GhlR4ZtYK36
tfSE/ZpEuFQFXVjzEtKGPfM5WowJNhk02JIvhNMc8wNfGy2d27FpaHiGVN3oTp+5
QQFwtGzoyAkaLY4yiOwwPXPIun2KnNWWBlBzDPtW0hVBa9hxP9PtIeMywKcCFcXD
FoqWAWklVHBUS/57dDU3hfAxPsk98BhiNiddBY7yydtp//Ly2faPUY2bmk7wkuE3
NOAisiyvpYG1t2phSSRQnuP78ld+dgJLhFY9Dr5mwLtUUfyEiyMh0ncz1Imlyyiz
9bySNYualGbVknVTay4HB92n0zggtgNDaOsS7FdSUhCVjkZh5Ce2lsjOcH41ViAK
bnF/YsmJxMPTc0YhmXWQSxnKqHgvAkb8YkIcWr9ba7VBTGy2DTl1q8HcQbRlJ06M
TTu6aqrR1A7DZSEpSL2yp57X+l9lTtVxkf8CyWt98LLXrz8v2N7Lu2Vm+XtsAeWl
XAsUaQY+CVcgEM5rFleyW86aaK3L/r3yoBr/uRbTxGd48KagOGNF8YyfG+R1NBaI
1KUn5MebCzuPC4b5q0ih0DpTvrh1CUCbZ307UN0mO0kmWQgeBT41afV2h0uNs1rX
jpi4GiOaf+ok+WS2MqMrROVOCV82B52OvvUIb2U8OLyJ/GFHoa1tWWam+vDuo7mz
UTmRJcal+49dKp0t9fd44WF3I9Gr4HIpBrd21tiBeKRk6IrtonJIoyvNNA+MIBBK
pIPfzy5RYNLtGJxzMSSaUF2pUsLx2UPXJfJALBhzeUVEGwZ3+yEPEKkodahwwVo7
3/SCRn5PNhk8OZJziGpCNgngEiXLlk8wrIxRFnBtKM8NvHaG9hnF75xGVTFQ/Esj
Ra/Ffaobyzqnqi0A2O0XxE6xXyflVtHM+LJBF0B/klaPvolJaWDVimOI2IbrApuM
4hqrjHRrWxMpvJjoeqGy3RvYrARgHvj8VRCEM/fnZttuf8euhWpLIxn3uAFvZmfp
MvsxkdHxz8jRy/HbdZx062cetiYnuxIPY4EaBkyDdiNZOgrQpVLWNo7mK3+l8EFI
kBB0fjv/vLA+39AgJlJ2GTrmXiaNCai2PQkNOLblRu7y7H278bQpEX558LXCVwnb
JQhDv+ezqwn4D0bAx/9NsmWcp6l1loUL6IunZeVVFxOkpMEsuMYYlrSObz57Ie+Y
CRkxpyaVTciu1KIr2o6BXn/QG2MxpjXVJz/ULir+Hw/C/0/GmK24XEreYZFq9tvn
5ZjuJlb3tnu4tXumT+XZFCI3G9oBd5CCmn8HoFgIrtfUGkMwvmDtTgzPDWyvvMst
GUi90YYSGhnr3YaQxVEMBpthaVTNGyUmUdg1wDnmwNdjHSzIFlXR9ZEInK2KKbit
2F90RwLD2JU673+ezRmjKs+N3dT9i+rBVGUMHeQImnva+D0d84D8HjAu1urkG5tz
Gs3kgc3QUNKJaaoT7st3GrQTandloOQt1DrGqLbb1w92rNnA8GzZevRVQ/PkPJ5/
vc8W4ORd7t/2CU1+VD06ok1OwrjfAVHL3l785zVy18Q8TTVOxU5poK2s5aggvnXi
POMdECT0Z88RsSCovIWfQQgM0Qc10JOFY83muLefFXLiuz5y/sOwjvr7vL+zb4WE
0wurK2L4nl8x/s3WbcZRi7ghH1BgDbXek3j/H4f9xMoLiIET7SQ7ONYw56v5A06v
X/+rLxiZdM0THYL5jiLMWGRmGShaK+SjgAVlDr7NIDPYh8jIahTz+u/i8uB2sECV
L5eIh1vX0iosBN35aWyhsuQGVeFq58nvTyzmyPxI+ArjwgdJBenbKGscV9aYxCFT
wVQk15mRLu5tEC4bcD3yo1Q/6oWByVLnOZjkbhKi7rVZGhqH55jJAJ+3ZtSrrbe1
kr2ox65/alYAcjYD3cIj+yyxU7Uzd4+D3cTVhPrlqDR0uTZ8p1Erkh46155akE1V
K9/SiSk1atlUQ0/PdbINfeJX3L2+KwXxAJpSnDZnIvbZoOvbI2C+fAMLHpKDs5hO
itdToJxUefu29vZ7VCgkMnANTWXGNNTNGxIbybEfyNXqcl225lpsvb1uJLMU2Eq+
SHrRCo4MZrTTtqPzKXmeqfoXtTw7HU+cvB76Qg0u6zAu+CgoOALgdZoMEk+31gnB
vk+s8Lv5/5uWTcHP/FvXkNdtbG38CbvorBWBAPkj02mm0AmPvL0L08kNAXcifnd5
MskLUTP6dTkT9wYF9OyZ1J6PBdvPSSsc+2qVWgfiJNr9MzUp0D4peTaQ44i4Kl/j
JJ7V3m5scqRX0kYbVSudWBQKxJti+/FK8vZm8kX5eEiaZuXtSptAXdai+VcqVkgR
sFTxvrrn0lcjEGwkLgzt9uxE8LFsSnODcp9NzZ1lx3akDAhV/Aj7R+Rw9cgAxfdf
/pTWo7ng76NFdfnQNo6i8awhTq4IymX1wVOSmzx/O23ELpJ0tSiCsEpES9AGkq9Q
wCR0rPsYKWht+/m35dnVJ3frU5Aet7AbTLNggs+7T/3CZUsVV33EIRjOddo+i5R3
JH+nCw2WyXVW8NS6ZZ35dWg7TsbCVWMNjpLRbdlYO+9k5P8E0Ot8I8kO8vO0PcCY
lV1N8fseLYfeHG/cN/x+Oz7NTJjMPEGHzq1MHymprnsPZkW32+k/8UuDD/1xr2mT
PFYWuXaE64r+Y0062V2HXfLoDAGmFs1x7YfTn2+uIT+kxB2jtxub1QdiaBles3r+
QZc0vq2PIhRctWS4lpvz8FOhnEykLQTqBI7TY1pukpug6Fii7UVdF7NS817QOBsE
5iA6MuFdhBJu0E7xCCUtlINAVjU2936X8C1MFy/51tp2eGs5QKN6+Sj3AEBy2+ln
vSaI2IiIHflXaFEDljWg/RtTh2uZux8oiVkpZ8iJG5rrAOT8gorXItuOKkK57seJ
KKwE9X26T+iSgPOSyoa3gumVl4XKbcwV0UXZDNH4hLMc5W78e/ItO+s3KyD6dZL6
Gzvm5fMtX9vLmwi96mzHIIAh+sGQcMfZTGNChRh2rj+Wr7KhZMwoUbZAJOqR90nL
zpwBl37sOszYXmF8zTlN71mL7UH7DXNB/warU4d00XqUkxScgrcRngk0s+puiss6
Y3r2xVUysrUuyAH7Uju6b/BCVnqpnof98uB65hZX8O8112M+a1KFT4RLvobkjxWX
Ri0RkOxRdNmKEtmtJCxCdYccumEHsxejB6DCFbhwZNMnsi0BH7fJzik0DimOG/b7
RAl2ftqHiIGwKXxjDr9tubjacbovPdcFiarKdPVDbbxEoo71I4s/jxHQBQclAMib
XAuK+7jyXaSYu3cBQMV1dJrpWg64jGbrHu5dNxEn4y8AdJt2C15aUFQPugqfcYXH
JNevB2roJE8Jzkp+OAZ9jZuhDkYCdnW7wNL6SU1Nd2Jv2JS+LL/5r6yuUuBcttet
YssoShN5z4XQBgbZmv0kyH08HEGaqsQC8CCaPT4aYaiNfqKRHK84C/fz1+2ATRUa
hwf6JCf3qJ79XCaVVjNVZJPYVz1RIbekit7HBMwQ5YPtIYdIQfwxYBIPRJWt6dYu
KRrr0IpagZr3hdfCSx/G8NXOxvRsELTVRc5nLQ9+GT25cTAHkFkTah8Oulw43P1W
hDweAa7/kxHd/QAWYsCekSwMbhb/o41JWPTAqHf1rQL+jaRcNQlvV8aoFqq3NuKj
qL+kedIWBjpQdKdBvBs2MBYGGK7D4XzC0As9AZAgsnDIjGIeoRAJw6Ra9a7UvhDV
ni+fn9+W/zBJWVegMHm6Zcwdx4eDkNA+OnHs0Bjk0sE8VWu5kkcjhBmk9tb0bGaV
+mwTX7IvI9zpfvuMy6J4iZWjC+J4Zev+MBMt0T8dHh9HQL07azJWfV0P3HpqLegB
qCGgyvWCG5RrV1YQEY42ycPiXBi5rqp4mc9jXr5yt7tpxCqCpyxIMlKQz7VMdjx0
1usOqObPRw+TSGwjPBqE+gvB6uRaKoUaFUQaTHzlXfgWtrytNRHhmfVLDCzG+F8q
tZjKmfYeCuO9MLnRlZPM4tc0W9jJ6EeOfS75g4W0HcUHFBUeA9GnXIxrZpB2ED1+
FlBm0BFGM+v6GLPsByW1hJ2W9OVvV2Xqh+RGBcXzMWHTGi9sHSX5kO7qVbkD2iqC
mAXsxGRuDDwFXx4BfrIl34JPwyImYzyOt4Ao3vEaNmjC6FuOsGPaLx4iK+wS8KjQ
sCvHQCF8Oa2nWoI9RX67cTiK7JzPlIQa68Tz1oypIx81wschDbg/El+E5gnBsmwg
4ZB9LPHtS+K1qC4Km5nRwC9JvFHtrlZHjPujOoen39kpXLOy54UN3mo7JSFRLRHk
XxYHFNJwfPmGy6X8DckaRo7CF7quHMbFlyUIqBaC1IZkOOD9pH0aapy0cRmzlP91
DFgqIxdqzXmY0/CnGsAvuCylG6Nu3mdD6XrjwNBUDHVoYR0qMTzqe99ZdOaSzC0k
TgfibbthiZfIQFWY3HoMM2kfgIeG8z9VgeEo13yvmCfLQ+Ergdn6E/zDS41pc8uI
gB0ky1Xtk3E3jNHPQgde9bKXvEKQQuBXcdUlxcoK6qwb1KugtvTZaUfHA0DZsQir
j66SPZWsrfPmjr81/WmvBIBr7JTlDUC2IvmZ1h1Lk8rU2HKgC6cqX7c6sjqvfY8f
GtKJyXheYrLD49vRnBnoPuU4qa5gZ60Weda/V7sVLcY7mZlvmt7vsnFnyjkdRO1m
UwuoYj/4gJWYWFMqETsF3KDYOHxEhw/n6KVrynPRTFQ2XS0ErVOI1OTV6LcVpSEk
YoFlxC+ycTJVXCiU3jku9Efansckk8g2Y5Yrd10pcAUcM/UFREH6qaBRRO8lXnGM
Y4znU0x64PuLpUwph02/+BM8tPlpHNPKUwUdsTyLLkA5ku4RqFhbF0gy2dGl+FmQ
n6E1xgRxprjnBv55INB2R2MsJ9p1DKmhUAbAxBbfn4PjSI2XTYVz0BH0wLi6PB6w
v3mY98pXM7LWglzVeeJTHfrLQ5RTG42EiCjs0S9OoEPqMhoHXmkNEMibbU3qnUim
VPiXkbk0zsQ3zYdMqDrDv4GAa+78n3+Yr/OcClNeciTnCU9M9TMHy4UK7iQwJSmk
JL/1FgCRLsnLSvknUtKX2N+3ddxIk//cRF6Uq2IHLYQzsu0P5lmQ7qfqm5tgEiwG
khk6GTqS8dQMUWcCW9ZC3WMwOhPCW+dwBNK9DHkDBtLZjGwQrCYl2tP/iAW7+OVz
9LQzumQ6x5TxTliWcbVL2zo2yJhOp6LRDRz/cd6zQE0+0/QaGCzViaK1O/FS1HAt
+7dSAPPkvJa5dpXyHl4iSVy2oZ7rLxkFdrosIcfpktQPOV7349htLGToIetAtjmV
UPzYsVAJ5Id86miRBJE9okkVHzsMEhZIQx09aJxs9xfuM2ZQNw6tlYec+5CninvX
BAK7fUf4R4FZIhX1b4FnkL8k/n7AElRaJYDyeTNoSaNcj3extnPBh/cu+bBi0LIO
MxoATNHG19Ujp4680MYJ8vJhWHzq9vnlhFDHzzn9nAcN3ONi5iRcxo9Kqhv7OUX6
cl/kGjvGjPWcAadd6Hn9k6l+UF7DX2IkYtN05mGrKqrDk6y3J1JFDWC7ayrl2cgS
8f0TR6KGQPz9In/D4GE987p07y84BFTMJoaEsemoJQ3R5gce0+fq0/4ZUAce25JM
NL4XZiYeom9bzEyIcw8WwOp/+bpXOKPfk6i7wEiuVwTWOkqf9Lg0KMgZyfQlOoPZ
zbZEBEuzh339EECOoMQ665/SYd1q/qyxrLc3A0gczZqmLw79E/4o1BAidKbNwdvG
z43ydAmY2VPILz9SuhE5uO/tVoDwfZUx8W9070wQDpxBAl8mFQnlLW4gRYAMDk9K
LccLHAynvgQgwqi9PFTuCFN+WN1CSHPMJRt0zx30yxwxwNrk0TirYpKKOUSwjs8K
eaWSaayyf4xG3ySS9h2knikdPmiAJ6YhTOFQwU7zszW2ubpL6hcUY96SHUZ28E2M
GPoooKQTlo87rXL2HvROPgtMSv+p6v7GM9WwEMySroM9f9KFHM7ydsPHogwv9aCf
bRsvFhfVSDJwS5lesEMP9jgDpoIK0Z9pEJR3/+XQL0xF54MdKwNEsQLEEcxXllFZ
h9Ru4YF3T1Hvnc20ObYtFFO/yHMVM7t+r7L60dYLllb0EGzm7KMFWmPr/6X1y0FK
zey3N91gniQPfDldI1uG7I0nt8j709aH2M8MSE7EHaTiSgBQoX+9iPpFQHPCAlbN
/NqL2TK8Oq+Y7iXO5g/UoFPBxASQG/ptM0GWA8KVKkYM7+sLOVBt7d116xgcOFhF
PCLugsLxPNpWBFtAy3QkIrpNVsz9yPvwQ/eN4bq8B8xqHsKEW48rXGENnsLr3TCf
/AXpqs0Bf+NNeTWWfFU6V8s5WzWM02iePZmfAspRusWzWcMQEt91niT5xvY3sVU6
k1/vNeVVVjuDL7CSpgeiSQ7WBAnk7NwRoYBqL0eC/UdU2ySgQO31CPI4mber8Yoq
C7Y3HzruKnn8kt0BqPmaab4RlCWsLJgQe+b66afBb89a8f07OHnFIJBtFZ27yrGb
4Us5x6McyJZhaISHiVNQluR5bs4ZE4tkj9sjUM7k3hQzLl6txu284LeKUXamShlo
qL+1mq5RQ29WfPtk7Tlkl+ebE+aPQk376oGH0avFCCshDLHtRacWchykO2qUzHBE
ONmzlN04nBgyEVIe5yBkJgqPvh7kfCTGFE95I4QsodGZ8cj47H1lcejhuA+PPOOe
jp5w91b8ifyRwY3MXJRurb/L94gABYym8+9ng4b3X1pIT2F625UvmuWLJRJ+sUQe
pFj25vpiSsW+srGsOCSzhZ/zO3Q0G0qMRAkz5TK5G7Ne/spZH8Tvpj5lwORsE3VG
GU22aAmQeuVjUCm33o9uq8lt7BhDT12/47bRSMSagYAtj8SF8WNsFhrSiL9pcH7t
DU/lmNnog6LPYHw5tUsDv0ys605ACPrxjt7LqG6SMX9U3zircyDJPElCGjbHBdBc
M3+cCjlRzI+NaSIXoY7lugcD68jANU+fTb8Sj9uX+B62R1zhjTcDB1Ujowz9/rIX
bS+IN04tRzZzNT3WTLdlzDMikr6Ex5DsDUSVDsn19TyM4gxxnF5guup/dU57y+UA
v3XFYH5zirUqW7dqHojFbulCxRVEX7k6xiA6Rt4fn7zEVqHEDNS9MhGb1i1M+0dY
HvqmXXToMZCMERYJQLOlumtROiMvwYFOKZL2iVNN6cka0Phpr6bPO+qcIPYCkYG1
Rem1TayeNgIeTseF7pi17rdL9irugGqhuRLNIQc6LHekV4/5UkSN1Fl0hlqRZR07
ICXMAMw179q87VAqZdZzyioNk7HiiaI4r/pewngpMVRxTkrCjw2BBD8KKqoHMyI4
7IFWTwqYHgMk0dX8QlmWo3l3waFxXx95zkOZ/Z7y01pI+TrFlIa1PAZDsGe/0Xh3
oGUy5lxisXiPNDKbe4C163ceBUgucwTq2dca18+g30uXO9J7Uv3z4RJQ+Torg/FY
GRGumshOaJMM1ldLVYXX9aGh4gHe4SrJPkSdLiShRL1P+Vo1EZgNy0iBOVY2TIQU
GLWtDBvgxCnTvegrua1CFj4t6zadgZ0dz9+QSLY9+AzqvQ+3zTWs2S5rc+E3zpPt
PaFlOhOu+kQgPMCl9Pv114VO6m65XrmR8bk2cOyl/npJ2fsg5A3oq+aC+ZKNgatx
INhzKI5bI2SZrDiKTz1YeH/li98ZXhTJO4pr4KXSIFRrInfFPov5zCFKd2xAm1MX
csw24TExSm48CXGka7dSowpLwLXe76cJxlO5PtjzWyMK8IJap1yKVh1PCE4378Mk
UJ4EK7PsORRtydfffV8+vcHaS2kxBO4DCdXQkTJhet9Qw4+AAGwOeuSxntMNRdQ+
DKLHR/zn/Jc8jVlzYYkKRus+V1B21zqy8Dg/4jtmn0UWe3FkyHEh/PP7/YM/SbNz
zOJx2uK5PfIGBjgQRurla58KWJ6AjC+7rtuTWterkBk13Z4Op5K16uJOMkMqXGe1
rc0OdAxYSRSOBD//pdBMgTdbD5ehZi+TfpfEnmsmkielXNVTAKYmd+HgN+0jT4MM
mABKI+rQHkcZPOcoRspoEj31dr3bmEqWzmR7Ypz4L+/ADd2iFwZJkenKzOrhavGA
+xX42JtVmaU5IXNr78MIIZ8cBkB5szLM8RBz9RuI/ouW+JJSGh6CKzNGsiezM51f
doWg0oC1nKdEYU8AFUpR43ZFZdHGQUZU/bSEUfCiCmNtaoWDSQEHKtFxc11K248O
BffiG14eBvOd3vdSnTlLE6tli5IU+08PsfeH0YvusmUhbTEOibIJidG92HKQ3Elh
cTdHeUdWj5xmFSkWfa4ZlRT+Uhi7WYw2scKvUaNHqWVCDaLI2aLrCZDjqKNY03Gs
1yXy0Qp3WwXeIVuCE5ynvZfywV2zGM+RC/crm9YTNRRqDkqsczxTU6GJXRHqq2A0
AG4Ic/vXs+l6+A+paJ4f7rq8oDUxe6qgYnhEMMGTCZSV92LAWru3AYJmvmN76KzS
I1rg2x7pUeKaTsBOOvA1zUH9r1y9KPT+5YARTDBdn/x3jWe+ddVlZNc5rbxgmONP
0ZAk+ASeCE5pReKWl1U4L7RMS4eP8wYsYMyITYjxmN4Fdo9NQAN4RcYqRiI3QZ3G
sEsyyB3DGs/1B/F5DlR2ZGlTxReswLtjryph373hZb1KBOPA+fyQbyyA/PEFIPFY
vkOKdQe1RkB8hkW6Pne9tJElwp5LD4g4CDg/TorZWnUW4LcwAY6AflwgscFyQgbz
nNZn9Bfi8peHn8MzkwVFipqz2KEvkKroCcA0qdA/50P/1hqwrifO8kQvnfE6pY9X
jIYjY6PGDin5NqHmYuYblE79AY0mFWE5jDCXq4FhcONDy7sT5bJvAzEWoe5vwI/Z
PeYYKT2A19IEPJS+VonSxSQYOp1da0PB8eXFamuEqxpDoTTEUnCNGrcOqnvkskwI
InmwsATChtnvlIy0KcjRdbVXI4xo9C2/iVljq0Xz+CC5/9juNdi3yV9yLjfoxiL0
Dfda8nOEtFWL1F+dO5+buVXsp9qo9xJq8qX5JIfaprONc3MqQ0p2TAkGIekCoaal
sOTq7V03vFs+k2zM+Oe08aJNneZplWzCfTRNVA+wiaK/WL+sdcdaXVx8gEdAVTmX
oY9JiRV55xMgGhEWnxZqFuuShEdKYPo+0ImVQbKou/aQV21AmwAiJRzI2RiRHvX5
RP0EmrtvKMXNhiiR4gtBY/eAniYyiu1kC0JRpt4PlC2RNEqiNWzT2fhTpm4mNtOq
nTlNnLFFZiJa831XLoKYoQcfcGyFSVE0C7JpSLyIsOaxYlIn3CHCpftqv7QRkUMx
xrxvaABIVj6zC5ST0anSJtO8EO9/HUHcHQ/vGEf39z6nE1XWWuC+bbHX/DJ/85ZC
aucX6n7qeZL5uEHDhKSCoh0Mpm0kt/WrPmtwK3pguW8YzSrCiacv9Frycq1LhDd/
D7d5miCA98pOh8f9PThxzIgvnpYznXl0n7FTn6PJkeKL4O3m6bxJsveazMaFWYpR
GyYkKB1Qy2qxfPaZGpRxRGsbktDzMwVgOoRhahdKUMXS2nCe3xrCXP7WHiuYXlkP
/HW1pvDIDc63gSTLPM583tcyjp9SdVvgpuGWTOQm8hE9zmR1U/ebVTgPxicKuG5c
CNHlCAfYDeNmrLerF5gAImW0SY/FwAgr74GwpeJj2hBHstR38ITdGRG1SeSE2ZkN
wwGVWcx+EQm7fUAIXDCfRdysCDtRixS0qQCsyjXD53qFAADVzl74PtKyUxf7JH8d
CD4Elzupf0X0y7DYp/ZrCJimq6IrUeRj0fRXg2/WV+HJf+7ZrTq84gyB+tJJh3aQ
mANO3BcGFtSdR8lgoOHz8DLtofndmRbXqQV13bsGKtRpdaL4wAotR8+2y03YVSHF
WqKXh7ZD+czq+E4q9L/EidouwnVehsTG0CqEBOGB5Kp5tKvIiy6hc86gbmITg19a
TbCb+KEhwk/fOcgHkZ7SD8DJ55M3BETDo5vM62fJiaYBncuIfrl899ARTIuyEArp
XddaZnB48/I/Sr+cp+vBg0uPXDyGWV+REhqkpioapZBC3gn/S9qNEc5TPQ39LvIi
pRvBhHBwCvb4d2mwkYAtcRTUPO6hwDZtrtTqKc1gHi4+VF5Il1s5rnAw81yE59qU
SbVxp1zzVnkPfKrw/83ykJICYWbaUGepvXHoIip5A7z5o61k2JuTSgorNAvNu3eb
aTXhearT3wRRJh2vc40Pg0voVdM+Z7U2i4GVUR6Zn2pJleqwwZO6OZ7liMN4NDbJ
IFnHNP/obmUoslXXEL0G4SZHCRSXsgPHvexb+Rqzm9zR9IzI6naMKqT0nMExOhMB
SZ1gxoO4YUdDXocQ1ofnEhDB+Ls+5C56jRfnEFufYdnTa7LWDnyYmeOFfNH4FlRO
bPuJl6rGmgRj3hMA8phODFK/UQr2LbhHQ1/dEDZwVTAx9KBiyvOS8PnRYaWclBnt
0JPTUTeDUmXLRoLsjIn/tUe0RF3T/eEQC0Am7BAo3WXOhOkskZtBRXrRkWgVRC1i
V77jcKJgm7m6Vexcg/5D/v0omNCHyN95+g7kzhSV4+lK/BOnsUm7q5AysdmMua8h
EoYTnwSojcCtPr4nk3wX4jrNhFccgodGTx0BrFdra9KBGTGfr8iLIWMbjon+kdp6
9LXzEYn01pE3CUGcBL8D8AzYOknHzANpWYPEbSAR7hREdw1zefhZOpL+sV6vxMaC
SfD46eE/Vv38GXqgQHdbQ2c59V5OTUL0RjtkgXPhP+ne6AIdSU9hDz4qQi5ESAcE
Yhuf/D5UwK2VhZNMa2K2LFyPOo/cxEV8kcwZQhf+AaA6Vule0Wpnn7JgSFHGGHmk
PzAeP9oKzDKIMoqndiCL/uEVoebffw66mE3TwlANUivvpeuK/+AgZl9+2btFMl2B
o3/wkpissVOKP51FTvfyOrNADZJI13F41hzjV3cJRbbJFD1Kei7hJP4RTHYHd+tr
4KSsvZp/H4pKNGHqPYk83EQTmWPL5IJSujUQT8bQMql1wX9eh2X9BaPKvIZzz9sf
AZuaO6beDgxmpk2RzG4MJ9l25D2LdMB5+lJ0G5qjZYEzwTeE16EV5qmzpKUxRdwt
qgWURfCbu3jk17Kk69oDhK7BfRUrZYTkSy5nxQeLYzAUPu3KSnPYTFJSMY/conK4
PFGczNsJQSemCLr/FsOTNS26qA6diy3Ko8ybNJt1TXcX0jxzLH4cr6N/6gMLYZ1G
lGwJ7iGFajeqwl9CD5/ycq/pCIx27umVlCJRo4KIkqZAWSiKYnOJBV1NU5F/VcCg
UgsREqRHMajCLCqnigxtEa0Is/ELYdKAIlaINnhLQfFG61Wd2ezIwqZtc4KUng5l
oJCTVanf0AJYQZpGuqA27LJvCoaFZMBR5X8SXwDpmFPJx8OXo42BvZSf0N00zq0B
KGr1UgZdRW1OCipNVI5CBKLb+9u+bXcB9WOoP5RzmC9hkp2YjKmVeMqIXoqZ5YIE
i6hqG1TkUQJ9n9fOTxENOksEapLx3ha1pEfaWrWLkAbtMZhjFBBreu56PyW0wUnb
tRYu17qPVnfXkV/mf2tLgC+3r1Xu9PuNLUjrbGV+7X5BZsojMB+LlmBjNbiESV8T
E6SyaUSkFKYtgkQ0KojyfVc5w0LrXiz/Gcorex0ofoa32CDRdBYjuA10JkJuAKoq
HXlk/baEURP2WgV6BICrsWIEBvEfiPUOyf5s3YsoVQkWMamTV5pYX1dkRbUIJ6mh
hZ3LgVhkyL/5dUCjD8DgfY0kL4G682Re6Eyaw+JU03nipeYM5qn1LRS9E6Zj+rPd
u5Q8avFzn5UkwIbC0b/l20bTpBNSf9nrliP6QcY+hDgtCIWn2PARySGvpFhdACZU
YPswVQIpiyb1FL3g2tqwOeVlbBxyIoOG/ijN40IV33pjgk1pm7vcI924A2z3SWYw
nUiH12Eggzdjk+hejSt+8Lw48bO/aLylNkBP+4znJfnMHQVZDsIe4eXvKSRARoEd
NKYlGGZa9IeZkohw+J9JbWKIU96QpQZyYC6PQo4eWXyV05GKqLV4vKx4qpd52FmF
L03vS1jHhSvch7SYv3fgH1bUcDxQ71a/FX1L8fpte6O6qodOLaQcbsA+Z7N9MGFQ
gCi+jvcX53ZqPs49fjP6cSK0c+QxRMJqPE0GQWUwanvmIUR1BjAAvJqTYRJJgxOB
HTE2qZHJ+imIlSvC1fqqa3+eeAknCBNYaGbpjK1oNgHeJ88LCJD1M7blmko2Z3vz
8+zEY0wqIBDsgX6OmNlYSP5JiiYK065gujEZHxQbuBAtpvpOegitqPCfY70Fzn/8
fwkUH/NWhvrqDA1f8BEmQjSkBsoDb8jpikawrBEnYMJM8HU5l0vMnGHTvQrgQyBS
Gtgi8cOENkOeNQY8tdSaUcqqHopxzkZCT/PZQUg+IhcSltCdOfkl7OsyTJqbr0nF
csY+MV/1a81wKAjVUtj4wTUup7glBk2mU22cKf3sJj9r/ZFVuo22/dMjxnXyCUKR
xDTNbS+vxLOmX4hPVWa2gVC3zkOr6yTbI3V1WJzRzTnEMFeMW+Hm/xPpUMBkeVRi
vJV8K8ccer/vJVR9eYV/8Qt+rRGg3N+VLCaH0kdRAAPytDXXML7Dwm9cBJ966/4M
IHpKAf1w0EHvQcfApfCTwNzfRVMRG6cP+/AsTN5g5qqP7O3Lkf7x+SpwEqG6ROEA
kA1GSpxNTgz8hy0QVnFJetaw4ccQni5WjzwiC3bFrkwX2qglp4ReS5SIMpyS8jO2
jDlcKYIVGAjjjgMyZ7sQ6eORj2nV6vO6N+AoxDMPwM4qGTsfHSTLgwResTPvCsmR
Xm/iXO1oRXZmJBKTvuTuU6FX7M0X6RQ4IB3RGZ366LlTgqv/iOtH1fGk9/N3W8Fw
DONbIFmcDjBMcvwn/oDkGGQemAfas0XfW8kk9OIasK4zYjPEGxKUZ0PO5BGgVuwX
rOeT4ptkGe9k5pWlrjTn4cjmtPyug8LV6eKmpwd3wEGtmzZKE661DZ+CCmDENJaq
h7uF6duLswKS4dNVeaV16u5GWGIItD8E4QVzPoGaH/7fDmDPI2ViHdPgjdqzAP4z
ZKqQED1RimRy6G2MX8IlPZU3FiAIqgnSwcJHO/UrkWuUhBFMCziQlehtOvF+9frN
uuEOfgItCxfVVYmiiklh7pIXOaUH4O3bVlD/AyNG9ddH09LuFeQojNRfUszMfODK
bj+pFCr10/r0ZbsOU3zk8NkhjoJ2xyxNAdSsBxuGzqcfix5qscsgeuoCQY/r/YBo
BgLZlfkAXx0+IyNP8UoUpXxIqGly1kQ/GIDpQ7RXBmahtEM+c94Q3ksWk7WSIS0i
5Mc3zn6Q+848D4gHuR3CyJUIF1HnJCjBInrbskds/X+tzftxx5jo5czQtvPhRSt8
9/742v87QDHOUzDyG3fJ6rcWbm1ckF+HQ6Tp7L1wy7UbeuQUP3GJXcYjUoSh6dy0
mp4TYe0kPoraUD2aUkRPCslTbJ9H+7m/c67iuCWpPRZMaF/dT+QdunroDopkqZ/z
9CFislKagG0KyhI14ap+oXTSjf/3YNtLlVGmG7vKiScJWThNOpL2FQQRZr2MaX8B
e/0IMQInEG+mqn9YQDqm3a1m3hl4Oj0GrpHYbsgePFB74RR4oZyh8TrZBPF8Wn7B
pFPfBr95ua0Z4v1gk0oNiTJ9+jcQM1HRDUODYVhoX5s0Iv4tY4LXTssMz3LEG2S6
o7gFg9W6k/ABNbCzGojQxGK3J3wxH91YSwoCwK2yxaaJDU2Ewh+Pn+K2tU8c/f4Q
0NXUa+SoEnQI7BIer92ZHC5QP/HNj8Bt7V9t+0ayomTfDDYz1E1m0TPbXZ3wYiZl
kfYhxD15niQzkOS4JP9Kt+DC6uIh8ZRR7/WQBin52gkhY7FOS0X61bFnNq7j5758
q49aKbMx1lcVijGCNI+jNuJyLWkIdAafV6KWNH98oY9RyM6uOt7CU7IBoF1qW6cq
hcUIyYb0yMfRw9WCbrEwiYbbfkJTnSOsR+1wG0gjtPKmhRXJVEbP0RYFW0zNaGW/
tNXg1fXxM/Q+AUJdITJRAFQFHWFRPa2VrTXv1FTLpO9EI9Ub4Z7Pc32Vk5TalmVb
wnqugr/HBYRftOgCm5l3JjVyFeMkWn1z7qrM2Q3eYSoP6TRlvA2i5TBALgQ2+UQr
Tqe26FUoxAZrFDSTf2Gzl4At/LxhXN0DG6bfTh7pwc4mKYN6EHrIlglOzwb40wkP
bD2YGxn2BIwiMWUn96lOXtYWRUPGj/nTXh7FEKVMFP6v65lwk6+r/t1MY03yI5GV
anNXW4uHwOZHEn7HhNX5BHMdAqOgXZ0n5gIk/P6AN23QgsW5P/e/8QdKd+ZIxCJD
mBQ/N+1+WUM5a2KDHHMnAYiAnrHhNwkt8xCQAb9aKd1TTdxphN30Z+ob4ZfzJi+h
dy9CNA7ZN7hGh/9yfO7ZQVJanqdWrNUW5l0sfnjJb+2J4vSwIpcGr6HyFeKh4coS
KvBdbXDqu3VzpvolkzZ5xsh63vx1UzizoFaURJlglBmRDJyjtbHw8vuZqD1TXBC5
KT3k/gSe1J+R10bSjTgtAtMHQV8oWLAqRstjoS/PE4s/bKensOtf2SaBVeidflXl
kYDmnApcdmQy/Xr+484apqPBSZCg1ygwRf8aukoIWAiXU/LMmDivtPMkB0taaB4z
75rx+UCyRr99ohGR+E6zJO9T06zvca0Ou/v6pwmPK6CCWQh0vgxhcPs3ew4E6ewa
80ToKqi9CyQ2WVxAJq9XjfTKv4uYHAemCS8+NzXiyXxnyLrdPqkvPVMd9w6uQTg8
NGslQsAafM3wziIRq3AzpmiHV14fSIxFUyUMgLmxKWV9HFjOmvqmuO9ZP29Kx9Ip
p4Vts3JKJ45eoRaPa0gykj0tt3+0BJkw2bOqoJQfUtHt9/9zts9qJoOOavU/Ui4W
WCkPtPmZhZmaQVuZBEoUzsjUg7PW+WNDIDazU22xNZzMWZGqDBJA0DU/vHFebayR
05UIN10akyU7DageonhwoERnBI6aGwRAWHcZ39fv4bdUB+hq/6LQWQUL8fn/xfB9
dFMeHIFgsf2SesTszuR/AL0EbSzLEnECdocd9BEnw22LHWlfbqQCWutlSZD8NfI5
AiZxj7z5pW1UesATHKE56QwCGX4PMsdzRqZrQuUrPBD04gBcZpWoJQv/Aum63sFq
RAL5DhN5TJzQx18ZPiJs5x5jOF/HALhoKg5k1bwPbC+cMvUMrSNc1lifI60PvXi9
2SknURcWh35Fhki6VBERoI5MGQFrndWionHVCxzUmlGg2P9a2iGbiqgUUsJt8mYa
1xkXyFyDqsgQT0emjUEmFYtqp+6Xr8QtQ8g+b0/kAKgHqsf2K57dGqusFu355nIz
9CohzfZwg3qKqRc1LJDw2FB3PEbVYfYpTSLZGkyOmeZGTj2Ru8mVndPcpBq+Of2a
kRF1ECSEoKypCR4unm2qUABIfGykDvgmGXnMgubHb30HgdT8tlppnHR+wDx32qYg
N9HxC5KOeoN9nd/SzSU0lAeN5OtROvkaT9Ha/gsVTgkCvLT6OSelVyTHAoW/eq4Q
BLeaB6xWuz/18HmE6DjtZLGNHhXgalUxCCG+Ex6aN254/cL/3KHGhRV4d23p/ue3
b+k4fshMXHMeFE00nXxyC/1kqc4Iu+IEJV+VE8vIc8VabMKo+JEZHjHeH1Ml69Tm
qouHkI491Xo+nvctRHrWPhSYMFRohFBeANJTmB9VEAizMqakboTLXDjjjzD57BjZ
gpOLVexdsNCG8w/P3BAHq+L2SVyD+JZV+hnzeEaZH/y5eGAiOgAXmUJ33tXkwZX/
Fo8mW/GPMUT9Tz5/Ystj4Ylzgfe9naI8030CoN7025y1bfRkvbTj/5q8AkMQkp9O
IpmHPmcvWZ0bHUuub0wCoXmd5AZZjVorBouqVPAw1oIBsBmop4xl9oOekLfS9EDQ
EQwREqRosQyXgvUjurNxzfIePotLFbm+fnlkNX1du7orReBgai/Uny9RzRSbAL2p
nh9G8vfMYwp7UxSH9+PuOqMD7UtuFrRS1+hftJhLCbdfr01jKA/BKOX5e9ieXKxs
QX9ZODtbbvuizAGOE19v1gZqJAk6s1Gzl68Hc56nX9nkcrMW29Jows9vh8CTmykE
SK+IH3F1TYiKwuaKiyrNVjkIUvOlHrfy10Cyf9sNAK6EcplBP6ZNZw4yxlLKzhGZ
lHtP9TeTY5UJP7plc/XyC9HlRJ5R1o4Saq8L32ksQVm92V04BzEnV0gaJUF+r12i
UdMUkupzLuYFbxv3l8MdEPYtNh80ArLbGoRJnz6UeSUWUdfbyRfZmVH/zXdW/1FD
MQQ5JC8dL667x1mUnNyG0ZjOHdupb+xPK9s5OrzVVuAmxWEk3eZL2aCQZJBEFlwn
4AlhrxDEDLL3PmzlP4nsf/Zm48m1EySSlNJop3UiHXnXBmMr6XFxzXJ95pHRPX9j
fzn55oxSSBvttUDponWg0bQOeCJXpwopU6lG24oYInW4pkpGbosz7hYinsNkCOEa
EQx6BGuNwabS7xytzZQhQGuGJUjE0M/r2jRDxiqslpa+kaeNGLlE9neYUqEI4sdr
G5CsSjZifdehisfdb66vdaSNnpItcPZ0diCNu2QKItH6bjtT+eueE4cCuW1RFnWf
cUy8MfgxVupJXLYtVny9dRVlIE0w87waATT6qUVCUHvELu2OGc55h9H8oAPxYdVY
3H3G23oaCm7XczNArUnEGKDPRGn+YSb57NlUwTVTjgfr8xl3ZnjJ1vGRMEQhLR3g
Ky+4Olo0/AJejecAlQAAG8fxWh8DDqDLjVA+XG8hXFaamVL8wTIZSpOuNdYyaXWk
STjjJ7yLKRdjPlZtNII9zcBJDDnxDelVzKP7WFnmCsaPXQj8uzmdcetDErYzCNqC
4QznaAGbGVob0sW7L4eGlcnDTSSJmveeQb3BlRR14TeIrCbxqaN0Ejo6kxRBRoaI
Gq+inXN20SIz/bQWjXm3tzZ5xKTk1l+UJHka1omEyaXSNp4XidvPCZfWRiQRubPm
6hQMxW6A4Ljcy/ukBQdpn+Cj550HU6I0vMAVufJ88aLaKXn9YhAt56cw+xskUPRV
xWqe5N7Sb04Wz2zxKxv2Z2mqNcdiNtYfyia5Z5/5UR5fWo3re4MA/lrBPj7E5Z4Y
xsQeMVYJMELzIXR+Vi3wInjsiNe3soc4qncOWV8AmgllzOux6ccPBPqRt7J5TDyL
EB8duz6Oe0TCj96uu8zBLFVYc2MVib/qiCSV0+SIlFDyg+QCVs5tITdARbAQ2T1r
ivZnXTpiX1f3ZSq5c4xXFfFYXUuvUgqF4A8N4TzWa+YjgtkWLBAzMTzd39FoL+SD
AJFxBjVxNVA38UQFo4EqLqWTiqNIdYvIxvwl3u8tqlsoujjoZFn1o/NOkbpONQeN
bq54woeTN0R8tjoXZ0CHt/4UU7klWJ6TtkNkyeEPcWX0z94BkmsqsSDXIM+9bk+b
6hpaoTfhg4N312ZSPHnt8RVfl1NYyH2zol1E5H3fAMN2ICNBZUK32d0r8JzeuLnv
J+xHQVgSFYOXcn1R+WpqhMGwE1+49dmBFBQAzAqhI7NeRbDqFz3cl3SXPFJ/Y3o0
tXOX4uzBKkG3zeb0dWxCZxex0cCeqKhKpBs+AsdQa8Y1ggPFolcj/8MbnCCc5ir0
5gTXb+sEWX/Rjr78pwVN9et//qpsV5QBuV3prmHAx2DsbEYdmGQzXrAsbaI0cySW
WV+9vl7QJCCaLixz2yQq5AOJkN44DDW6d8LvjB1ci1lO3fwSaL9D693v+iaPSdHs
L95bg72nDhgN9eLptwiLyd7VC8ZF8UrXTMek3eN2Nwl8zBLVuGw/laVxlEhnER2S
x69rhX+zLaz05KbkJWaMMS5k449+2F654iVqpbQMkfWaCmnTMF/Pp1RBxJbF5anV
KaIUWB5/tVoMW38pC8V0ryCJLFGBfhHdwFa5OqIqPYp08IudXlS0h0nz8CdY2+Rf
yTgerkWkt+nEgQSl2QKOKvL0wk+hV3njrTPsKGWB21S9bxCgcASHZpME09eeUbUq
2Ltvyti81BLOYKqa53k0SYPdWDIEVlgpvweLC1Kbu7VnI4k1x7OZim88OnfZnjdY
AZnRBnR6ODHJoRFHZ1kFbqicsk4ToLIFRv1TxmRaCSJ1jZYI7vVAtfVL7upPZXyk
z9tvJwdjjmTGJ6TCyLXHnzdmgw9fE4gwgDOZx1sQE9JyOcpdSOUqCq/262phnvC0
KOYToTYPlMHKQ+xtf32Ick9dDm7I0hqEzOnJmTw1J6ihwKsp4ZiX+Trn0WuVZfJy
a/1C+CTew8gBmB6joyv8urhU/Xkmr0NqigdhWJjdr0NTpv39LGDQa/+a2mTGfNvd
12jgoj1WllYzPFGx6HO9bYKyAA7x12jIWX72F8D69lEERPXyOFopyliiQySMjFdr
BKwL0whrEbGZPDzND9VcEAG/AbhflJjrbTriTMSBIZrYa763U2wezaOQm521HPyZ
ffW7FmxqI2SkS+iuSvhcTFwxJLgVJhNPUgt7TLfQsNqph8LSrtT7iMI10iJoIut6
e41lDm+l9KvnquDk0jQV+J/C50hqEPjEE3aogjVtUQu9tB0o8F6BHNT3ydHFNMXH
0QBqxtC3dkDgr9i6tnRGTSVsPY+jGuHEvZ79S6Wg735BbE7MExsr7kpmLA/h+ozQ
+blai0uZ68q06K+nKyFaPJ262zdAQylh9ZE562cPBNzKQYtgNVycfVbVKqNKRRSg
mXew9yEGrAJ3ANACg+scBaDPXnFn3sQug1X2NTwLmIXgB14VHkpe76Vox9NOavfB
q3Ml1F5TicWXsTPJrp5MbeAV6PU6Lr8tnrgSy0a/3FGXwEfFRbbphDDoUyX2ynmy
7TEJSsIn5e6MZRQe7MZ/q8Ak9R8NwgEez3C+lqyltf3vR9RMtHfaucZ41C6ZP/4L
6TdLkvHNDgc1Yd0SgOn2bkVjQWnsWzHB10mcmCHiGMquDLBPMh9kLLRroqaO/m5v
3FJ6bWlsMar+5t1SC4Nj4f/prlpAuR4WZqeKmYjb5i+p14BXU+OngieFqmgGsfN0
8DsWwFyA+0g8yTmZkk3TLcvKFlBusITutEU56HbxeV5kYnd6N3CphgpEPSgM/Tf0
RwAnCIIfZZSDKNaRdpi8zRwmeuU4amgMNHEqsgvix0CMZHY610MqBpPLBjoodeiR
/uBjsHyjDr4YvDpsqMMdzuY3hUCh57qgnYSaWaPwxwWjm67X/H+6aheKo37SbcAj
3+1NecSuR9n1DgtXxyzSyMcKF6OjZTP+e4eiVpX/ZtB5VxusewfkcPiHnGY4B6XG
7431yNyRNLGfpUHnhKRvyiFYzDHFa7jkOD8fcsSF45ST3ChRTQ3MSdD0igjMl7GA
QvQiEBOOqI8xNihTG1kEAWIOM5dQ62cMBcUbFAHFzR89TBjdTde3Ioeqs74mHgbQ
L3agf1n9CGi/V01qGU02M/rHwxUwYpUtCXG00n4tOljl50CP8uV3hZN9xuC/eAlQ
tLNuNHGwiOyTqgEfoSmNUDlD4WYMAvCc70+mPCMffRObsneFR9ZiNtD2g7EyAJkJ
HxRkfHxw1tqbu1+F4oYBOYseJMClIHDssI+zox1Ofw6eV101ybMjZjIGe6Als133
iJcruhuWPTatGVSn+OqR/z1fcY4rn0p6URs3P11hStGd+Z6fOBrsdI3jEnbr7Oil
0KTyeQxmbMH4/Bqr8m8uh7QF/PTOyHvVMe8NKkT7riZwHpdRifubciT6DQw06dKw
JcqIzlmaYwg1euoLe+VNatqa2JvME5tsNeI5cxyzAamnT+6pR02j6VIDih3/IcCg
7NGKRdiZaZmfg/wOAHXtXs7I0LwYYtAG0Z7a4JLgNXIJKO6R7lMnoPV8IybrYqLx
UtTHeOPvGqKIr1Ep82rDeyggE9OEO55PPyQU+4Jstd0vFH3vR4Jb9tv/iokdbkz0
iYg4mWC5FnHeXIpVZRNB7CGd7D+5lUkpxrrC6SiWSJwAewodGICufPUPeRNwdIed
NlSNzAJp7DSiLnCX4T5NJ/JarVRKIV6P3PuU1EQSz0gWKVSEbm/8opSNToN+E/k6
ekIg25+z7FCLF45+eQ8oKkkY/LCk4ixR/ltsVlMA17+0oA/BmewN6eNM/oWOaysU
ETQJtFrMC9nT1mu1cKHKg8rfjeg4d0hLWLUlEEqYSayu9GObC1qi9NwNqqSPoBXg
4xS3D23pmouY2J75MHDYX0P9Fudxu6/PnS5nfcFvu7x9x87dSRx5uAIk0AAFC7ME
qNxNzxU1JpGrvgpHqnSfpRk4cklhEsLarClFkXWoHmigVdqWIFsQtU2MrYlLf/vY
OWZCQsOAHhHpZupxNU8KE8PXdF1169OEHuhp6dyiAzKMGoG4h5WLC3Zb87JH8k1Q
nz5ZAtNOnOUTj+c3qQWN/QhbO7VD99Ce7E56U8byuy5bVCPJQ3CR83BqYmz4l1DQ
bx9H5lzubYLSeGE+vwKhpB+x2ZB9Kdumr/DeFYnu0ofWy2JYB+DcWH2WC+1S0WJu
Yqx8W9OBmOxydQ+j9rO1b5vwU8YNuPWKlQ4JRijDp8Tyg2v9Z/wjq1esM2JOtyYS
kTNddF0A8APKxVlxtqwxii7boQAdGDocXzT/H7jKERY5T2nmLP9B2Jo6hgsQodvA
WzK6iFY5pYa8rBQxmM0piztm22QMGbokMsL5Nj/lZH0OLKeCJ0NBW34FJzsZ3Q6q
vZYiVW8V15XLL+6zFGTrRGU6V6efJTzNOlBcNTNGIMQSpkNCpQfJ+SSRgOQdey2/
1ROS0W56iilal6h7J5g85zHNnzZggQGyJLyjF6lBDttCzKMbz0YvU9N2vlEkDuWQ
Pp1S6bad03oM010fC1Dk03UQoYb8mxYoiOSdK9YDaE3NoSsswoYdvbvkFtd6mvhF
GwNiX8YcC2RxovzGoX/pr0jGAii7LSxFcfLV00DI7vf9qQGF3bkOUT/uIRK4IYkC
DtsMA8PIPjjlPWwpyaLt5b1AT91eF4RJJiCLOF/fHXgxs4pQ/rT16tfdDhhCcI3m
H0EFs7Qc0INoyibjy17ozdcN9rRzz2vw1QVmxg1q4knwFT6EcSIfiJ6d7e8gsxNp
AJuAGGESyo7yUgjw3kygShq6ezg8RdT8uMSqDKqQldmUbGqID3Q2zsPisdRcoYqw
bcnesG4KFcfk6jIIRbGsvYVWFQ4WeZ6uJ+nTwmcDcWMK2SPsck4TMa0RP6HUsg4F
SevQe6oZcHNW5GEr34Mk4/hU0CSi6Mw7bKf0mVbiu8LkJUo8xcYlR1xzZKCniV3W
1UDzkzbTmDEucuwslzkUk9UxetylPgMe466hyw0iDGhuXhjGYMClSTKkS5pNuzsF
zqQCbRwUqNOWh+g01qSDezJ/Bk/pDDJzod+Q8GvcM7J6wMrefRYlK67MDRHU9Iyu
faLLn3afoLG65oNnbMD/r/n8Ypkz5yjO1VJd6jkI7+asnrx5TKaPwsCQda3lgp/j
fTjxEVCwrH1xYcKtl5OsfbJSuyllS7uET2lX3Y2JfG5hQ23/UD0hLc095+ObvDUE
a4ylsWSPdvch2yZr8eEUCfpjJ1t1RTI/h91KjOqTECskAp6K16Q6QJH06weUbvfa
r9KyC8FgTAskGBWef5JBYKiMHbzw3ama+Drk03/NTgunLFLjjdgzqfosTH5bq03U
ITc0Dom0TylMl5aRNH558eXH64/h1ihYZSOHeiOUx31rGC/cLq96jciYt4t+0PDK
NUfrXAPBpJTB4T7BrPB3TXUxFyr71Z5XoHy7cqrTAUufOr9YiDuCPW08nNXA0oZ9
fmKJenknuGo5zWEK5znm63b2VIuvrQZmZUFSl00KXqCUX/JAOCh834IA0fvSAMX7
eUKKo6Wf6voJFgTvysB+YNom8kPFZ5wlHzp571TpQbMVl7FgO6Ext1aeAJFwMhKt
UXZ2m44OF06qDlUCWBzcrhVhCT4EjjTdlelukqKr2NDUIuZLRE+1le57C0dmh5sI
YxCkxsaGubMiZKTyxuXjeLSKYav8XtgMlY59zUbN71xGGiW2Yywz8UiipQS3g1Ps
3Kck/nn7c96iytFA7aBlhZ4bWz04Llz7D64oOCnYx+oV0OUxufhT5l0H4NoBfMdO
waLcggyRUyV1SqbPsqTnoK2I6iQJ6/0qBGKEUuDyeEiKx348ykq1dd15Iuxt4YpT
69b0JR8IIHJdLRtHll9Y3c9Rjea0JJhnqn9PQqpLpJRmbyHHcEVUf5Pb862Ps9LV
oMdx5j1o7tjmCpqrYwV0heFFCP1VeISRPvSy3Twn2asOLh8TDKmz4f1446tQGaXv
du03HF1AbbdW2DuVYxpHCwaFwe2llHmGWuTgk23sbSQHIC1AkedmJ/iWM7ftk9Bz
/k7RoY/zBHvLHvIkPazbYAB7080YIDrcMvDGk8/Hu0YDuOZoetn6uoQcMOa2hm9M
mMK8xDIxvrJr2HylSzn46W0e/WDde/aIGoM5notbx/p/4Eir35a42WcbT5Uo82Fh
65QZX7DXCQycUDKyTVi+d8OIgt/liXGsaoPK3OofFl2l5J9LAcP1jMIpWQtlqclY
SsrJVWrlnVuIHl695M97/D30NVSGhR6cg49iErLPfbVGfMGrz069/7Nu5iL9r0/Q
VgOFvLY7qQZcVqJR6jaOuIPcVqKPyJLzSngaAYxrcivv2ONHwPy8pGy4NG3uCcZC
XI6o10TDjK1ce3Z3b69YZDyp0V0Ku5tMckCqa3+ZW0d5OqHsgRThTCH8rFdJfr3a
KZ7VgJ0Hel6CBy3KvZBhY1ieJ8WgU4F3wRzbAk3Qazb9engsml4SGBV1IRCtVy0M
FGa1XJYWS0+4S72KDNU1NBRLSnZPqceNkikcM8etnFpZRzGCy+gw0Fv860L/3Hgx
5T9kXlo5YStAsMgT26gXyzvhxFyf5Wzza3ytt0slTIrExqwPMwz53wnaU7+BHtgQ
eWDhRRoc98bluizGW5DyTStG0iePzlgeDKTDocQ+vjQCwj+/TKgqebbQp+0lXVLt
cJjOYFUK63RAvG2xQ7m6kEJITNeOtu01XkoZtZgL8AjOh9bBIVFlOTndKrv22D7H
eArB5IP5gJGoftRS9+sQXwZLcTcRhS2pB2MPXfd+A9awVmFAbQ0oSH9oUG/w0ffb
7yu44ft2qslcWa/MdfbAanJQwWdlULB1mcp/D5JFChphdQo4vwR9NfAHEv0vx4Mc
mbJW0f17SpebHVJ2hSEbFg3ET0cxC/jexUR+A1hUkCmgh9w8lEF7EyZp0QEg/pKk
XdZhHU1YWKKzDx0iJdOIlo2uHxdla19AWRKDvXY14Ot/4+zvT2qlUWn33eT83sZy
7yDVFiOZ0WHBNrQ8wZiJZsuSb8wh1OnehIEoa/QIBa9zqgymI+kqd2IV+KvikF4H
R7LWKpCQQv4lyA/xJ8RCNJ2jPgLLWYs/6RsEMIutxFDYkVDNsEaoh/Pz3/H8SdXM
Lj2Vc4beNub8ibiSvT6gBkww/EmLgxQLGNByQ+t3cQ0xa9BRZplHVNOLtqVq/BGl
poqYMHRSstzZn9n2in/6ZOY5vtU+FiPdo6InfrTvG6C03/Rio2VyFgr2e2IfH9bo
hEHiduciXcCUP2EYuA9EJLNvivEowcHjV3zz41Uo4cNGrYwOUAlM3K3Ry6BVH8SH
Efy0ImlqSZO/Ectj6xhfy1+sM0AeezOKSJ0ThjiapOMe85cy7DGreBBUF5WC0tsd
1jMakTKg9EMhhAllFKVL/8xqUqCNEnpxba26rM7nLYFPNZEgR5UwqOXnznxZ2ipj
aTUEm6PkH/bEo5rYUY7/sZk1snCY9dzvJSq8Hy3v+wXVe1sPoFR/kXqUZF2mNKec
YTCiC72P5HEWhw3UsF4VCUcuUqtzkhEJ1KPZJ7VE8XXsR22dY9xdeB/qxvNCiLPN
6PSEfZyIbf0h2qMjjSeRE82jz4Vev3BEt9Ak0vkuvXW4UaahGPqYadUX/UXQFDe8
IgASf8wN0XPQaD8ZUuVd5wMXe1tosW3nShg1hJIAU2EnYCdnk4rFca9ufkbgI7OE
WHOufFSoE7z5O+/w/jNyt5Z5J5ggiCmiDyjl01f8oSWIs7XOvcFmyJS0ZtIlYLom
KeP0EDr5SNRdPOz3Q9QgozE1HAJpn8Yj0og+0JaHaPXtnbJ4SVGhhDSZtUhRmQ/6
/exl4JQ9jC74Uvosq0XqlfRuuezoTjqVwACYcmBNfaXbmDKi46F+DMy3+wFA+S14
jnCjDftBokmh2XmRl9Pq0z/ptru5OQ8fEMmvHzG0W/VrcXN5Yn6k0mTB9/5tN824
qigpIKbEi/kkcb6vpD8XRms+fWQCnTtLun6whT7oLJNUMU1Wm8N4SL4oUbnb2Qu+
K8aWmWgQ6zs51mafBsDWTNJqds2ojj9BY1nmD6Xq+1Vt2YRdcWJqq035cyebfflz
8DxzEtxc6Q4Ts5NQ2PniIneo/8xsma+YLSdqSeBg6HLoyxLr3ghOXezdjrG+Q2ms
xJzyoBzKneaFVYpGhXf1KbohePS6aq1nYUDvH+BASKfnvADvvGLeoq+Uy1P8QHSl
ZpR441eHgUuPjqRLkonRvwfuxHaaFNvjpOtwRphW2zewc4Ql8aMtNtPmyjmdbSYX
8VBpLApLIxcAz3uJMIU2jB8sCNgZwjssC8YtpvjW8yCm45Np5l75Ok4Tbeb1BSBc
lVgAmMYPR0fbUdE+ev73Gqi1T6Os/YU/SFBy02yTljmkQrBpVnKjLz+ELlX7iSy6
Mx1Nw70fNOS63041VKhqavuUnrY0/uLZthv1W1gNraodMaWjjPbKERYKwz4CNtIt
TWz1IuwKJCTEwn53GV/zGFeS7OwQ9E15D6J5tU5nHsu7vOpsbIs+kARW+lBBTzmz
/57RA+qRFL+gpRVLkr0B5YoMHbpiKlM3E5Iypb8BpR9dHS5QDvOA3jfxB42h4mpK
giRLbv9TMdXbGjEiL3p+ftOQ8gfpPfMUNfwWXXqOWRUXdh2IGZvudkwgkHVIUcP1
1bW6AwpPF9D6pISgqHWbElz1k10kmoGvGccYWQ0y2cxmNdOYEUPBZIslO8+urBGV
LeafySVdMf7ijbsN2Rg0FxTUEb7Bf9urPfEH3SNcFmuQzE6KyqjxGD0W7q24oO70
D8ePZ23LcKwxz4vahQBhloSopkTsxWLbPFGa/9LfWdU2cooyWLvD3YM/LLQW4Yp5
QeA/hw4e5LTcFwSHqV0cSidtjycx9J7J1vEs8ojutF7oTSGfLVUhREuimk8QqKYK
kk26i0/ybbCDSmNVi4SNOoH0E+LkrfmY+lD7lYo7/XdKZOBqtAxD2ccbYuNxhTVD
Ied9omuS6v4SQxbO+4Ifj58unZj2m1iU8X0/Dc/3DPK9iu/ecmdrn0WOIVAiDo8U
lX/j2nL3sA0MbeRvqqxijgTz9oHPLaZHWULrd5Lsc2+zxPa5/FrSgrTpL4FsP2g3
z0mifW80NBxBIvhDAy0ps8skei88KgxkC/vFM/FK8IKwE9Ibs09SRs4m9eHgA5VM
16DoVvFZJJdWnaXts/vtFqw9+pl+PpMhdUE02NOrm46ibLOyGg0sOa1pu9Ea/Hj0
M1ilfsr8IKx1MO6lu7jrcg5OKt6eGzPKeijh5SM+sFDtdAJXWZrlR+C79aGmmGLj
cwUELksK/VAyoRcuU9pyvNNGRBifYD12Y1IIfcG4tr/pdcpa8i8dpOI15Gf+cOA5
DW2A153Dw/zI6PtGs7tFUCrg+9P/JImIXWuEzZmhF1DDaAMikio7ODwMngtjOhSN
AWROhpFbCCRcdIze1i9LYohUhi2coIrYqst46meLONYdfQuh25L0YoSXVkHya8UI
mmNQc0pFOkH1uxkB6LBVPEOx7ScgX1kgVClQAslfZgTCgSYtJc1mv+eGrrq6aKZs
SNLmS1xJ5ujkbjgbJ6kKsUxKg4cBKFKzGI1CPoHnIrHgmH2c/wG16pjOSHJwK7Xb
0KzQbf8FTCiuO4X9u4kzk7CsrH9SOn2biHEDIxqKUhJf/9cgCHEvmXbYumehRWUg
s0AzfggcwFgHe0HcWDGg8NDnAR7qzWKpHlu7sNPY2mzrt1UFMS1CP3OcSiLtHvc5
MEAQGQTpiYdkgAoRRhXC7N6Xi6nV6NJ8nvp4PCqu+KErODBXDRMkMjfgJXFsS1HU
TTFyL87mE2zQ/LNJyvcWcKibq5ZooK0s9PbRAl3v8j0m1Z+SIugeI8dsTuWivkLd
nugY1U8f0golGc4gd+32PjLsRdPsz8caOAMSjJrB3riBaJAiiFBTSAluTvZL8wxT
s+sXGMh12hq8XaiLl9kk3X5nbtWrQ0o8lSyxvJ7++tQd78rY1PkwqsIYskL2gYq5
N6c4p3pHoNow3Fv5bqsAdENu7o7X2hQDy5hrEmPkOWAmDJ7H2vW4PQ3U0r9iDWO5
U+/6wi2aYI3ZkVfaFpf7xtjzX/cc3b4gbetYeNdw2algnaoOa83gNhk7Mt+PCZT/
/XBYz9POXHcwXJupgrbyTGX8vmSUTY0w/e4TLzYf/VrR4v8OaWUBW4G2/8t09kp/
33Pr3Sd+xM3PaNhJTQQeIk6d5aWZiwYb4g5QpXNsD2Q8SI2XODoQCJjqPv3nSqZE
IT0f5m5nsuykxADywuuOyp/xX3iQMAUS/OLFeeBy3xf6jIms4nsRwNB0hcyGAOK2
aFsi4QYq7cnHpXUOCD8UDWJNnmWEV7wYQj1JsHY1iz2Y/fGe0KFme4YxBYp6FeZc
Qsv8CnhVRjPynwooHc3tmqEOqBXAgLpCGe/dXTJiba65inHapWshF06gHa59g3ZS
lJmiwB4V1+BBbO8oFPSBq0c2HP4WvlZMYDKVDruFx2XwVx4vJd0If6mAbeNRO5VD
HAgljj1SMKT00tPAvS8apQXjJxgyP8ulReMeWStLE3QBH1/dSpLVMG1EjefvzJF3
/JajGDg9AGJ6UdIFWUcvL+yCy5yV2hTfHa1oaJkhGMUZpnh8MMUS36XdXF5cbWS6
LH6RMjL0ef3XF4MAkA6LdYiAJVnoob3fwT1Q7PDtnVpe+gHyV7ij0OpOs2cAApF6
e94iB2AUHR35kBmAIsqfJVT/RlQsERT9294MlqnVG9+HIKrgg2XzQxUZ7o0Xfqjo
z4oeXOnq52gzJ/8VxBOdOgsD5RZohsoRzunGBKE8REz77SItRwEAQChJqoV7k5ES
WJUfEzAG7qvNvEIV/BLW8+qBE0D7Sd334Nx6vmYCCv+X0A9z8RBCxR50R1PT8amW
T/LXl+xGCsoEMbF4RQRDRSJKKuVgzx1575q/O2p7iCldh9/unevPC11euuRfCThq
8e9c75pklfvbJILFnchbDpMCKcWW5n6ZYOfu28MZHvog3J+0Jq5qqVwlU5V3pVDz
kzcb9r6xpo8GfEe8nth6YkYd32ykQsZetSRhRwsFA+RKsl6B1LzPWH82vHX3KBUH
53xRkIBlsgE/WfyDR1TDaJz/OZTkJfFWPZ9G44ZB4M9WwmvL4AaV/+ZoINpV59UO
nWmuFl/y2Ev5AX98B0eFDlZ8WiOoSpAmTvSXolL386NQ1gb5mPXKgAYJooV2TlhC
cGipJW5DDdNGe3Mt7169jSIQSCWUGXh185m6MXHkJ3fyogOGWKItOciQ8n8v/1d1
4rEJX2TGvHGKvWIOYIl93q0ZGMFXUIVEZRVbETXfZFc31kr1dBOG0D/+oa3V7KfL
CEVHBE3LoklmLI0wUGIiV5TfoVshrMVPC+T7HbqwsCJ/Tu+NLWswJwHhkQcbaKl1
zIc7MzReQO0le2pVHgAF3D+6EBfE6KcET3ZDwxQdbBhM8dmHQ6QvB82FZUf5AV3G
GG8afWzWjvpjxfpiZwFH42mz98JzFUjjGhzBnsQn5g0SYAPgHMKqISy/yPkxenEz
Mn9rsrrXgoUPj4ZTALxtBElXKTUub3IrfnOEnoNpKmvcngmTFMsTiNDfdADhYR2Z
o6VtxAZ8ov4ykjxXciu2BenjzvgCVfomzTHwiNbFKZwYTgIRFZTFx0cXpn+eDUL9
SrvwMh+6L86mgab1s4z1qOoXw9BL5bjz7Bk0YSbj57wBb9pAtAmI6RXBE12/Hv8t
STklEuWivxy3bHGShPbvRFOZo6F2+1jWxWn/6aLK/73Tp5Ld8DI0xZnSOkm5Ziaq
JgM3fkYeGfY701I+cbSfcCPhU4VUDAqxdAgH8waCRPZHhyfaWCfIE2faJZMcMIOB
39wsHVy1ZgbxIJlWeCN4YQtOsZzMDKDaehMjhbeA/D13WUB3vEjsIPRWH2+kqmUx
ucy8C9oAOnwUsRg4q8SR38JCjfveiIw327mP9mQjuyHG4dNm0On+IiTYlgq6qHzv
yGp/B46KuZZhq/bKezRwwHzry60ea73SqkGTJj+OX102YecfG1bG71HcLcocF22v
vXgFExLQGKMrUCtEhBhMzxN1pv/wCNBTrLkJ5VHOgfijR09Liuo8y54dyNqgnxF6
5MyHDwFsZDILo9FuMoEB2nquPOXBohXpVYvBOBXXiG8bVx5dbOkMJSDTotlN5hxM
rPXEWcqAjTlEktSlvhaFlvWQeRJdU7Ogz+53tfmtDhuel0emgluGhVBBSto1GoOj
+85Qc5fqHFZW/Vzqf+lOFYVwZbXD7MoN2f43FFkQtCKTWaBM7qSbOZQuDptkoxGL
X3g1HMm0z6Wqs7vmnEkQ66IDUuEokFbH5BXnAkC5L/t2OihR9XdSDiOK9cFsHGev
O6KlOL7kuuM+Y6ka7qq26suuJ3VOXoznoEk1PDSuWzQ1+AYp92wEROs77nrlIsVM
w9UfHprVF3s9yPhhyo/TiEmnqMh0TVhXY9pqE/GB8fYqD72w9O+0lmSdCS9/1A+r
wwvXfdxa0kUKCwzWDP5RlsCl/vAsDo+ZTuY+yKsSQgPZPQZIli7cvubn494xw3Uz
MsV9alM3jjHAOJYWDAWjJB+5dSzykF6c3I6lNCHIIBy7EgV0+Drg20+Ph3Y7Ulag
i8ZuzJn0H+aeFMz8DMkE+M0adpIIVBchUzM5LBinv2G2tS/FTq8zNE/895ES6Y30
EVc/D9hc2doexELcYSFkrb214ObFu82TjvaFkfeTF3WQpvqIUHH3p6GsOAcHqeT+
KlR+hdYkBuL3Bz7AHBO2401DsWSPn9IGb6v00EihiYcGPPdaUf6X+s461CmF4UIY
J4mp7ub6HfJFNky9lx2Cgw8TRIQyhq1SqxePlJYSgwwjjbvF9VYKsPoJT30Ilxpf
oA3iz17IFijxBE+uAfioP3uF0P2JutCrolSphIBE+OJWuCDRcC525EocQDO/iQPS
nA4aPCjdbttvUYQJOkZ1+DC1uMvCvS+SblesB/wWqDRvdEU93HoZXxfJA05L90Sz
N2KMqjW/tRraF7y4dF7upYFbsr4exu3nJOj/SVLAGo4ldE+kxM2CQhujyfQxKGsr
rjfEPLS4VVgnR5AGm2dqF6rI8Mew8+J3CQEESotOOMDVucD21FJ9e24+ruiiDSp7
rK7MUS0zolTJbtXVmM5IfliToEh18+xtugA5JspmNSJ9oPvXO2kv7Hfkppu24KgX
Rso8tLgvYaf814oMOF7CEprQuOPkcKsfQVnPZe0h/XeMc7/FpgN909DORoMYyR/7
BLdssDpBzyyNjXF7Ts0KvYOLrIRpgxyYHL/FakTOtXXcWpfitf46Hft/A30sC+Ev
jyRe70Hc93GO7cK5H8WepQKTyjzqSMiHF3BrsMt7g5mkuB0xQPs0r1us2zx21MIa
fPikHkmllNcPonfWTEDY4RIVv9oaR95uUmqXCWvMatHc0IzzKDd1KPRcY6J4Lp8o
0SwVDt1odNBGweL0zjrupwRA23fVopKXNCP4bqraGLQN7pxcljTgVHE2CFXbjBuo
ZS+JA4SPRf2RyNqnH5HJj6UM2vUOxqgXmIVne3JzEIGuAlpGbJWNabOvvsh0ONse
l0Ufk+38/YO5ot522RYusO3E8WAsb3JEIJYcdw4+hJykQmBhYTYOEthqu3/iolkl
DmuXiAZGdacw5ZrNub3AzQ2mxL27pauTIVCyj/ogIFCFcc/Vm0ggOLBk2pxQzV53
QSDXbM0V5GMFjZsnO+yUXqeDNt/b0iH09gNuzQiaDlrz4s6jcf2uNB+aPHHcSDuC
DSdCfFwb7xDehfEiEk99cV8+JMkQTaFYV4fW10ApvJvC/NIi/FLHzX9kmz5/uPl7
EmWrghzXhAmufMvWonYRJ+aDG0TRcg3QwEF+4Zo0PiB7W7A2BqB/BPL/AOUIoSgB
rPCzoiR06wIYktJx6Mo2Pr/Nrj9YHdNB0wY5ipk4TSgqb7XNbT5UYPLapVZ6cpkw
/Sjn7mfxrbewTpBXGYJKn0Ib09r0jw/2ZYv7uiR443CIigq3R3K3I+G8EaoCxNoR
pRwMDylRXqvG3E+aS4bysfx0V0qBZXQEPlXqlUk35eQPjYnoeyRvAO/r8OhAJqdd
rSUtWlVgQ1fpdoDPgndUArK3R5N6YINXNfPORndhcCAJh9GFfOsVvMhIGgRERJeN
oxV/SY29e5dvKKeJAXD7LjsODhfI0mMCNCdam8awXIUxDLb1MCIyaQbXxWDMoMnA
87UVWOOHq5VBeVVCKf15bQvFgKr1ZOXLxDRaOL+G4dPZDMfuiOwgdDlcoJncbCCy
TGPFtvEpnTAuqWpnr9BphnnuKR5S26h0SsooKWUExVWr1r3nBlle2o3w4Yitr9IT
knktWqBSIzaq3+CXViY127J2Ywe3TwG7Y6chWO9KngbiaS4gj6lnABIVIEe6x9YO
DdqLMxMrgzPdgIz+97DDZ7tyofgdDWYVsH1Y9LQeIU2jrp4eEt72pXZC1cfiQ5yP
71Vk4HnBNlviEBGbiOJUDzQ5BIbGVYUU+0YCAY3N9jqAY68kDHqotbnMOzO9XAIT
wddJvIJWJsQ9p3ZzSaxPgriZEKYpnrnZxF+l1MLiR//HpiC8W1g6m/3EP0iyQroI
J2Lgh1Y5qqnO8zGhygJhP6whfoFXc7956DuoSPAYNA9k5pahHAj1N0ExH4Z0ChYU
FKwVfxa51Ht1xZh16x9tNU5gK77B7E4OLQD4sS4PgwLW1OIHSRPPpBC/S1DiHRW1
2pfONhLhM4AG//gCg8LhYxxvWjfCycYd4jsw2CJFZQSsBAUkIB/9iRiEzpJvvPoN
KUoRLqOaeFop7IR4jzsicB/2bQzE0P6BOcHaGRkZcWq2MO89ymezRXOkFFDaj+2T
tPxcfUiRtbk3sI7uex43Yb5aPPKW3+MSfaQmqsdt8aEjbY77cL2F0uPC/79Qt5Tt
KrpjgHrokS/jCGAoUrrpuju9ppk+SPyLdA4I2A0gHjizPn7x+obE69Y3s+nMsNPg
+9Ilo+x2thgUwrtryRU5AOYRoSjK3z0vDfTqSuJg6IWPnfoKMDgbCUMyL8GOUeyY
+CZa3SGvhuz5uzJlT8uzsqUJl/H5MxHlt/mzxf3fZdu7nrvNI/eT32qtFbi/Xszf
IKoPQoBrbd2DniKhvat16uKJNn4+akUujGoOdTsleGY3cXh8qAL+03vmlKsTkRSi
fyItgQ/7Qza2/eGcuq+DLrTee+/KUMTStUKJANURlwxOXYpLBpiiMHp9XWeAfySm
Lmlj3076BVB0ljKqU8n6LFp/VdBKgQHD/RZBbVRii5DxlauS4elgeAC41s2ZI9JV
e/9jdS/iNnpkrrkZ8GzNvDqF0DG8L0JKAaDGLa4S5Sb3ZMl9m6XjHB/uv6HWcgky
rJpBeUQIV7mrV7Fp0o6BLgYTQX0eKB1F/qj+N6Gagd9fD/mw0uPhOtZDeWDSspRv
wTEQlVVwJu/Rl4HSv50C0GzlXsXTHh6z8gVu0x+kRchPngsrgzns4kQKOUj+oWyg
jUmlu/zfr1DyrWgkoivyOGSvhNx5eiRbr8bTuqWFOrNiM78mb4oBoGdzleEqMtCc
cTwtLa/xU2kphDb8p6mmtCam4VVTLZaUgtcZ79NF1yxGYwFRWXsY1k09ezfqD63N
GhiT1GD3xPxejARETKJ3c8EnSD50gsz98lCiUNylGoH39ApcWGRWuDl82cAfZ0p6
cGVSGtXmZXgwosFmK2Cy0H9IgCGALZIuW65xgE4HrzrNgyIPIEh5yb2NO6l7H7tG
HNgbd/HtP2uRiPZK3FxxNz+WV3tmW98Eg5Qa/0GtSkUpyZGUYVT8GudSUgxn9BCc
rI5fD335eTsOWYsNHAi7hEmADS55sd+2/jLa/Whf7lEznxQUrL428By936hMRHtV
lcHdAyw2vTK4URgyy8rftLc8d3fQ71AyVH0lX0+eBsLBrW9l6zeN6+shG8TwwR1V
Enlt4pumMgVv/ZOnwZdWZAlbbyYcrb8i+NMtS4jiYX/CJWN9On/O3cBIR1TaA8cZ
gwQsJn7D8tUOMxyXVRmueLgexqaES5CUffIDYSOhOhbvVu7dnI7J/53WMzw+5q2u
NzfMENimIF42VlM3yOB8WhiyywZktxNMYSVso9kSt+wP/d+8Kpncin1Z1ECldbyk
Tx4gla9miR1O1muJFg3ySoPtv2FqdaGloz27oiJPeXgpI7x6v3XbRX1gTqthbO9r
YfRvIp+YCstHeOfriU/RdViZNA3901rTSTlWUVR566r5BAkY6THPvImUmii8zCbA
AMH0UKntXjBkIuUm6UIFHX7Lr6xyCScoVHOCqWfNNbNWDpcKaroZHSPXXX6rxS26
8N5aFvzwiQc4YpQ8SSx/h9hLCahmgg2lfLORu8rUt2ky7+Oc3lrX6pX9Fk3r/ecB
pEVV56UkJGxh3KEiALc50JLLZmgfvn0s3hP6Ra2/8AUDcH5INdl37AJCWEpOapcH
ARvzI6SoeQAZqdSyWp4i0YA7Urq6aE6nK6uwgsWrGh8o2wVDlwc3AV+SqVfk0tSD
02di54V5m9tEmnsOSfsAgLCf6Ia+cDiFIDq6DNXQ36FnI9TuBNM9z9Kbw64sy8Ms
pOBBeYneDUz6IV+dgH9axBGdbpDsYduOJYCDMkyCdpx7P0uGWixw7rwLHp6/3pnN
J1o89g3nX2D7Y+V56tJgsQaZWfMHk8hgUfFapJhLD9xzcMBRINJelW6WPwJz3U5F
61UWoWA29C6jqZ9k1wTVQgwNEcfD87J68s9ZwxpDDGxywyNS1rxzNtp2ykujHTZq
0l7WRBy2j+wH2zy+pQLcXa6je4yNxOppysdbIxm5LQRKos9IKIEztR8RQ4psuc9I
fw9DmrchQBJOlYc7Jux8wsUyY38b4qnBQk2iT+90gnm/kYXns+L2coAuXHrRJoph
QV1Hc+ejPihuiYxYp0slbQs7mcC92XRLQZ+ITLZ864KCrULaG3Ktke8XnhIcIcYP
B+ubfl2jGo49c1ddqUsahOits0tg/fonp0WlBv4oxtqmtoBsmjkuvSe0cbr40lPJ
mW/rTzwgY8TzGxDN/U0Q0f8w6gyk88gbLpA7eCXXl4RAMlvXTRXx8t/CPKbR6Vvc
kQ7MHxkBbTAPAjVnMxdMuY0xCzQp0fsj/WEubO1qwspLRD/ZjvEQxLik/wHyonCW
SA7reCo58O7Qy8oKhwIrwIpO24zxzHP/OOBFG2/4+Of+3J1RAwI8bk1CBUl16kT4
b+7lWQVy1QtiGu2owJ4OJuibqCo5l4DL5xkVz9Vrzdp9o0pZp6HBSz2eGMDx5F5j
PsF0wRYPjRTG7UIjpgYPBM+CbmI75Wnt/cE/H8dAy8eP3dxH6/vLn5TmV0mXZIPW
iryn4J41nkfltz+8+M17KNlVV8Xw9cFp//QkCfptcnwXihvLwbNX4VaunG0E4TaD
d2ioXqEU+lYnu7YB9kDXaXCes58COpFjDEp1FDH1P3tBgw4JiINHJdJ0wb9629q8
HzyN5pHffDuTzhSICETm9AhX95ptMPWzPxdbSbLfsqnKQ4+06lw7FhqASLtodGa1
5Dam8Xv6cAJb+wN36EDf1zgHRTLLhDZwatAZHuVnpsPbl70CDvppWVq6iSZrmSht
IY09I8OJYoq9PrslcS0bz0DDLMde/G+lOczX/pyCNuF1oRJELZYUC3X9vKTfZJEX
vX9X341N5PKGHnH/x8v7phDX2qFFc3/MEJ8O4WgogRqBJEnL9Ojla1/I7K2g/xEw
pS+Z6yrMujrUQcLGAw+OlR/Ndqnjl4Hofm5Md413eI2W8idRK+3ijL6TZUocCu38
hUc/zdyvqWSuYCsW3ywqMTX7pQEO5gJX8ZPxXDlDap6fSb0t9tu0pofklpsmDGtC
nqiyI+gyIkkkPLUDOr4cUhzQxO3e79EqBKhZMjFslD3aV0TU2pXL7/CmmLMa4h1u
MnGsogJE8kVOBbiv64m7oo/sI1H73n2GVNwGON2rLVNZ91agJr9JW//WKzvOiVsB
/0e5KEQ1co4+OhwyHI5LHkTQ4wPzYJhs4guw8zMnBEN8wERH/Q0+YMpZwoqovSmU
av5yJ8/HCzDrRhsP441YQiDJ/hsCm/RZB2oWWPULc4MRSAjHiz38AVgePWbJcgdK
BK6Xuf7DCcskbkhSJgCMsft+tdOT6ID5wdbXqNj0pvrz6oPWGJB+mpUS+VDCnOkl
eFaXb7NdqaTaUfDGOdiPCh/FTwLH5xZZHhUDzR9jQecuTLOFup0EnHxPoesLlvkl
pamhGVHXgMNXT/2MjRumke9kWA2iGOmfxFJnEi8pKNp5L44bMiTF+kwGZIYAV+GX
da7Z72bkAwSq0C0umnCvv2nWA5RFf+UM1iodEQvEq+nZF3/tZ43XTuP1X00oB2kM
eTlAquXB332M1SIupS0/qBuWtWhpTIeJsjmihdEiAeyQqnnvvlzraC2Ae3v5ubCp
vlorgLZEpN468C3lKFpp0vhyQ6JfV9a7oj3ipke97rTt0gSNZok6I0Wzi4p7pT00
yJ/n+kG6g/la5ED7QXQWuykLez1bTOGpSFfck5PEnQAZQKcMvdT+aT/qXxSdKsHH
SxLZ4Jzcx9WxB34UST9w7gAZ8onS4/wxlzTTLQL5x+M7cs81chwc2eChmgpwOapX
1/LaoadyOm2e9v8Yq9BUONXXLvrCmVO32b9N/uVQLGSkqrb6wokO7zebPs7DIk/f
O+7P7xLkQ2Xb98ldUXG3srCR8y8k8FJcpJfFe9Ke0fMHQihCqOpL2ED39Svmpw5F
/hbGsHMzzZtkIFBSjR0i6BfJd2Ec/V5Uz/ss0tTfpRM2EmxtXkG1+T/LDFyf945d
jJ/Gk8Iz3rPsdtxay+fQrLofSUObAP5Hirbl7ynczbTlFIaItucEvuBClMkPlFJx
ZRxfw8DR8g0e1g9Q/ZIvjDGtHreHhFifmAkYt4TtP1e1Lh2gK8aNyT9K2Lnvhy8F
cBQt4fx8Y9dgJYp3HjbSYtMEETpa13VBX5cr0fqA4PJkJ1jevuQG2Zecge3z/zVh
VjtsJIwcbZVyQbPpxpbSh2xDK0jtsS9/VThciuSbuv4Q3RXRZ+kaXopxRZZZYYoJ
/Z0h531eixqycYtrYgEjv6mkfqdvLgQEAMvnCj+SF6p3J3omk5F5WqvgK4fITEvR
Xew5ZBXdyUWQMZpl2vtownGqv5rgH4drBsCfJ9toaH+GfdmHB15j5Q1byWi4EVrA
vZLN2Vnnms70i/MfuRyRqn8L5QyUIW1kZ37UnDBWDC0RvMLzk8Is6Ix9zj/Pp/pM
mWt7g2eb9T/AxgBE4BEZpVYnFekyIcYPJdMp8ugf/b/E/YTkvnI4NXlO3vhvioEz
Gkv4HKQx8LmLRE8NLn4LHBxSg0hzGQFjRzaJMF0uRYbxuchTtDaaUox+CNcOTK2j
0fH03wMxr464BOU5G63ECUcgoJUdvS5bLkCnuLUIyodq0ygnS7y0SwBJcEaojB3J
Idw0KvRtZgtMa/5K05v2uDWRkU94CyV6EYd927bow/Y/p+KJYjEejW5PiGwzYS73
iPyCvaQdUHcEYbtNfDX+VrSIZtYX0+CcJToON8AK985uaqTcqMSEzpuqVC5bUv3b
aDOUQWvx2KLTHY8Y0MFJ7wggKI1oy4uPjI86jqW7JBvE4ZPGmujhinslsc/CY4xe
JjIlaY6g7HeINKBssgIDROpirdlgj2/LgN00HR9BX3Rx+3e5rC3Csq2Y6SqPTmWO
Be4qM3AfxDEn0QkmqG7E2WvtmtPJ8mecSofnTLowk8AXnsmnqOuO25QA3XoRaCvW
/GugLzZ5nq967Z9bKlqZykp9jfelDcLi40Z2VTbX8gQ76RGSAeLzLDCOLR+s4waE
EL0O9vAOxypmG6mvJc6l85n2C7Y5mRNPaA7RdnFMLQBdVC+tOCtDsc1z5i5Kt3KA
7O3NJSuPZdHtDCelb73DYp/6rAIcnRLgNSNJ4IXkqBIByofjqqEnN850KgC8yuks
ZXzqf2gQNQOesfyPoGz8aUAg375uXzvfysc2EzWTyrcjXd4V2ALU4Geokj0/clZm
iIYdjjl34+6gKZVarfUXAVyopGjP7svL3zo3dMaepOpFkKP2HiZtBp39lmd80BcE
eN7kBER9G0Pvy7/66nZRYn+jkDBWa0kWV2rqKcvMyMaNmH6A+c+FHn0J2Kj8fsyV
nuGHRXWmt6dZns7sM7d0GIV9y5sVWW6PuOMtc1QvR37+B25vXDGKeuMxronxhqK0
oY5VOQmrHfPpirCEzJ4L1ru0LtgRvpw5NBwx8tG+GrimN1nty+03iEb7C7qI+E4N
f31FaaobXXeFRU8TwPqyceKzrIzcWAlVBKe55cK86m3N1gW5uaHwiBrINILiWD/w
gq+Exv91LDMPwishKlL5G2kZ5zBWpw0G9wSoKro01218jpCkyFKQS41MR9JV0/YX
aRdwWxqd4xqUnKvogJOFm5gHpqwHJ6bz1pPl71MRYVFI6DXt/BQtnXhcGpMVccfE
9mLIzh5RJZESxfh2ajk64GgXNXIwnTWHWB30MhlXo133VszL/zDU8Vqyeki/3PDp
qIQQp4KSELdq+Xe2hmkVL+ZsZt6qVtzfj9Kw0c8wTzmbMhNm2tao2kmegQ4TOW8P
/yzV2V/9gbWJgyGPpLQNU9HDlercjcVOWlql4Vm2BQ42edHiBCqcwhlO12u/xEAj
ksMgUAWeOj+nyLvcqSIrj2wutd6knyNP4AAofqPZO+lCDQefi8zOl0IjCk1FG+G3
y6R/oHHT7MSwjapQ1N/1emR/6ZWch8NaVEc4aG8jNyU5wFb8VA89aZECtTe4gEJE
hn7YUVu43qJzhJTbiGqxe+GxmUo1z7Xmi3iSfTDTmOkLEkC5/kXOYrcfHNhfTNfb
VQDcJYRpd+IEVXd+FpcceFIun7auD7ZdDFJGFG41U/w8b5O2PR0URaZGA0xAFEZS
ZQxDG0anCD5iUv7xm564bWdacXa6EmWsVuV22EhwNumCmhNZvll1k1opMX1vHTos
sCc1HGBdi1xYOVIKToXdJosSSHC1Jx0BicfSOzIYLpAGEBgZKr2g5Av0NLT7FAQa
syd9wRajkkVOduMj+FpJZ4fHdAL5e/Cg6G7yunqO99qXLCk/SZWDFGOC1yUvczXy
CWctjZzsZ8cUTYKwVD5z5JuuHqzGVRs6TlCPG3vKShDIpXXg9gzx9eQMmH3ANvcg
DtrQFqLAGKyJHQpyNIBWUDr9iUQUuN5NbuUmPIXc5kjSRdlF7UEDT6s9P2awQiNJ
CqWe5JNAgfDG8Wp9Jau3Gc8sDo92ILZ9CE5u58yrCHJUUo4DNGy/SxUJr8MprDNk
g4/MGyntWfmoH8vJjAf+kyB2wCTvIDEqLkuHTiBvlMggdq1QK0D/2dYYeTV/M6Yc
opriJYV5n5hIFdD6+Sp0wVLVQ/bqXp4v+XhFhSRb3V8XDzAwI+rJP8HXuEEwyWTF
wWDaDjWld8Fkx6GnRslp4DBCJ6iv/YS1b3IgWn7HE/nNTvkgIVrxfKSVAIupoE3/
UhOsJw/xuxgD2hekORUBJYlYcTBmp6U/ZiCRllBhfkkemq/L8OwL4uck1fhyS3jU
jEROxxC1jaaCW6KWS3ED8Y48c3GqeAbekWQHBT4OMiuBm2mK67koebL1/uRJi1E6
jNymW3Tlw/GyXYrxLkjjz7ROtNysssGJF5G2CMxeFKDoZFrqfoWQgy326qfdYX3U
JjsaJ6VpnRxGwx0z1wCH9XgvWT8mum2l8xb/2G/Uti2AE6MDrlK2i66JQo5ugFf6
O0c6QIxIKlsB3wYfeaCpLvSODrnN2iUvYxHdHA+gWSdhQuw5YYqGCZ3wXDY7RVvo
8X8ocsV9njfnGNmlbmqLAo9PbZGwBTG3xzk6NyRHlaZqAP/ldPXrejesCQXGYi+J
L++MOO5K0IRkKCIsw7xIxqjFiU4AWfDVIKyoGmB4GpshuW46s8s4XJiAnfmTjDMD
xQXRkZ1fVr2m9i9kHJMQzIuGM9Qi9gJhopjlT4tBbtN2nfl0yGrLScsPr8lpC6hy
EuRjxeUKMZISsHWgDS/12gwSER6IxwoZIcdEYius573fuztUcG1m9nxvx2ihPoa0
kDbEr5tW7j5Gfbwh+7K//uWGGrGY/Kr/qEQSOBAjETn0CAv4aICV6tnN7jeH6GtP
0s8cBgX+pSI+s5YkAPL/0i+j3B4DQgDMvdjnLwCbNuYnlEy67g4x1lRVqBvDyrG9
nDboXK3khJSvu64BhB9tSscSN4naklgTuCeMKiUiCDdKM/jRD7QlpdIHmxbDFDRR
65GhS32COBW5G/vI3BDwD20bPpxDmPlYaNA5yJnapUUYOLJNKUpoOk2J9rWPXARw
dGv4Cppmo/IEdJG7Mu3e5BNvISRCNi3hea4j46vCaUrlVEkROXte7QRNRvziWUOT
+XzrFlzHfMUTwowuzpGmcAsNARqGSNAjBaHsd6CV4Jm8z1DtW4Urj2rswQCMeQca
cPWOPeDgRkenG/5CgmxxmfDDtalQW6jZaRcUbnHj8m6ztwyiYZhKl7HU6Vc4shlZ
daVbGisRcUiP1aTf31+DDzR6buINjGWfY1TN3/FDH7E/ydPkdL5AqMAwXfOKJzch
wDV79PDOFol/e9Us89ksU44u/8UEGBGtgxtSE7z2WLotCWQSjY97mEkKBz0o1L5C
E5BDC5NkDzJAtqsHkQlCEYplPdJmg5ZREny+itkf2kat3jwFxV9tgusSkiPimU1k
i725EmEST+SDC8Oi+PNb23NPCDQiA7+eaTqZHn5wiNo826J5vi9NQAHCqiK28VlW
Ff7pgOLYaHvYI5K8u3a5gHNPFdmPtMdi3e+IyCb3YefrVpJuhen5b32noRKQWee3
AxTB+VlVWayeM45Eqvsj3FdZEkCzinPSRlKRGKI+lisiVVWqYw75KpjpFMPKfipY
LQ1NxY8KXBaKSbhV7b/MT4dnAysdoyMHa0xJzEkCAaG9zYinZ1p1CVjIh3lxvtB1
cjHFB6RC8w2OHF7r2h8XhX/O/K+8wSRvdNU+5FVD9Rs8+Uuv9vBbPBnBvNdwxZNE
667IVIpI0Pu2Qk6DwE23/WaGy3lTVzKpBTo23/22TBXnZCLw0bNLA/lyNXu1ARw4
DwvVkg7qwhQ4o/+RTxrfNXlAtIyDB6DMILDQFUNog9KIEAochH/BqnNwE2Hp16ho
Ekkg1HV7dwA/hQ8exvLJY8eTx0c6NDaK7Opx699aXzWFrnkS97bqZOHwkcOiKXhR
2K0ul+95SL2Sngyis3AqxgaRtWnm0157L2gzIGfXzDDzWPdyAHTCVbdzmKnsUlxy
KZVaJbUBhZYHtOoSDiseJxl81A+rcStg1Kzw35eTS5s0y5t6xSMOnkgbN5rvf5ZU
Pi6mGKHbidmtLlXOqJjpCFfEb5XutWWSVg/cZ1NV6LBkzimfXRJIK9zVktrbHEHf
bXLn5Qwq+IfYQZZ7r0ITso0rOlsBc8h45CRt4ciU/M4XAltiRWXOj4oFmljIzwoH
nCZrU4NdMmWPQeaaG5YK5hhc6vAP+k5+dG9TUvRxjj0HXtPTbmxbMF8wZXR88ohF
xDHUW/4Idx5YqKlt3P+MQ0zLalsSqXt27CeFlb35E5rrl2JgTyrlxsx+h1IbBoKp
9d/vgZGSjUqKW5wPbOYVyKg6JcPP06cDwlf3VBuF+/4lO93Hq6wL9z7tGXLDX5Es
EjuqzN2AsvEb3txFoHuhAGThEWeL2dkMb9KWcjp5pFoDXv/IjctidoilQRtypWs6
6Bfl25WolbUEMC5E3jQKsVUsTp/AGI8v4+dJwNzor62aDfsjn9G5cs5PeeAy10sB
ci6SGc6keS3STXVTCmbvUbguD28FQPM+Jt9k2JoNJfzTUqm2qS69eAP+fUSJ51JW
2VUzZ2iEC8X/1hdrF9tO2hTnS2Hat9caiKqRhlXeSd9Qem0f5tU0+YQCxXvKmuJO
3XJn9xDUQn6ehvcjUXRVLhxmf5Ah9XbjRZ8sn1JMc/SnYZRis6a49gqOtNomik6e
ax5dSN3hJ9OFDCFvvSSQlpWqgbD0hKlJ3AqpnQ5rxKlv7h8ljCzx8UwiSZvcBNev
4y9pQ9YHOPIZTrCQuHFOr47cHac4xJneh9Y9QpxjZJ9SNz8ufoNjiSlWUPfHUeb+
hwZxylBF5wLb2/Z5x2FCUc1Bzo0Mard39TmfuLjsL1bHUSmezUWkUF0Qubf6RHSb
ILZcuH91DK2uoxK0lStrbeEPxjTg0wUrQkxSFki4T5awvJAPrIdQagvaH6pVY3w5
Xi4V0muvWfyuUbfVwx52XuEebIjz/I5CKeYPJTe5HtF6z1zgSFh+BAe4hYhu93g3
wVVyU1xVGitN5oARvkVNuAvJzBlhnxkxkzaeCaOTwmkegx1osayNIgHXSgBleqG+
Hm7EiqeaOHeL1B9eDTPi+op24rsZV0SoNJ8+/zbE8D2btAnqDhs+P/zrNLM8OBE0
Oq8w7ertDOHJ0SwwSee2Q4M+lr2ENt+BnMC8Iv/uqlZgyLww182Eb+PszeryTgvI
0MnOaJ17e8CndN16qQzvN1JDXQhPeFmuIIP5AyqPiR+hzDElll8FWr/1HO9kLDtp
6uk3oULoZdE/W4H9TJq4rXdQ7exRaeC/zSZ0gxyfAaJJIIhfi3o3MmovfI6+fDOK
5ZIICgdFO2T/YnBAjLe6nXic1/GR/Yb2hwiCD9OH43XxHg17ASKk8QR/DPLrNMJD
Q8Q7vdIjLPTPHwE0MDVxNxcj2y60rDsR2jv72w9gxGoKyZ7psJ4dVGQCjib+pSRD
gxMGj4ajBlA4urzNeIKadm6Y29s2Uft/zziPnHBdDAwOuJb5XTw2mcQ0kwHnV0/u
JJn8Wua0Hcd+5N4SR0xhZ/jKVyLikDItbhGjj67jwEKXPTUBCrQnONLHhyyNx9Ri
9a1+6zQ0J2z0OPlqaayX3kJuUV86TJD7NYYiTfp4iM/tpN4siA22B6X0M2hMLJ6g
jszwvwNYbyeI25lXXLwaiMA/4CxKR5aRL0zrHxcxqRNod9oppNVsR2Ct4I2YPVp2
vhVvKuXw2oLd0m9lzz8lnPjqNuEfdtXOEq1r8GSn0a4queNzOYSeb22Evl6vRHZL
4RXDcImJ5/FecWvfncybPqzU0kzsR5dvVFPsUHzZh8V12NNt9R8Y6OzMfwkFGDgL
SNiJGTacz7UaHulmWJOZoxmOGWTH05NRRgCCnlADUt+mMOxyH4nL3CeDaTCVSS8T
y61M3Pjfpt9oyQS4xPg2cbWiLxxDinXsl0DKit5Pl+WSEYEo3dLTHLHj8br4s4nb
HKQTltP/8hAnOaWsQer2DC+1eHyzITBqWl4AyKBBRreGv5U2+qwN5DWahGWOJ6lx
Nb/iIZ483ts1iFVdMe7kbumlPK3xSpsixVWzjdByxXFKcqmYgoUGJGLc4Ag1jZqv
OPByYYjEifIHv4cvtPvHA0ITGiHL2KVRpauuDBfq/vaQ8v2HVE9yRtLkxjv+Fzt9
0r6pnXn4RwiUBPadi0rMkrxv9SowJ+hGzlIG9UJOPkdetzyNFk/qNpHyrm6Fcu8H
jLl6Vy3lP/7Ni7rIcdkA+0hTCZHO8YfB4jUEgurysNKUHDWnM3u8qCqAgk8n3837
j1A9ueu5rUDxMqGzrl540NBwB0DDbeMV8JsH3ZqkAJE4ELZqKxDt4vW51/WHY5VN
Nspr/l+OYxuYkik+h1qvG88dtlhyy7OXHtR37O2HfaQLi3xpU4Pc31EUqjwqqbNi
WPejH/KkhJIXQEQqZcHl8XrByLq8pQvGgRQUZuIcARM++DZ6YYU9h6ygHR9IJkSw
RQDgN2Dd3xwJgNI9uDqudF3ek7WfPDPkSwfO7/uSWJJIR7y21c7hvlYNY2iBWEM8
43rZCVRq7ZF5GHoce2KCsBMKYFHdRV84N0FVDjbGcnqg1U+FmsTzPFsaNbgm63PE
YZyLFHLly36SeNQ0OITW/V1VqKKrmBXQskAC8zQAKsHq39pReqPTd2BFseZWsrDQ
pTn3uD7sifVRwrgZ5l6h2s/hbMnadbNP7SE5URgfDiZ9RkQ048kTvvIXiy/2EPKU
Fcy1n+xiGl4B3si997DozTycrDO1YgY/gCJPIZrS5yybMzr+NzhguZsLD1RzqBZM
hTy5u5cjdZyaG4hekpTGyyBbPjGUModPGo6ITlsr5qfIRDgybsMw8pLiVMOBX4SY
z430qXkzvvvWGxF9Z/UqOFgP/5bMgG9V88Mw+TvfsT/enIuvCw4af32ZUzBB9b0Y
ZkHz4QYRR1oDiAT/QeftuzuNe1g8gUpr6UXoOjrNOv6+zGfGsRuYm5fQizgHcS37
BDY6gMMsTL8B6ipqQHVwezMwZkmxvo1N+EJvlOK/5TRp0mzk9LXNGgpjr9dBvtxW
EfLAcqWbRMU1/XN5q4AKpHeDidxiaiSiPOzLy3YbIlrfrMWCtkjDOfZ7xoJmr3nS
4E0ah9DSu5pjAr86M0+WzmsrPcMNgaW92VbPS9TzADz71n6HSe/2jr0Rpr8mGxB5
A8CVAfai7wGEkksG2sXAsz83LZIH/EvTC+qD9E14hRbas/dLxJGTwOBeHrj6KrMb
YK1tlgyiHsN0E3ri3MJWDtMHzNo/D3exE7AVCGcVYFvGgixz/0VQjq99eKaqToT5
y0ED7oMzJz/cs2gldOpRsA6CuOv2p1s5I9oyCeZSxLTvmOz+nNlHDsnRljHVkhOQ
J79QRpn7z0A4VAG8TJRqlD3nm9b8HkP0qAgiGWfIfhup9Kvu3mpvY04EDeZ69/eo
yX403hXRftD4GPVwOA2sOJgDP3DvDi2174OlOUSnlw7v6FPkanuIZleyL2XQYxmf
QflG1KRbqlriqYFbtXOQcAE5ud7YfoyQnXQg1ubGKsH8HWcBBebaT2Lw6kJSVE2m
27rMW8x1Zhs8FPPGb79NH3i9h6Sb5q2NIAOHEI9g8Lo0LqwZSNOzSQBQ+hD6KrVx
tbNW01FXsu/JnbLLgPDRL9OJfJKwUyx2w1ojeD5Jz+odGBElnfXAw161q5jJH/tr
h4kHKCB5kUGU5I5JpCmrpFLpmaEGWXzYAuqMkdzp06sFwBofLRnbDwEv47vfYDxK
peE59QkvoZzcUSrwGPKIYPkcCuJPADCdmtFFkz9L+aAavOT/byumexzfUhF3FzDR
og3Kda9YEqewAHYLNO8RG0+dzlKPavf+MaBarNFxYvhPxiXxE0ypMc2ccXKgxoxT
jm4Aw33AMWC2mCFZozqdjIe3PN76KU9il/BVlUbxBpND6nj/Iy5RGJLPpeaAlB0E
v3MT9+hE+US+bILquQwabTS8dPErZwQQDGHbGmz2BUEwWCj2K1R/7qjS0r5Y3SQS
rso+0twpFuFGG0gXMcIjZaAsjo07EJbNGCR5NIVsHjDcMuvVIw8YAAXSpWoOlutd
O8rYMA1HU3YtrX3J+Zp73A2RVzxyHVQ5A5R/wzhTcEEsxhPlUHTemmLNw740cavn
EH+k3qwU+PoHW7K8HjYnRhjVB1gxXVxx9g35X7r5MN3R7YGEGb+/EbOUvxT1xD82
IMhRoqqr6Zq/fIlpcIXQZEdzEZEaj2fxxKMckAirBIa/0WW6gr/25lbjqIqwsW+Q
G8jjoDlh1lm3WjjcP4V4iCIo1mUDqy8PGqz4ZJCEnnvv+qhJwfVvYLpGJDDcw8+R
krz9Q3L6oM527Frhu8EYwjIgwOe2M9/ARTtmy9w0QTg1mjeBE45P+KFzqHh5H7ss
ib4pSlLFL1tX9tuzPCDjqG05Ojp3PZ4+UPgtayPhfEx6vjOFP/dHvJB4IJMFt1iG
SUloVvpc1I7la9YawWdJISaSv52n4RWsCcadROphuvVEjJUyYsl+cNtZ7r1eCCD5
jktxSkxIs5CSjtTq4sWIRU9aKoXmId+dPU8Qii3g4X6No4weQJruYnQ6w3oVONw1
Uzu+0s0xFlp+CD5X1nZeoYDqNdJHNaqLZuUJNQ2vVKANw6YRBTKpuEryh9jdCJD6
KcaJR+ws9XxBjh78zhH3NnLVpF3mX+S6prhJw4eTnLJPMaC9wIXEsdNInANeDBR3
u2VwfCds53zS6x/XqMzHCC8xtLhF5BWXiat3XCj6W8vrGXAhz1QRWPHmv19gl7l8
LD3rmVwamdgaDRRS0GPiC/CiD0GaXMOPKQQL8oNMcM5VLOoCUmv7JtLLLn5J+2Os
OVxA58LPmbC9PoB/RLQI/nbG03EVpBp7Jyjh9pOYwiHffC9daEceNmem4R3PZG8w
NwpszSaqsQqB9wVC74uyoY7mQUHlthzh3yBx26eQcWH3hv438qNFDyTzlGHpP9PT
yGD61gzY081VuHmfjkK47Vf99Uq7Yi7f1aqG8aQ0TO5LboxlXyIUrxohuI32k+m7
SqaEDVmaGuPdznL5tHphAjANtylH70C44XqoOxt1I6XACM8ExuWvnXamjdi+AcZU
NnztFArHSv5oG4H9BEg7Vk9IDmDa5xptqP8rqukaYvJKsfRgKd58jRpdYebs6tL2
sR1JoDoL8MmE4ZMQzwLoKtWYgoUKvNUWhFJLAqmhSquQmBQZaWcXwj9yM47YUkgo
DErvRLUX+scR1NJA4OGsoRwSTXrs4fLXWqsgcNJ08SPUiRMrd8lBpW32B6XI7yq4
FhlQ2BnfBqRvODG+LV/5qISq+jvS7h+h/zFvZZFJSXbFc8+w15map1psokdLEj8I
KYsOdFW8DX1qpPHctJJ0rsg2CghvWtEWuxWHaelysUp9z+MgHFKEhOr3xqr3WOWC
RrxCk3XnC8LFw++E+GaP1cS1y6q1jt3fCyk9EwySSsftD7nKwgXWQtxyNN9W9gvv
OgZsXu0wyZ3gtAJ8n83vCAikdImP11VeKXQFlWJsWWxzkw1OB6wHThcB8NVRVwbB
2dxoP3w3JfmBXcmRwX3Rxe6qJfV7BLED6NEgcC8k1H8QDVYAZjKpW0VwgyxL+uC7
BDUP6VcOY6KZJHofTi84CQKCOJxKWCNbVoX1OIBgTUjia1g3zdq/EAK9o+3p0P13
WLqHxBnPADbH2gmyX2za5pcCL0GsiTkpVLJ6/HzsgRTTEw7MoVLyh4umbXKiUYlx
WOMLs1Ui/+9vSFCC6QMOpc78wRKwEaad0AoGK4U1H96ojh7PR7xHnAwHuAmG7ERk
gCQ0ilMqw6qN2isAVj+YhyDaZndiTogXIU202E3kgcmejujB7A5ewRovyzbL8eLQ
VCUS/ILXAj4Ep1N56PeROa/WTfSR95akfRbQi0+b6RD9pjsRApcY7nU/t756gnlL
/qujSQshklXV5cByHPZUtsJLAoyCWvpvdEoGPzXfHbljwenxJW5fJog/sCO3sPDH
NFDRmNnVrIUXyM+QoSD/GL3hXucNbHvxSFbuOoPpwzf2mnis/T8ZlJyiSsiFuwAH
RlcIBOTOaxHfvcDZVVgJwYIkv1bXaqPtvu1fy5rusim+X/LoY2WsU75b2Uwvk7RW
fCyrw/M3sj6fOeEHTWmaBBgEg2i8AWBN5XvGMBWiqfP+QDGB7Lmo8LJds/vk5Fl6
EwMfPfXWiw+RC3XkhhBnRRQdQ+lqb4icML36KC+XImFUneH3zOgadTjqGkKXFsgc
YaiPd9B022PTkBPHHAmO+GEt0gKEoVeF9OSTPbkEc+fibdgeijdeLJJxQUyGqHXO
QqmbrPppLTQdq5TqqsHdyrILh84RKAY4emNoz3BUyuwQGU5TC5+vXSt80/8v7Aj7
QLISrV/pIZF2UrziLpSb/Bbk1nNufD9TOXkpyIiIN6pxyki3cOILOuJ5uYrsldeY
Ob0T1t/xWQcGhV23tvrNefl4/Cr4sP+0UwkS5P7YByVfujHNg1Loazd1JRFP4YWQ
yObQNHz0P0/O0gsIPN9m/DWgP8rpMtoGCsJ9LbauFXPh59o2sCiPwD9yPe3MLSeP
fdPOKW9DiEpdthiUs6bvmxv1BWXh5HMKISuUFcPNsFSpy5I9v9vUAjzI7xMyrP07
gnuUOncwQwqApbNFkd4zSHcXzh/IPLIFlE45Qfl3T5ETN0B0qFISPmtVu+YwSy8o
0Ny/PTikUwYDeshMlgXY93Qo0kINsN4qWAnASMEwd+5VZHjdCB5xRffA2lfC+GXq
jQDNQWi029t1gxxo2zI9v1nIpBlBiZG0hamJLYbEON88ZxMgn8br5+2VkifoIWwQ
8VC71idbI+pcGZtGrbI7HkifWPok5QPhp/GE1kG1Py0uyO97dj10CHrr8eiyBoE/
UpgrhSRKphYDinu28nJ2HahF/KunTODuH6V0V8ToPyDAgOVykCYJkivn3+8JkH7k
+HByvu1LjStB1tcaJDc/Maz2LdkYkza+lVLD0BTwfRwIStH/CowWlWNe1CUbLgXO
NkfPfh6yQZXC8YT3+FXoCo2uEXv8DTRVaQtAvYERgyhwlmaDOj1R+bd3mKKqtXhD
WBvlyrQ8RCWgOvaHC52sXJIaCTvmhY9C7rBTU/fdVk+p1uXRdFn2A5fu7xMYDsli
czb6uaUpQs59DlxSDJaBFamjx+RG0xLPHZx5T4MGSCCtUl/XbT+OzDgGqzHjoBvm
sGO7GhKj3x/tC7KXhZ7pEsPliC0EXBRdxiRdl1Ft60WTGkk+dNN6JV3wAsOjWmB2
Xgjsy3q7xnIiNNLlFOA3RijQkJ/lNtA3dTaQb5ddDtNqZkJtso9Hj0NMDwH9SVbe
BRMq3v0mpOWvb8ss9DQ8PUIx2kmUhl9dhWetWtZCBZdG2GoNMcaWZyuyyBCHGpuH
JxJtIzoBlL6hH7nd7H06qaHEDV7HFxtgKCp+vuIgdCU5qYIdFldPu4hR6/8YExJe
GIHGvoZLCKZgNl8zop5iuyg3DyoUGA0Vx0bs4pGhyU9yCODenWGyxPOGQs1vCead
itSlhfO26pA3Xs0yzdFvodJe/RIq+gJqhUyR7K4F0UR92WKWbrx5SICdSY6znl2a
5xor++vmJd6BokZunClfCjMzim1sIde8JJBNMuDTltD882viUg892swA2GqhE7lw
gnFtmeBiJev87RpBUsAp0FCtgKIGFzGGLRPCifpA5Vd3e4ivW4F+xyTfKkyVzAsC
t6pyqeR/7P8T2uE1H4k5Ofyd5DY02l0IVuCxuCZrWKr9x8wJvbz2D0HELrVOdqSO
AQm40faTIGS7ZqGUABLaTinPOkbWvu2K9JCigDh0healvUNI8SWsvn+MvZBYVbUn
011NWyraXd7JjrSktIyq79E5yFiiCU0NfmZty520+uZQ8Ngnl4rwK+e3QwfslEzj
aJ5vgqOT7jVJhymWgdw3wHZuuDGYRRTVDPTSSkJL+JyXuwFg2kQA1k5G2NQIm8D7
BNwU6H6VVEdRYQGqBMQAdhavzcYyzcw0awoRa9AMKH4zHashXKJ8DpUpNFv+xDS+
0NJUKZ5r0aj6iWZRTBAWuPCPAzT4SygjVytGwmoyINNVBzOLHkiYMUZ+ziUtVaYD
a7aQmzia6UODsiChS+EiLlIFloMgsGHehUx1MxohnDUUAelL0ENKKxGzmFGxMS7U
4J6giRb6WHuophflROiBA0VX551ZzIHL0ESukcMwKbg0Rq/PfXBtJIJUaD6asS2k
PchWQIXKDpExeW2XqjAlm2qYUmdKNw3Szxp8CnLMxZgleFt5til0WvHkhPX15rXg
2RRqNmKPHeha+t36rJ/gDyepj+1OICk8xDsehlGG2uEl7PKO7gKmwN2oORhcoiZP
HEMvmbjw6krckGazH9lf39eNBscUlwdLeSxMkOxKs6BFBUVlS/UyNpt1OqClJtRF
tsymSjfmiZ1O8/E3hDi5o5238vOgd/+Kh77GW+vUuR8G08Qit6n818cUrozWrYHE
JZstga5rRZSbLbS0rZd+Saw4ky6/bvhC58LOZwd6KXnn3m+9Hd12//sWXf8mdOWC
eTuK0hJw7buurnrs8Ta77KHIrdF9B2QsHx4M0FABg8jAZ0kjIMVp6t3c25Be7DUU
jkdfIhOYdIU5Yx28TkAPcpP4eVIFSy1ycOC1cHcLY62vQRarj4bCvMKVJZpzdKWV
VvIwElrZHzpZ5iclZrA83L2P7gPLA/+tjRA8rxml4yM8R+mfRdVyczmCLZbjogmL
uYCCgtLBrB21LsGv9rmgv6yoEN4FUlUQMrlewN0TPAsDlJQax152+EJD4cWXIFNb
BG0L2K8DQXuzTvv5JPn0kZFi5NJ80T5jDJ+x3GMLzMeGA/+VFHVt8VWtK+H/C/9A
RHomcJSvTFgyzA6W/VXGCAVVKHwu2sTIPCHilt0lIjXxddTbiPwV77PyZdkiHJTP
8ztRtP43GbouRYOdN6IIRBLObujY6aQ48cvkMiUyp0KPDsraeujk26tXJuG6bjLy
JFOCpNyl02cDREh07WHo4/Xqv+BVc+1IJrq19E8c6G8WB6sh/cJVHDHgLWWywb8r
J8OVZhAraai/MfZHiojJc7DSsaQTvBZffZsEeVq4O69mxyEXXSIL5PYtFxckOGwm
V4HVxIpIvB56EpSFahZH9ZXjv85fX/L6rt7qGIHEPL6PFqnaa5pfs3yu/TQUpcHF
lsur+o427N8SQC5Bi/qM7W6vWxRSf+MCdtjP1M285gq34w4KZm5uHTsemwRz36uM
mZUy/Z5j9UxrzhbrxMluM5DM8dU6Bs0wCNgGtmpX8OZiD+Z6nccqmOCy+qOrxtFN
5II0xZIRBje2RlRx9nvkDNVG1o7dmYZz5Bs/uWSnawhSBKKuzeeEUAqzqfQi2m07
MzD2d1gaSQcCr8hbwPS4cNmpG8n5oONqMWG6Ejq2U/mDwM6wkJtV+yyu4TzWy78r
aHtUwXSiqaULNZikdwno6FBJjxlNFbDr+OmqDC8Wpzey9Gy7IFVYsZaSyRQ7yCYG
ixucp6y0WaKsSVmgcPvqtHxohP9zqqy4Ajbce6Arbdm6bnNbctJMhE+Rys1XPLkj
mWwnaBSve1qPL32ZJDn3Lb3CBArGdPOuTWSmiLtz9JN4nW1HCrC8tThTJlkA9Z0A
0c9ZSPciTJn1AJK9UKzAFP8kCOS/XIKgjgNRSUPdzSzLkuIDSw4YewNew+BmgZGw
EUmduYAy1TF1nk/SZsA1lmy3F9FiaFpi4IGt2FD2TA0mDoKqAqK9d0fELEwxqFlg
ioCeMUjxd30arw/5eaNf+1BfKb6qaQzJRW/xqga39g6SVeLzcrpc/wpJNLQ9xQMa
Mm54NkwR6B/cFDuAt5L/QXunyHQQFhHzRS7kXbJ7ORgZbOKx1IlrXJmTG0qPEsC8
2SeJHhzd/WgFR1GrvdKsHlPnfGeawoeUyBnMc+CuquGojascNQZGGVXpELn1wH4y
xSLbB2gYweSRnrqOvlgE22EnOobComyS8ZG3GV9cfdE9h84ydq1O5jc+YYEy/5N0
dLw6naZ037WEw875Il1V6ToV3SykYlABdaMcetcBvtTBAloTN6Wq9qw8XJZ27tUV
WLPZ3N29aCk8+nslai/eNm0C7xn93X2OfVFVaTB+trImNy7R1Rc+dB9VJI7wFeQB
NRIaGJ5KucKANLj27iBBOy9sptaugoG3JnIp2U8yUO92oVSP2Y1qM49pdR2sbTs8
mcQONG/a8c1NJv+f4M72amHHp9lu1jD6hgBFVTBv2ibr8EB0Err01IonKWOViq9t
WMsK5XJBRBSAMn9fqlzlIRm09zBRw12wP536tTKwYn5nnm5WiWOS0jmssPDOedQL
yMBaBJt00HdLexjp6IZQ4sNGCacD1BBlyUTYPIJN1kBLTOmrqb3V+En6KvdvX2zj
o/eQkV5kLF/93MOib7/wti9E8NE46LS/OKarfshsQx6hc5iEIDrUkPpf8+cjuRU0
hK211WlcFlGM/Lp0xtQFCX4hKbbdK97T1nE1oBLQ/Ch6YT9ww8OIWMQ7WOZqWUgp
9i+nTj22qodwmvSjFJiHrxX87HzbBxnqF7rKpYpybMH05GGQHFDrfiEsFiptbDh8
RsR61LQcqN4tT2AfrVl8kR5hEs4ucRg5ffrxqMvR5YiHtPUFh1ny9DRpB7OG/caY
ZHzCLSc5HETwcWKNZy2AjW3Dyqq0EuqnCCxijDFHOx5F3QPvdAxDye1s5Ct5Mr7e
Vkn5jeZxnNiCdSk3oZUgUWktcQ5jWOQKfZMUN14+CJp+YuZcL7n07TvjKMAGRwDw
G9EiNajvPDbW+OTYILUPB1Pi6L6WKfu/l2V5/WHa/upMAhP3Fc2ePUYmcwJ+UVGw
UxWzwq7r2G/2NaEBSlPpVrBMCYgWKsdWjO6oAWehn4c/4CEHbtNzl0tIBAVuby43
yZyQEQ9aZbIuMmQyLmn4uY1URdxCXR7ELvZFMlcGTY6ykHcYfDfLSCj1Ogoa5peh
ftvNyfUUBEReLbLhIlzvZp9zV5BQ+6TebDISx54VRPuZac/Iz3hMZzlI8wjs9rcZ
7JmQjycXCpNaFNPWe9ekuShPWohffJWeO79MtS58/Xa+neVE9+x3rCwewHUtA5Yc
K/Nd8wYyczZz741EZ56ZookrjkzQ11hRACFeirbJfWr6QQcN22wOKpTMslYetWWc
MKqvSHD4vyE9fIUPB7WPzzQcN5B5QwD1ovl42z1jIBF43G23kKteH5bV9BTFfvCl
+lrVTvuKvcDd0mtoJKRQ7FGTdoOxl/zmavYp09hcHlQBjuJlreNqhcLt7ybhfbLw
R4AhFWGkXTYaWZK7nfAw6b3I+a427+aecOyWHii2a8y+mbMOMcQdTLpl9pMyhtUv
hSfjdMBtTI1hsZd8W9Aitnbk+hS8jiphdSIIl0Pl1kIbbvdDBvPfce2030W5D53r
tOH8UgNHm3oYILAl9mSvD7Uvqu1lcmjdJkJK4g6DIOOfKb/fGeCIIJT/mOtKcgxD
fakIv2m2FDWZMDIpgRfAG8Kjjq53p+PcQrcvKNawtQlSiseEhup1EMPGnP01+MFx
XLHgnsq2r5rKi3SA+xRiLx5BXcKWbpE7yjCjAv4Ai5t0E1xGAA7rc8J9pSF5CGKu
HpPf2Ch2jXSTrZZNkvNRCc/Ede481DGguN4lV8MELwXae5m1xmN12iypq1K7Y6wB
fb7Zsa7Gi/UcUhl0EEptzFCHPdVCpEkN3oueCwPJh2PFC2cLyn+oOy9ZnqnDT+ml
PwQhY8vzPa9S7+TnATm5suuiLwM3T2yxnjvxxqAQ8cSiar1okal+BnN9YQTJ47c5
MNLfXe12wUql0oSlcQmJ1iJfNXL0TDZOsBTbwU0oUPjrAUsZdXB9p9Vm3enmJsyO
swJrZotN1wpTXgkqiP6o+C1XlRGFY0LKOuXAINOBryTkCKvxj6Ge7lUKN0XKEzPO
vusbL4OGId9HFj4zuYX1yXABgBnXGm3WwBgAq5IYg/9SKqJ/5tYqy91IRv3YLSce
Z6mH8fNWVqR/7Z/gOZ3lZlVv2ri4MTX5/CIF45dxkLKHT7qieyluqzYUTehSB9sC
Rv1njvL1nEHH/1dWQ9KLFMd/83dFuatv3nODrBGWOEvi9LRfBUYWerOtJstMz7qA
j7K0ZiBJJFeYQU8mJTc/aMEqEVP9cxz2G8yZ1hEc1dd0hSCdFfqKXqu9vrFMSvRI
jVtyeD7uPqnytCPJLTPVXY4Lg6FI8MYGpQO/ePN45w1eCerNpitxH53I62OxmXn0
+Fay7riylw9CPUuwnz4EOv9I3YSA87+Impij7j4vUq2j0JYe+/IX7R0arX/4rpG7
VJbzeeCaJc7e7teRDdN6vYMZKr1hqRffc6s+zuCLR2itrvOjy0wpEeN4cULk52iz
x4fFX248/+jo7wBCRzhQI2wGdX4pN94mPln5qneYchqIRlfx4WJQcbf0gW6caLkw
K3hOwUn7Bk0yfm3ZT4/QGZTxQ4e8QK93D5g8Nh6gzXNqjSsyRAkJaulV+WILmTLH
UbzW7P7PPeGWGalPzzVyvW4PhWY9GE9wiOY3zE8LMQHOGEfTCHlnJhSmuQodLULt
b9r3V69FkR4oNAxqCAfQmoz3a/8nUSthL3KQLK7RhL3fZ027WjsWrSUFq+yk6Mbw
9wnlOEV04SjEe3qkeuuFYH2plgG0gmW4OC/xynRZfethooBcYwM1BlBZMNPhuR29
c+uZeBH2fRBtbPKYorTqAbYbS1C6hua9KRZM563nt8s9udfPGSHSR5Occ/c03yQg
+A/c+dLYw67j3pyOTR9fU5xjU8kdouFDAheHZyhuvjfk1lOSloxFS/auMDx0jVU4
2fBWEAyf97tTPCPTR5Dp4rIPp7xOzD9Acgv+2LJOPshYouUeLZZY4fkTCvgZWroZ
x1vstknBVfeJOPFRi4ApobhqdHqxYNgDBw5uK0r2G6JVQLiwN8Jmaenkf01OESZ4
L7wexBq7c3jzwYpIofwSkW9OAMo+iwVA88qZkpkxsHApjH08K6wK5U1MBs/TDavw
do/uo0B7JLGlYx6Xi7IVOwO5OAQHDPy6DKKkBjnjX4xyzgydDIwt37XlOwZNMMvR
UmJRDVvJyHvJ3iE3rd+xpizVamHyXPY/NjB8m5RVz+VWE8uuamBZIm+59NobJri8
baLxKnuXrNUhVVfycPlg7gEXoQK87b142Q774fVOWm6kZ81JG3jNift1itLx8CTp
G9/6lBJsjT6D6jr19uNGu9IMqQWHnjAYqJe3I5YUOarzMuo5akoetj+kIC8onyUR
4ArLUJ2bUZ3SwBTXAWPEe+OznbGwqoLLvt33ow8GDsw4YVyQ4w895y8s/vAr7yhS
xQAgFzHr9pzSGKqIFJQn1n0QxmcwgU6Gqook5rAAZddY6AUaLf2bZ94PTkZaBt/h
fFWEYsiEtlx4RXkvqLer5oPvWWynYAMGH3Onwri/PDzEUDWp8n6rl7y1k1BelodD
7YciOPvlMvu7iD560TnCh77A2p8evjoq+2HP0SjxEXZCo2KaJIif0pj4eemTrDCp
m3ai4lep4NxZ9ZGrMZmOrz4ug9kJMZjAUWyWsjycWBft2ze7hmLclI44h5b2ljnM
yA7etYk9CmWv3SFv6yDSA6Rl9fgFK9VXRkwXbTV12BOilwgMRMrj5XZAWSeMumA2
SVbO56MMdJa1vPHYCPxskbY58aRqW67MFRGYvVgRGc6+D2QAFVp7EGF7GMoBuR/5
tUlLyf64Nhpr6FJzdDA5eH3JWrVeIRKilIc+qwfZmIghbM9vrXdmfjbiqWu1VTPn
OaFxK8me9/VKZK95+nJAt0gxIBqxkWbWlj9A0NQYdpcsU9L+06VKgHtgRFqdfnb7
nRX0z7BOp+qhxOKLjKu51qOPfNn/O43WXofiveJq/6byBvH6gU57gFoN1AHiXv94
dU6uKXvLoJb8RMqeuFdlOrqJZD72W9NWR6x9qzLmIJbB24nlbxglqRBsxQUdH7SA
uQxKseObssmUAtkj7Mu+5htsKzV1qp6zlTudsOZZwtv01nGlr1xDJTcrD4mSnvlh
jpOiKVjQNERKhPLd2qpOY4hpw9MLKNHjC+h23sqyNVHlA26F6dc9POKTlZ0oIoXb
nBy+69so1GybYTZ85l3B9wj1iM0xSC2juXpvlVb9kMXRHz2WSU03SBDNVujJw0n3
Vd1xODuaZo1raY/7UqUtRc3hLRPWUPx+pbTmTpvqbABWJ3ZOvCOB+jR/PnroV3cN
0nmZ5Cg9xL9OGnDyHSUa0zFFfE+jsBpgYcvtd+X0ts2ZOuFoYnAr7KLuOMsV2CmF
+LorSUYd7BvfnBzeN5fNenBLFmqyLWaBYPK04dTPi36mkkWfBTXHRuwWS4o5tK0W
pUEU6U2V83lqv5dbxlr/ugpLnGpPA26J3JBIXGchLhwWIQtvQ4anvPUQTGOJR0Xh
aye7/NMTmSt40aCWiE7ahZ5zTVuYMGxTZca7gDHCvsxb8mG4XXvfrEIfBCBJocOG
LJZQTMvPZosK3bsd6zA8xDvOwLwghtcyBysfa+f17TzFxsasdEwdA5n0ENCOHsTW
cNwcvp2rGzqycy0PvZ+cDy/IPU6m5MGWJfGGvuahXsKDvL8nWpkPbK3cDgVcrRQg
n1iTT3mMRL7iu1icjYd+DOfAcbXI7pM4UXlVwkmCSM+FcMN44Ubm5K5qchc77EGa
ABA649i9NnFRJh7qCu4bXuGhsbr4vYOaoKpLYoTzBA7SOo86ANsn9WlrL+Gr8Cai
8M6O2hiE23dLCqwL+y5BtqFm0whMN18z+z0dERT/BiPcePnD8C4/x+COiwu2MVE6
iopH6cMILbBpbjNeQTOwSEmXYhCiLriXwqV+GOh9VlMnfymQC+AhY0BcrThjdNWE
xtPOZmzivk+HgXNwzS2yIROpY3onWtJKGFPNX8Krvf294DXkFdvQ2HEzgVaAslxU
ZnaTygFykNsvDhcyBfvuXGZxe54P4Szho0AJAuNv9DhwGjLsZ4NH9IjchtwABims
nezSqIipoQfX5Rv39iy9zpsKoq4WkuwUVo69NK4S2hydfpylERciQJSxl4+B1so8
fLjkvLQigNlkhn3fPSFtUqwHmlupXklOlOtVI+1F6VrCOdDTNRpuYyQiyVyRzLqY
W95XKYDbnD7AleJMrGXJw9mX8ErvTArUNYE762cBQ4PTaS3xRBBSyN9+uBbqg0QT
nI/XDtMvm+iaIyCYTjN1JICUwFcAYboH9n1cMURsfUcZdhZNWhT67kXuSajy3jVn
e17uzCDY86SoGd5YNTURhDQso6KWa74N3L3c0Tpa/9l7SpW33PqfTm1xOF3N2l3g
eizBzAIRUexwQtVFuKWza2CHPrnX2weKs4UVKtacqhu3ERPoEUR4Xch2bVgAI1Ns
8WDP7+h5FIl5oisTPaq1KhH9514ywGeANx/usAJWTaOhWFhqp0DXNQztSCwAwXCQ
Tf9r/p7hkhQ3PDpeDIgyqwq8HSs+bqJNcTpI/l34oND0zrcI5K9RKV0BiA7IXFLy
sANgwIIAYogYvDlCHdfULOYOFwYO3gi7c0BMEonpMVxn8/aqpw5r9XuPEZkNuAPL
t5h34YkzDyU81Ds54JpzjrGMdehOL9E4XTDmqWBEtiLpS0intrF4y+bHKQmZoKzj
TNAyy/B09rWnZKm7xr9/4zaWfbycQqzZZHN/oWD/bW3kO2YCkV+vz1lPXtjVxraV
fzVnpLRym8Z9Zp3FBPpbgStbTFtAk4fmHsOrTp8xhoP29gGMarxlWIA0X9HOqWt5
2loADk14qugQI+s888JwcX7SJETHlW+X5HqFBYPG3zoldXCsARfS5oiCQro8+JjG
bFuHlH2ZRpNLmSUKcFj2PnZVqunnXklKun1rLAI7PPE2CQjLaeOlRy25dtGhgIbq
QzkaZfrfJ5ZsVVcbZlRTrcFqJfsR6TwqwbemNp1n07O9ougn9V8V7cm8opACjuDu
StqQz3dpnQe4sifQIsorY96bGBZykeir+dAXrcDHZKXnApiMN8ao4X4mdahKexdD
IuYg/qk8ZHZ59Idf9j6JYgWS8yRGu2qpf74wzqOYeVPvrgDdwZUHcY/3+p77dw7q
LhA3s49cT5eczYbBd+0XNnLGVOhvWhAgCoH1je7tvZMPy/exX8XFo3ip9i8TUDXu
iaTbBisFDLJ2hsEujyyz+NmVA+doUWHJWhPlO77t46ScR1p1h/+XuOzSeqzWYBjv
TuOi7gLR2aDSMHfB6LlVO/G31G9d4CAaXsRxs858xSvyPsL9en/wYX6OV+vLIm+l
7EjtvkkKHd+knWtZM0jlVu9KZzYHv8k7jkZZvOUeEvsmFhpo8es6ile8ywjptmws
gvUmPIMoxDNQ8ey/OYNqtVJnaLeSvJVJj1u3zRl8/kaBNFWJ9yFf+yPEYn3F2y7F
tn3L6DRmeq01qFc72xhJAAXd4XlQiFA49KZ7OBPd34ftYITuwIpIoBoVQDQWRjpz
AF4SjcQFaKbImqraEk5O083zeG02bfAYhl7LC4zIzLfYgIjeufF1nEnMaQgeDXRF
n5OxoVI2eG3MlFybiwmpmyNWlDlXrZqt7Q+Id5nq+xBuWmaNxzmCkX5N7WLSl618
bH0UU3QpCkfztUS8d98O5G/Kj81kk9LPsqOQeYyAI8nldqwpUqdwlRFJxHvwWeRg
p3v5JjpUEHGJPIbWo+125pQTx0lKKZRTH08/SI2taUEEqOAd7fWiqEXnve9gQ/Xn
22qK4TUPeorQitgoxqucD5ua2A2jPv7cvQGysYfyLU4FSRQsBSr8dqBcFJaoJ6h7
8UPicbzajlLfs8kgVoUjhpEaossjLheLjGO6CKfcUEM0i7wXxKZXOn+CaJ/l30k/
Qm1bvPAV3QK3H7B8u6sXluBaWqr4ckuW/bCxNewG56KEYgB6QxRpd7IublHal9zO
mBo3+CMu3tF8K7TklW0XXIP4GDKEX8eUzVJ39aamNF18uDEkRVv5zFNb7EQWCJmm
pU3Y7C80PH8OcUpYyfV7NT8eH4OxPUlXRylkS4AlORnRpI0LEdV7GKm4xJG9opVk
YfEyUOkN9VhX03qGo9Y79uqFb0Qt/8T3zrFAr86fPd/etaX/8rNqoFBIJvz5itmJ
6MFIp/S0jSIy/epc04pIZqeGBTt/ACyVi9fcZV3iC8gP/enLxSWal3b4I48qAOj0
XstXaAEt3zSqbKEdxeTE7rHu4M2dwRGrOAOdukERaLXMsqK7Bb3MvDsMAYw8Ez3x
bUlLo2hEcCcO/j2hcY1SUm0a9vi8hBALbnI+zXooH4d6FTrI9oRvCtwuayK4bRVa
3EdKNCvk+L8k0zgIylVNNpg1US1HmN/TgWz2Y/KBzEJuP2F1CUOSNyFyAxEzHJ9x
DJlRqPadrdoiYpQaWm0f3EoRPxXWJ3bmndgk/7A11GZkz9qwi2zdbZ1suaqXbIC4
6tedvDiv2A570467tAxUeARZoEE2J1aMwSma4NIzVEFWiMPnKQb+0EkudnA3hNEv
QBbuuVBI3vJ9Xz9XiNF8cK897rWYOuUJD9voq0bmDPl2DjfiUjk5GT+tgF92JCJA
VCx7Lrj2rCbA1VezBkEJb9WKpkCFxIJzHEI603SceO59BrAdsmm7RYnNGwUHPEEe
MLcprKhxbfvUAJopT+abUj5fF2lJQ1BLmVNUqid64yXY4lDUKrD5a+H+jE7XTYPL
C/eeL/BuOEtC1B4GXQ0yanV2gfWhHyT/LX7ny4kSnk5wzrT3L9BH6EGyRoq3c9MG
p6OpCuxBLHEAP3m7FTUsecUgJv2FR5BbpP/qXMmpa2+g0/p1qkgtTNst37RrHT39
hIvRsHUfPtfy4j8hkhVeIebt8sdxaAQ92vq1hnPDX9H51JD3CMBH+yTEsphaNJJb
pvopSKV36t78U2z7qTUZRe7tYB5+DnENsbcPLjkFYatINRgJdGAvfwQTPU+D9tkx
L17DcFjFFg3suMosSneB3xOGzKJKQcyWS5wYBdV+wxVPcOFyfJ29+kYBEIFbuXzx
J93SULd3KD5ax/LJow8o2pUO6bRuBmiRoUxc8g6h9iKspukk5py8S5Hytqq0orhO
IHTxqZxFDxJDXoMdObNOl0epwfinMDhX3AELYmctwYh3pv3HOHZXN7EnUOxwIQEe
+JGXF+mj+BVdzaoF9wumDz9muu21lMOsUmOdtR4pJTOM+Hubcc44cSLE2pE6lEfd
3wUxgPUNyntMdufXJVxh2pnIQ112a8cTG4P8L8Aag2SaCuPRp8FGKSbDCKhWl38e
xfg12acMw3EPAPf1WCbIC4yGYKz4KV4kpHNn8ADZXICQaLImC23IXJ3P58Mjrf7t
B/CxSl4jGo+7HKI3S7CGN9KXUHJVdAzXbnVvI330oiJI4fCEQqS5sbcvYmFI4GkM
9/D5JHuG9JU0Mtvo1bWyshzLbxqcmZi2bg6u+yvUQtqwZptm9pN1KAN9PLiFI6Mz
I0lhqmmLczTPxcPwvS4fStTKX3HbJS+Bs69dl9qKYR5nc38WOpxFMC3Om9QJg3UC
1H01Bdvgh6KpIAsImoey9LC3MkoAykxk4IHemgzYbj875akrzR4GzantZD6zGbH4
s8Q4TnRxJ2c/CnWoeSLBekM6iLedGKrI3QxHj1wbHcsMcm0ki07EraHlEFCuvwym
UDZEm2RQDeuNfpFD+9RzCQBCxUWkC/iOFdT8gKGWI3aVh2Ry9l/OW+3GdcVRbSA+
VBGNqH+fOD/wfb61K80/7rHtNVtkuFg5kTcr7LbcU4dlZDR1P5taf+Vf+aRT7baI
Fjs5sIn4tPBptLlnyUaxQXXRR9f4HU0r4P4xmTXSndklXbSQ2aTIUWYV4DDLiT/3
KKk7nHLQOKXv6dKApiD7cG2Y+SQyUbQo8WRY+pXnACETSenroBGikkX7hu4NyfLg
rT6x6INnPlQhhjBLEe0476Vv4y28hwn8GEmUVrd4TM56q83PSJkBhz2x4NfGUXKy
HDEaqO5KgAAH5ce+SsB2SbjISO0RQygnqMwPQM+1UMPzVmAxfsB75XKF2ueZBlBH
thgMG0bXKzVwyb29lXd2UX4YddNQ9K+Po7YWnTnGDFmBhPb7Scrrt9/HSVT/ssG1
RkzLTaC+8W5mWV2Q2QYHPXRk5WFqJHLYxHuAZpS/XW7ZI0qKbeA6xj/JGWB7teKf
W8AcQwYiDgqtVdsnzKY7GA5/NgIpJj6KSdK3cfygyGoJbANTMzNDZAz6Gh0IfhsX
lQpKKYZsnyg7MnirLx7+i8Wmn6aaXPDD0m5CoSanE6mIQ+NRyv0WIb8hW6/u3e19
J6Kee3vYPg+8SdM6go/5E5LliTBK3WJo0CUBxKlC1ipu4P20SLNk1keZiLrhFBXQ
Ae20vxdR26d4qEfk8fAjclls3thgIxxMGhHIY1lSqeXZZmyutGl+vCP9c0gBY4ny
zpgABKZ1YahUD/t4HpwrQ/br4AL3S2JKiiEcxbNFwFQ2M47aTBUdDB3ak9vtHSzl
gNKuAO2XTIH+Ciq4bZGcZjCBtiNg4duRtUZtKoUPmpC299MTQq98hAN5yv6GVrZy
j33TNUJCESvgnhaSIslzNApzxwBmcn6GxJdquJWJvxiur0ednWrqqxuVzhh8qY2M
8lLy0iiDoqUA9BcHGBgzCoMT68VLNQICWmtJaD8u/ptEeq/5gMDsgcxFDAxTkzfB
sP4Hv8oz+aFAtz6XNiosDRpp6xM8KuyRw+UaJ5hY4w8a2Gx3b0GqXM4zKDl++nfq
PgRxYKf2bmprbOjXErHmGkJ1EDn8s5QhGQsBN2D53PUjrgapewcI91FCxVwrMK0K
VByH6LLpoSve7j/wRDZU/4MqwxFwl3VZaRr8S/4MBMsuaLas+sQj4rkeSPztY5Jj
D4+WXS1t0oePLnLGbs97jPTRKkQgTyLYCDLp4soBHteOX4ozqWubncmCelW0iUGd
h/O0kUNm8uXWkQ13Nh99C01Ql/QMU4voWTTf4O2E28P0OsTWxZ6gvSpF0/xDgD/U
+pVQoyLd4atJaEVJ52HlNNBIrTx9YMLQN1sKRaUzwwEGn3XGbdbhubrRfwfGgjjQ
WPTitJNjNYlyQvNoPboVVpxYx6yyQ/+TmilSEoK1sVJ7VWjDNjFHl3BdHX5ibv2j
hrqlIbJmtPsSzOv3lrM0WaoD719VxNHTL++eqnsiawe/3QisRVbRhxk5q0TRnG5x
t3j6j2gJV8vEqHy8auzrqqSEpBu6ht4ecGPbi/i//L8a6Hygp3RWhewb5/HcFCEz
hke8/sgB98dLWOuSExoRSOe4R1egqrMkPa5YH+DvahtgcP9BzQNfdD0Uyeh/JLOa
/2c6tT7p/l4RTUYONY1YH+3IBsCQHILjThHqcJCx33jEg545V5nvp2XEgBU4MHKn
xDKa4OlQzggHbSSoK4Eq4TElQXLgBZrWP4mcjA40r9BzbSeFLvUXjYYEYKGjABI/
I5iyfr9wpwTTpTM65+eXpiDhhwMcie+7FpsWjtfyYY/G3FpF/ZC+1A0vSOSaFY4d
aWR9x4gvG/x5yrqyOqpxIzspnpJLwaOHJMljXNi2nu6IILdWWPq52RONoWrz7wdW
F3MyxxBuE7IjOk0WUxb38mmtMcQ7xGx3j3+mVR7voSQoIpNAByhAV47x85MKEZ78
YlmnmsuzqjRjT7EW8XOYQCr3GfwJG75im65mumOFWFbJmloqUyVDEqrwaIjMhXyg
7IrUucvOw2jI9G/Idv93tURs6v3gMhVsjriG3jj65m/cRB8fKQ41GanQ0Tn5/pfN
IcI9be/h9PI9iHCfqIT+vWQnE7JlToHNU6E6K3G+aMkC8rIuKbWqK33lBGTQxKgK
roqwxTrQDlLsNFz8PUpJZfLtAQwxZmgNXVgT5W0cQmQa0E5tw6V+W0D65AzJW/lH
DEocri8icP51e0ZP+dRBGI4ahanqDKlfPzGh0ydQaMHvxk0iZbkrq+GBfNA3tIVT
QYdz19SVe5hqT4zJi06/MNJZ00mH9psZT5aW5zL3/jlns4FyMh49HpYaaKYJsz8a
oCp/RblDKMsHN4d4yOsYHALCrdRbEj94cTYq5p8bOjgP1Y5iI/sYWXsVGPdbdiK4
rd6gIxdqxruXENuOcba23O53y2ShurDMrbr4j++ONKC2TgaKNHu41CruZg9kW2FI
H7NkJM/56djMqOXemYkc4wsoVIsyOEMnzwVIo5n7UhESL06u86zWby+Y4NOP1yPT
z3VUi2IU3TW2EmlgTPZZha2bmqjE9rI1jisAaS3fwgmsyoeuXqO5EE9FZdMSjF4m
rydewsxJtaJg3swbFDiN3gZiMcIMm0OH8eOArO3BMcGqD31np7e0LlQNjiWd6BCB
FzQHBK8a2CwcrEiQm1f7Mwc2+1rsCNVD8XkVG2i/5oZA+xVwguTvpF4F4miZV4DW
xsTMauy2HaxosqgSvj1DZfD9Qowez/lnmr1w2YMZP+pOeanlID0jljKXEzBILfMJ
Wln6KqgfRjTjQQfAIdLk+JO0XaOVfXMPXzFinhqhc0NZfO5TBE2uXMfKLFW82cir
MTtPPq1xeaccpc6zrTfCe6wZWXYMrV0YoalX07MVvJdDVkhjdN+2lU5a2PuMcJUV
Zvc0C3QduHqX3ypbuqHikV+ERZCdy+9oiALSiKiJRwtsvrZcWnu4JbapjmOXG1Oy
k2oEr6h1W9rxQTEBd/llV3p7M43j500UTzNWfAX10gFphvY3YSmTfNNTHQvFOs98
3xC201O5GTnkvVyvVV87ayJy1BwPRsiUK8aryxteFpGXd4m4MHctKgzleDxB/tUJ
rPZT7bpkySUUQgj0SDUlhrcBvgWsi11u2kZNQETQ3ukNKJfZHX1zgno0RTYgqziB
Wtzw564qWgb86kdCFX5JLS/SxlhoN8ftUJAoDxWAwmgdvk9r9SPDrUTwf/UbRreK
ltLGflAFqaX6Szr8eQD6KyqTfFQ0s2ofDJOWnBQ3gHgSOqpCVb10oC4jwYXZPDNe
MNG8CNO68kkLj3pU5pmwSPuCWrEWX8g4W09Y6Qge2UF5pjkrHaf/xOyE/l+VvwKL
g5VRQCbLVx8gK2mVZ39oQ/Q5a4pDHdgAsGNeNYSXylUGbpAMGDFuR5VAo+CcWTBg
rrF8173N6SOPaGbE/LI9Wbt90rA+/DtadpZrDPIAsiizuZtpnzTmO32uEEuWpQon
LDyR3k+BblK5eCw9224OZ/G+U4ieGknFpeim2IpGIFm3rXlbHAJY4xwGPWUZWTMI
8zi/HR9bUWuuxVGGcuV0GAQudFOnI+j5Xogd5X/ELa67Zq6B0Wc/FRfcKoi+a3QV
s3H6C5R7UyRpPGb1EKCnACW8kAA+v1BmWN3ugQTMEFHxv1mphN0xz4Qkj5fPk6mE
U3aC0ddWssvLN4KEJcP/o/Iw4EJKntBq6I36MmgXvldkfJXVbTRW+nC7RHlH6MER
M6+RHmSBmZM2Mr68WTVVCZbqmCqrpXIqS1Z7+hjJP6K8AOVuHDcnzV1F92D2+XAy
9YKDYfDNrzsxB2vRttmFJHYHsYDsynjeRIqE+gmmEybUUBsyKEQMbzvrL1Qvr6Ex
zFmECB9QOEKZ1O1IoI5r0jgH3nnoSVIwRbGrO3aKxzUxaQBuQIS7ZRcOH01qyx6W
7yAAuSj5ud8p7f035kfhfiqgeZ/cRYPC2VpkJ7bhZTGP7GZ8KakC32dFNkeIAfYa
W7dbRViirLpjosUqOrl5mYVxaIZvsfDqrgUrzf+zkoJDpkK8Aq1JOwLmtlkpJaDP
0IkrQRBQP6Warkq5fALrIDNmArlGrzVN8PU4ltE3o72pkyPGEYef6+uXOmXz6Vin
oL1oEjs/1piCbc/1UW/V7ZLOsHDHQQPO1gHqGxFVWHB7OQl+K28Af6X7p5ZhUvJ6
sgdSVcTpXKCqNnM8Eweaos/0PEGYxA4NUAYa4luSdMs6hQUwgxuCOYA6y943p5R5
mbpZicyg75NLedlNwTlMHY2Coqt5rhm+VXI/pD8QMz4lQ5bM5zlOHevFMxOopoaD
dKy3qZeUpXtW7CMqyPa0F0nrlG6b0J9HP3VeTRWVIgbTeYz5xDzSs2evanvdkXpT
ws8R0iSOqDyY6QoGb+yTR/hmVoY6FbV/+y11lqFWgoonBzSL9EL1sTE9hJHEsB/V
0pATmAJZSgtXLIAAnCoPTXTBPeJrpnvjeLqjm6RACcrrxWbnQbw2CWBLbuEymtLv
+GaFrrRYBpSBA9ypsSOwBNk2+BjB2bAyjhb1u+fq1/xPOvqU0HPtrqqlxDNdRoRa
8m5oZcmHUcnAZv8Gz2DmY6ZIuzKbHpCxeWN7d6EYKSWXLXJLpq4aRiAX1xy8geyf
e9o9FxbssApIkVPrOSMORY4MpXbFayibKCWa3hOWgBOl6QSQvO5cDYZHTNBRMEpK
Yyjzv7LYKrqC3Tp/zz/25eSS9kgB3qKenEu/R+56Lc3onezKFtMc65LIQibPDacV
D0VeWGmNJSWuyDiW3MkOeDGkURVsF+aNsvxUiGVQj1RaVfErTIEg4Kx9hfM66DyS
SM1zlVlLaCPOe79LciMsYgxfaNSKkAUnnCJWRCoutL21cGUsEuLPIqAhTt+5fWbh
P67D5Xd6MNZVyLJiiyXEyclBKpylF84MrDAAOvly8orKhlE7ah6n+lsGP4KAb8Ci
NWwZr3Evnd4lsC94LkY+nLTlKyKxKbFDFio4vnBQGikJ56LSwcF9VSlSFGoXU0Lt
C+FAZiRTj+uBxr0mpCboolTm/y7QiBt19NRciXU14EuSze2OqEK0d5SW7YmNPDJ/
iSAGL8bGXUwjya/TdrhSmt3LJRoiIIlL+Njps9BGiamUh9vPUneZFRZiI/gEark0
mqKokm1uGXaEdptzXLywYgHcdqx58hzbL5Dr92O7ePyvtvdCk9qFF++E5/Zha750
b/wdHvp09CQiSO4XvTGpG7kjdDZtedpGuG0u+3dTjXphVg2+ugakM2nbAAT0XB0H
gGPta0//gELefYmeFL2BzaB4z7RXbF7ZMY87PHm3I1NNii4aValA/fQWicNxJl1Z
pnZSblzii8sUptJHgGYNnUuEO7IvRJE8bjo1Gy26PuCoNpF+F3upXFhPMljBHdE+
Jfs32/BQ1/2TYcVY7xyr/577A5NqH9V054a+DizKCGmzL/tnOkuBHza227GzmpT7
h3Gg4j3kadbkYiYlbbzAh4G8wyzZE+4qLkMye4JJ8aXq7r2KKPxuABnq47mFtMWk
IvWOFLbwlkLh4dxMMgWwW4+cEWPlWLHifglGa8BSOf1FArJBLdhShJANrZFJ+hWa
KbAKemOegg2K3JDc1QltFuVCwdka1MwfQpbR9rsUe0ucugfhQwWT7p0spBuxdxoD
GEogqxBchPyzFW1/l12a5OdPCoNXrHcQ1AF3fnk5cxmfqqZpn10f7bShRwVCs1We
yEoBKyNPuF7cDhJZQUZ4HAcPRE7V1vs8RgjPaUq9cUCjopttBsVvSeaHlvKgqYGQ
pDzpfuSSUaOGOwJo8xdTU9hiOjJakgTlcxEZFT0YWU/VOGcFe4z7PXczh8c+dnhd
IEZyHpX+hJr2IrhJaG8hq9jI6WlAyO5e3D+YXiIlh/R4ABIWhheExsJnH/bLWQLN
alvAg0+IPvP2FgzUAXkF3c7qT7g5t8g8QWvgj6nJKJ9NCDzSJRmEJfigTQioHEw/
TQBn0SX6WcunbwuqQ1JhMMHGdJLmGc+jyDv57T0kR6CiPEQfWvQzMQFtmnfQzGhK
NMCy7ill0mLF2NXOsQqj+tobwWMhS990WMGrwdxLlffYRv/Ju8xnBCA40Qr7+lfd
KsOpunRyBJw8gO959D4tvEKFLYq1PysGmxbbD5qsajETpioIfZcDAqCOG9YeLOG3
YkFigi6ylxHvFEvmxli6ZejP6hXocfXG2x1LD7IfjlSAeOAgzx/to1xQnGaW3quB
3A1kklt3n0ctaUxQhc9LfkqHVxtgqxLLqexAB5MghzJkui6zp1ve6BiNS9ojtEPs
fjM8Klfg8z9dL5AvKJxiioRs9Hd39fJ3t+Fprs73Bl5pJsQOQ3r8S5Y1htYEY6Im
0aMrSKlKJ5JdEm+XXULbqQo+jAHTz7+4cln+5NDrl6LTLLhbDK1yU8Nh7FOR0Y3Z
KqTv/+gniKaA2GPEIq+Nosi2CuedFiCDeBtDfYXJJNVUzsCqEzsbmctsKCR8zBPo
00TT3UPUXp7M02BC4wgymDoyr9XaPYNmEkx2BKuAYRakhNu41JFriO7HqG0QtKEQ
Hc+63vfUrgwrQSFpFdvMAymS2H1QIkarbky8PcEC/mZTlNeb1arZ7MGUuVpWIzf6
wn7kuiTY/Z5IpMKXXDcRosF7wKN8jd3mxaTZTiJ9jYDsX95DuWAT6PwTdAL6Dila
Dr1K8wp1TEO8eTiBpjlnXiGf7z7xnRtmC2lNIXJXod561bV2JCpWJsIGtEpcCVI3
gqNDZ2iekQ8fOcjrWpNgqphB5VFTzLCgzmdkIRsQkLEUaZttTidy6DbE9cjqu55k
2XYuHmiiB95E+rEWcL5fZqV74GtmRbCDWtJFc35ggo7kApEGZMAqZVXJuwe8Q7uk
Dy6fXXJKCmFRHo++9IxuJpI0E0XNEJazKDlVdDpebcWxtodYbQwNnztCstf+c9PN
m7JMx1wypKu6POuPX4OnQibKE59aydLMcWutpMBXNhL91UW1eAU2JrySZRKIPLE+
IWBfL74YvlfSm3UMikNcXHRVby3h5EOiOMDP33+2p8rg/1AFWjLS2qAmnC1+pH61
jCQv9sTij6h07xL0aQFEniOVPgUxO+0UwqzkK4XYr/5/ZU02jf0oAlRV4JMdyt4p
8JxQhBjtpvv30DuHzqmZLNcn9pZLHF7ARKevPIzW4hcLzoqVD7xzk+c2KTpRnYMc
kjZVExAxJe4yGygNtUBtMYYhbdwu+b6b3BFZBD+1S4lgcBotDPKMMtPh+aBXqK/U
L/FPkfq/M+xOOfRYNWQ1U1eoNTrJsznS4ZOZKsFDYCZuxpB0D1k1Vf4GnGQT64V4
euWWvXf2mERRHiVBhR5Wg5I3oa/wbpQgIyrSxytZCYac477kP7QR6ryhbXOrVfR2
Wr2Pijnvecpaki0ofig3Ez7IkqcF8NTAM6tV5GWrR4iOZAJNVhIXBNxhEvv/RB8n
MPsbw0qLLJsw7cxK5FreVJiBWDgbMbAPrN5qblhfOLq68/zyETVDM1PO5SSWRu8y
pMcHi3Z8Aj9Gva14vXpb+ur42MSrGLeJaHMVXBtNTI6rHAgqo8Iql4gFLabwSELf
lJfAc2pGDnXi4cAE2EEyFDOW80uYHOKEFt5ChRZ4uyJPEyu5BY7BJN4zQlnJfGoD
ECIBPj/1jRyAr8Y99y2XANBmuGRhn/hAcd5IVS6a2J15JU/6Eu2NVdPgavQ2me7T
W2qQjGabMZcFZpJQoHqeICn0vpky538qoRt9um0JaMrf4BJ8AYZ0wa4E42kVrPqQ
jeO6u+hWsjyGLGW8t04t4cWlk2V8IRO+N8XcLtAk2VReh2j4wEFvtKN9rpnKWOOj
tlZQCNYkwAZNbVI14jgiyZixUTaxKasvK23xutphD0GnmOtfoEspfP2G2/BgEj9N
Hwx0ysYj01mv0UB1pGBzn4/JAzdVzMyO3ox+fwF9+0yVrLo8W1UO9qhZR+rstgWf
eesoqKZY1gHefx0zVxRrNHDn4SoxRQD2tmr6gljSgYlVnK5AVhlAFIs1Uyh3IybJ
Ob/v9A+Lw8PRG/Z3ssOT22cAKjTctXwKR8iGWoDPTWUaDTjaqN2ujEo7pioVcuA2
xQoGV+KCl+tP7bSeIeqp7Oyf6czHGI0M1BQWzVFz4m8+NwOqeMFGQ8FGzQmUKtJY
AduIuXGMHf4NbC4mEf+Ca4fnv6flq2FqGGgm/d5myvUfx3B2o3UMKIq7qSm7TLxp
2P77pAbTj/pJc+pNrCZuc5y49bpcrS/cWOpFaJ5Q+UytCo+FwdjV0R18dduvxoRi
1+Kn8lTigiF36DTITQhlnNqdsMNJEO2MHx/bEwwmcefOlD4QOIb166aNG1Y1rlx8
RIb6QD9NqrREcU+k7mfwi5GOkPfdzGbMgWK2+oscKjNK+qJQAJk90J06VUw7ievU
DnZqFWooK72fg6puBoOCUP/iG6sG8Bx4UbZCZTkMnA6CANbWon8l8hr9z7ApE2dh
rWmt5NT3ofQvyg5vbTc8IReFPazoyNSCCHwgG8o7MTwHk7ylh/TUiw+N6fmPsLe8
AWt1WOd8ej9KSFHnfkzOfkinH6U8P/mCnaSt/WydxtxNNHf9gm63d+eBO3ITVHGH
QmMPU2TWIRZBOnFvB/9hMXv5tPpbxHKNfwSC0kSxUyNwdUnNIbRljlZBt14iSnJz
JVKmXlXdYmxapfOA+A1eK8IFrZiYNw+aZb0PC1/Dpo+qXeQreKn9SBJp56lyRU17
vK8jLCDUPovsNhz1sBZwQikGV87fxS+HgqPkU8mMx3eJoQAX5qRGrEgSNMJD3NkP
lMvstnM8jr8ud2ZHuJAvRVOEnnQRDqjAQBKvFoKermnuYZtQzuDw8urxfkdTFda4
C3PxDgzDlLewMMA7frOF0KgYcNdZA5aUA/5VzhPnRJPhubFqJAIIcFo9USgJ6mts
lm4nt2f2Xdd+fVrGHc1znBGL4C5qQXPpFoTxnDqJx8fjSW4FtP7uycdf93Mnt4Yo
TDbXhZ4lfFGKgkYO00RPjgBnlnkK9YQXUTv4E5iFCnujfzzTqLxkaQP5jDhPGszV
os4dY5otUAh7ETj1T1Ydu4wv5tCQKoAeKIRDkYMwgvG0z/56C0MSuGsn8E+Zh940
M27VVkgvNCQQjLN3AnqNB+n+SzHrT+YuFnMobjdxjAxG0AWrZQvUQBbhZ3KeiaAj
xWfnNQMCVL26lKgtDt6QOQrjUP6YkRiZBHJl/mzVp2Ujcgb06Gvt1pcRGGDgCgr+
/Df/UAWTeRabO9izJBFTX8+BzDqkye75WUU4Hy/jtPDUdL8diCQhlijjr05kt1gu
/eXA1J/NEqR6PABcMC1oQibpH4PMI3Xnrvk6ptNOzCY4K0NWEwLI1+hy1kjc5LVF
Bjt8ONwqeHp0WbquVFCm5PvBUjjh+ZDbmoVX5un1TyY28v5NviNvE19RhPq5zaPA
+uOENEDq54DybQLa+p6Vnetkm7/JyvYAgr+t5KF9RG7f7+LSgSMAzBCmPnPxgcZi
vumo9SaVaId1AXeE5H61Z8RAQ0dHJ7m0nW605AkKj1SyOnGbaQKqNAFfMYJm++kZ
6zQVOJucORtxfOdqtIGat1fl2RuwlBe7C25SuBJCJfG/pp3dvbN9b7GA/AvvuCCf
rkw1an0nGghHiluT6Vn+NVOUiu36Jy5VhAXLhznE7J8RSlQfEh49wHfP223+xQKo
rY9Jk5GSj7SmmSXDTCmI2Byrdag8bbkF70H+nFty/bWbaEfBSASmD9D64+XZIfAS
DgY8MsNdSMjgr8wiJ3wRLwaBoaNH9/sOFPhWI18y6b29G3Zs3DihQMd2oR4cFSEa
Ij6+mGX4YM+6WWkKpRRx0zcoXMobDjjE4HFnREEh5wO3n0FLFXQyIkoJBTs6rYWj
jFMI/0CAYhNrLbrnSvmfzlR+onlGZGAP8s5deHfXYNHD2zAPydOXYHKVQCmCG9HF
pShffV2YhwcfOVB60gV4OaknnLT2GGNM6vbN7hBSRuUkTB8i9wbT8HAY6w9Wg8dW
79EQG/DbBHW7Y+u7xM8zNiIavWF1cAtsNqjM/EVndnxLZ0sygVa59jTvdCTgXBic
fY+Ae543sIfwEGWsMTBoICqhxVSZNOCw1oKA+oBW0Phyg6j6iFUmdVA19ZEb7djv
EWcW4yUxTFjJ3txzI9pkh0EqfvgxVCgKklTpRb9GD7Yh/RmKidnOKxYWnA7Qrhpw
UodBorJfdpulabFcDuAznbN0jxRrWQILfEgcWJ6e0HqVU6p70adPeQcCofq46WdP
550Afx6A5chx0onMCdbOzkue1ehUJq5P+lsv2wyxEM7dqMTiG2gyBbQvwZcXdUhB
yNwrDspBHtG0JsWGIRzhNGlh/o35wE4H0dNWVR5lDI0Z5P/1guyIb0bFTmG6TiZw
7Rtfd01K/wAUXEPlhp4AtyO6xm67lPZvS6iv+QcKIfTXwViTgkCyQPiCAbOxjSpa
lwxTpR6XhjMgozz6wzYvtXOckrHs76vBdTNM8WWSHn7Q3wIflpsDSLolE1V6Hr4H
1dbSyKDl+/xiXjeE4NmmnHJf8t95de5ylj5Ta3ZpT/pStvbNvpe90bn9TfcVb+Tu
s3+l5w4RCPyfSVqXYBkJxUBF7G+hO6FtLrZO6zWWPbOtZq74JbLt56BbuQYw/aXi
aIlRC6ZvMM5sU618Ocn+XsCOaVIHkOgQWEXiePTx8V7x8k/ExAi9vozahmaOInAI
s5vPEIbmpeZK5W7AloCYvkxZfXeASZOQ2fkgDjn4gr6ZGeblEVdowd+WxrwHVL3f
kJ2Xsj/fSv0oKBe4DCxctl1eDl2oLveAAJ5PCd7Vy0o3bh3KM2CkAbg2VbKYvUQi
UsH6sALfx5Gn+DTi09olPUeXy1CpuxyUyNKprTzjkNli4YMrLHHgFxO2SjeZ9xDo
/482B0qw1P/nMje72wHMmtixqzKEOKRfEGEwy6oBvf4/d57kv+G8AChTSWNBGDoW
nO8vPTxx4jxI07/XgiMj+lb4Hn8qLhdRAyEoMER0WgjPzbOVoY7zwAPUkcgKVwZf
+xaEvz4Ft6y6Pi0u6UBn5DplY12Mx5PgF4Dr/kJPsfmgFQwuO5irUXGx/9fB7+4h
+414nPugfDfglofop374Wj/4iQaMbsgfVpNx/2KbRr2D5tLhm7WImfqxs5qW9H1L
kOVu/npEbDftyWo6Z2n1ShWEvjHKo2CAPITgUGCctqR8UGDJGraFUV07oVl7uRN3
w0jk7ESUEYTiC78x9bPKcfzHLPpGNT1zMk4WHSXokzgDXvbazpuhqxaNcIVimZ3F
2tB4ke0c3qriyTXg7aF9rOT97PRH8Q9VGyD17uNd9kUQ85ECG4fCA0F9eXLdgXwh
DdOMQ91GeK7RuN0mBRdu3UzW5qflO2/hWiBbLVj1iZJ6GCBRISNB6IB4RZpkYnWQ
4lVTwUIiSMkPi9oHuwMA3M/ryr2yU66eHLtUIc+LuelF86j7LGL8TPG4PRpEUTqu
naE1vpfuTOJn8m/7s6i0gJuuXQchBIu2jqSEi/lsEeCWAHkNf7FgD4B5UXLfR/7H
nPcu2Gjlfke2ZlW3DBYaA9MjDeEulKGL3QpkQSFZWGSs/coW+Gs1uBIAomGIDPaW
yQ0Vd5dnVLU8MHUphugkAfh+7CYmG72FJWbQYE4bKLzoDqjh04tdgd/RVokdzQ98
aDysib42J7WfRncd8FeK9Kr4OFJwQkUbECA9EI81moVy20QFW1IckyY0TwzLXez5
4UJX5POFJ4bInVecYORNgMCgAqGnNK3lNwWRy9NeTfa1bJc2nZXNUYUtenP2VIBJ
63HB9ECSlWC5tWBFP6y+uhu1umaOw45+NneC25MslALu8CtaTlmGNiYnItHq+cnJ
V1focRW9EimHORqXV2hA+jGLNRqXWNeS9ZVfuh9646YhtTZvWTkxDxRbaXbHZKLA
YFKFLMaRozzgLod3cyhLZyni9uaN97RZ6UB/5AyH7ywXqXd2QixldHwlDMAxOc8k
mVSIpHHEA2dwqZDsc77yN4RzvB2WQAjtOTa9+iqjwIz4xhgoWSSntn1lA/5MWz3W
NoUeKKcY8kVjlpl2p+TA+O6BvCDPY98JHsAOmKQ8VmQvbWjkvfWT++KaCPGIOQFy
3qb7EHKGOWTAeh9zCH/u8Kdv4I8O2LgJuiZbGylORfv8GxILpwPXtUCVEy65Iwyd
QnTe71NAJVzrRg2ZMNZ/9UHLiVC37jm9asOuBJtMplppksg2pXqb+nzsBGeFHSOg
MP//gLiS5WKTDE5XwCdq4WKHAPlfWgI0Ps1YbEcGXsmqDOSnFClhyRBd9cCk28Xj
QzezUz2Y7oMUWgbNW/3v20XP9OJCnHMxIeRLuTtHykI6rRx5zP7BxNvzvI9tN52v
07cicaYrKh1Foo6m12BOoG5wrKwJWQRjijVAC91y4S3YCXSgYt9i9LC5E6hZ6URp
iWM8az5tbx3tZQizQBaEMxTvwZBoMUdVfy7tHUxF/ZIwaIHr7rFD3Wm52b7ImBnR
Xr3PpmkgVhXsNhbHc54jbH0MmMNQevOMmJ8QdhyA6kxddXXE4D/Lb1ydEiWeuaKW
JQ73jZzzMzDTyr6TNqGuIXlgeU5NJk9knjigqM0PTNgw8RAVHm/ydwKJNaeggwV/
us9V4xa0PZqIILMWqzSWGLPu66ISMt2P+IpABQlXVlINf3ZUpZpuj02Z0myln2Hw
KI0GF5wdmJTzQEPsIWXr8imkuNfuPjTKt8VbGlGKQbmUiJT+VoXA2hiVuCcj6YAz
wYNSktpZ+dKjrTxFzT4DMgg+bSSQCibdkEEqklg5h+oLih8iiVsnJumeuxquSxyk
TeyiuOHqgACNm/qDT/+FR7uVOMfeOnYyBmw47+hiz2voaBpRwZ7r01cU/byJ9Dxm
WTGOu90lyJJoinb4pxQ6ZiKR9h16rIYnSC9UCDGwGhXNeOlXDujo1jr3z2vPjrBo
Wo1qwedQ56cn72wJbAzDAj0cqWFJSt9ZFdiVqA6EKOjBEuxAksGjY4IEIeZDGBGE
1S8hJi1wVQN5oe1lfQKJwjJmEJLsJIk2IdLUbTTUSc1qpnCROVU9TVvs846r17vj
IXrIKzMqILzMs9ehPyRBXfcRGYPp3ki6upwF3OTvYsVZA+tOXaEGypd7WRbdzm2G
zyA+j2ok8Ch5oODnvnqPpFMSb1bLgoe4c7tSDqc5bsXsxYWumTopK5OYM+tClvU4
zVfG7TM+UtI4ILTXLxFbDWbQdSbpNLkG+aAKyoizMfKsFtYLvfiSMtCWZqFat9Dd
NE0Fr2IrFl/JmVuQPrbfQ86s07aOzR5j8STmJhiEUq+quAC/C7BEEhJYdORUKuQ1
gYFrFTO0wmLYydxgufyTIAxLJX2S2QuLuTeUqNBHkDG1Entbc4iHzrlUafDSb9YA
yo62OJfRMEhy+k9XvStBLBUUVvpbFqX6xU0cUxm+5L1QIRjipQVaN1Rt1zbVrhSF
ZroeL2Chlsgicaht/y0vI4mn2nFZimusX0LDEaklLXNz+A9K/CvjZMk1veebRpYK
nXBv3nmr3KN5JPZFaWaJXnEZDheSR9UB1P4exy9eqd/C4G4MfootVQmJBsJLkPbr
d0vFeioPt7uDboJP0Ms7e46qUzOmkLPwXcs8/e1oaPUMpMqMis2i5pGtjSyKe3H9
uo1h7yhrJgvjvRwiDJSUIegQZtlRelc+9IeLZ3BcMnQ6MRnj8I/4lLtIRwVFI838
W69YCo1xL3vDOYJaUg/HuoHEr06/rBJSeUCNYDV/pIAVPB7xl/MOwn7VJaACfS0B
X7pnE3aWZ2ZcM0/GVgeWOFxT7H2D2Umbqa2YfKitKD44AYbMduCfaTZkj0Rkconj
iVVjPQwYwUeqXNtnHCGEDKmbal7UV8HYGU7Re+u01haV285gaYc7Nk6gu6MmQDg9
34fYntlnFuVMaxhK7mRj7chkRjI1Jxg66BXL3pIULsYuG5p7wBybgnJHphDom/Px
H5ZHjiYjm7SdI9JDSO6C64Mxqgmy6wvQpBhzo/FCuv0sJoJT+vgYrhVHxkGtem2t
+NmGuXyKERdEOziPkF8dUedaibK/ILuCxYR3gRWfgdMCRatL3NaQA0ZlvpT79URG
pNxsoG1lQ1qHfjA0vLWTlLWO3RJOVWYl3Aa2GmokV28emQq6umysg2wi4o6xHZ0p
lF0QRymBDaqkDxOYfJe/U40D+w6Ni76Sq7INc70Krup3WQWry7sCfvSzonzZ1sFJ
ZK/NCgYFIPjSP5vYNWCsDOqHmE+hw2uAxmFseJuuWW9GvSS6/Jlgv6MJeS7jt02f
9GWAPkogU0Q200M+xOqMalIs9u+ElosPsi1s5gs6zHTaHV5JuJHCrHcIB0Z5t6vA
YXGhxYI4rONgkqJiQqrP9OR4v3dzZY6GhtTvqz4vo/9ZL/T4WswQgzVsBWGaAw02
/+tals5nPunZh8U8YaPEVW//3gjlTKVpXTS6nSwU/zu0pz0XbhviW1FfI8oSpJpN
C6O/8SCSY7otTqL6S/Y3vRW77eNRYGs2EUFsF1Ck17KKMfsQvpOu2jO4mU3Ix0eM
SSLX/zpzI5PVv/NX4OnbvoBknJ0D06HX+hhtkE+/OELM7oxHEv9pAoVfuEHjXf3v
K1cLUhLWPHszLXRcyu4rY+cuc0BHYrmEyegR2M0oqkO2OdIC6U/1KMVfzFz5e+RS
GY45GPQWhpSgjr4ZPsgul8HkmAAc1OPGB7Kd06Gug/hQv/G5P4SeRGWQsjsIFwpj
VB6DgmNfyYT65c9SwNj9ByxATXGRvKPkwx6rDnigmTf6+pPnsopK0auOljLRT7Ak
xpZiSy2GNQuDIO4qpKWHvPQ5hyc2qdBRbhbwW4GL3kN1YP44mlYvVjh5XC3h2Ki6
LwtfLBdAD2+P2KhRcCoTLskrpmsbDRPusMbw676uOTpgP5SAR2ul2adqBl6Hx7vI
CC8r0uHZKY9FXahT9sIxtirBsXXxVl3fxGwSCwGxuI+6HLJzCRFRaHh1XBDMMDzw
eVMHF6M2q1aNRVwXA5QJhQ+98ayr5px2R6vUGGemzsqQ5f4C+3GfVwX3njzJtJfB
XiIqN76ukotDi4IV6fx9hsCVhf50+TzhUFtmlnSoRsxzKMVgnf6LtvgdA84GHcsT
oTMtY+y0fMoZFTqVtpFZ4pDJYIjUbSIIgj75zORCBQj5/33mZt8TPi+N/EmQA4e5
T3MOF8RUlyDSjXoT+wu3rAoCTCBkwOAKWh3HcvkT2M//BQew38/NkI/415mqEybW
g5KQF2FS3fEiAejWEkIrqcwxIcSWAVnDMz1i2yGaArmcaRXWRcDxJperCLPwszs8
3NDqsarjS2Yw+hpYEIjjXwInt7F+JZMSURliZRMX7lwhDTE4tVtJDTZqGy2v4t48
tyg7lMMwTGIuGhbczRUI6oTE5RF8bfesv0NpFihshb/ZafnaGPitxcam9c7SveIp
3xJGOsFZqOVmpYpIJR2bNNqdAPbW6sONIXnq9x7E0Ig/Xl978Tc2PXUsPpPb7Ffh
QQoL/61AhoOtWuswGvmJm7Oa04+Uh16ngLHVovQAiPlM6EvQPVGThvR0OFnIlxfq
IquccQKS0tsZmU6e0CIBpppZjzxJPmCQxI6Zwb5+Yt9aDTfuWbcZlgVCAsFnSD3n
oyzrw3IRYzfH6Bydb10Fr/jG4xoUgX5LobRIhLCUoUqsHfxfXncP4Nr8l5k4DGBd
zI+L+OCRW/vZmnFtDZZ+4WhF4kkNYRITzP1iaKT7ezotMlmxV13mtqM5U9K5n4Uj
F5V/aYpKj0kE5BmKKFU99PlqPH0dy7F1899HqexQ/BUzABu2Uj49R3x4tsrDJUQN
K9bRNlTZ5wAP9D8IF8/s7R1oAC96WHieKPjZaTVPEASf4oZW0+sEZEm96950k+Sz
wJWoamKBh2Qk/WPJa0JP64t2N8JkEAy/GIDWIxvRwBhpKacLikD0jidrMpGthJhD
++LVQ2N4QVBd/PJ0jvUlK+RvtZgFe1HrXijUqEOIBkNchOm33YT95QhRMm7bhlXh
YruXmDTBurJIes4zQzzuWyZffRPDZiYlUCRhNjW3oyCv2RyeHme8BmJcBKDYqHw7
lfjhNDjy8ex/lb5SwuAYKJ7KIsfeS3tA9pVvLF6VbXlD2IZHfJBCBxlTWAsZJskf
Mov5eE4VzrZsKNi2IZpYchTKFenEAjbTRjIGJKztwXnKGZpuiRxHxptII4mLyvlA
OXbQb/2GMtEjmm/55BYWwXCCNzQglDX96N6ZQfIivTB29As5aazb089bS62tTx7B
laSxpwoVMvim+1G3ro1xqhZyjzJw36VZoljkQ9+uRQ03uLn1RFhZaf8rzSzuHivX
zvc8Hi8KoDbPTRC2wChKJdrbPSTXUHOkIvb36P63iLCeiQjiZQWE7Gwmnjex6P5u
TUnbtnGf7jfzaWD1Zaz1K5Cobd5mRxi8IV2TFtP7X5j/uJI36FyNUItuPG3c1vp1
U8DMH9M11Qwe4Cm9uBfd8dl0XsTOWTKA5HPMHf4N8jr1f2WtJI+Jv7yOCTFSvaFK
5/AHl8sK7oRubJd8e1n65TvVfVwSkZaESjzLnLQ2kryJIDxZVdK48tN9kDEWD+7N
BYIk2uEUA5kLBbGXhMbeB6AadYhxKVOOawkELzDdoPWlRtVheI0Ai5Ad+Bt0eJFk
E6D+ugpeSZ+pJQEjgx1o56E4dKISXZse0GbogT0Xy65N8ZOzN5jeH3yhl28ZnAkt
pM7McMwPBQvbioYQuLNc5Es6dHPeaH5fQejXVK9zjVyMvOUh6LIZWmAqQQPRX9M7
ibmI6j/LqCgQn8x7S3oLEmzomvU3ih0EVebORA5V65PiFGNtRbqimCBbZjzVUUkD
e/dXbhwAWxs8241EqXZxjxr6PV7RKz+Erdg2rmN017W9c4VqiC4Kftziu0AXnJLd
8R7QoG6hK0/9bkXij5tvchw4uS1vDw0Cg81WVaqvBfOBBfh1LC7ri9n1oZ4YbWfZ
yGe/cPbeHBeUlh6JaY3qfK5OHdK6ylwTu5lLZx4uWQWGfndBwMrtYB81AJLQ6ELg
zDN664N9+pMXRwvLR0/TNPIF6UxA2L5AUpxK8/4bEoON7AsH72uDGwnsQzrtjUcZ
63QkA1OyMLzpm1XFmAWEv0cL0Q03gVINRDuTy2RZSSsjHuttlGoBC1WvpINOAu6M
nPXW6kuWfsfQ4pz/ZYIxEJx/Lz9zi+wGqhbueAiMD/GVywepGtQLPuCeM6giHBnm
ndoGAOlw27H49lI5XQQaCc+tY+zr1YuAK0BOTtsjOT+38WLHfJ1cefMovad1HvXL
FhtxKMP/TT7vT8dpLr6XF2RztsUEfv9w/TcBFAdFADmr+naB2cBGie6gxdO5W2s+
XDXY2nj6hs9QH2AZGvt9UUuaWkX+QfooDx8E/Oxe5IC98tw68ycBDJQZJ3saPSfH
puYxMojDP8+ve9V3vN6oSZfGAiYz4AYvcIuKLq2hUJmS5XZXCAOhIkpOUQ+aXAm/
SrVNjOLOR1efJFLq9+4QWTzIygvniXHbk/xQvQX/JN5DHumIIy5W/dJnMU4v5j7W
Egd0M5BpUSYkssbUYhliROXvrdYvyUOYHAefJ+i7qR/Gdku+e263OFmyZ3tHR5f6
VoTDxfLUsO1sURklqu94DIWXV5RMZbINwCYAYEk+ZJmNWRCPYlPxt0wikHvduw5z
qsx7I5ZktKqBCPIEJofs00WI6hZUsVyHn2w6r27MCBCvybEoGYGznjExesO9HRIh
GOTFS9DSBLWtLZoznyvfB770664e2FGYbWeq+X6H29qhRUwzn0hKpzRDYlQA6MwK
H+E547HG+uqwc1unp9dPnSPrSUYysFVw27Jl5exGPCIf08Na27VcwnWV28G6VQoN
8VgnE1t1Jcby4y1hXTp1A/ZC9/VFC0Oglkr+PXscDaG43i0OscjVHyWKE16UiEkQ
Lb0XJ5KdORLAt2UVHbEkshEik3zAhWI+IyPVyu+nUS6kEjdSIKpkNrd+r74aEDX+
8ZR5QrOb9HNcp090HjiAPnzqsPNOYYNWLUuAKDTHKHnDIJvc15raCxf1m75t+min
r11iABSabrM5K2j1q3iZZi79G7mQnp8rMpyXx85tLumRwYnaIsaLWXpL7hEYbULK
Pj5IayCNEKS9Kp+/KFJgP2QNOsgXLcYADoJHGZ6IzilQ6c14APQX5Vua1UHYWbWy
RyL8mRP9WMAt4p4m0UH+Weeie1ZSVjguQRbTfjPSp25hEJ17plFedFkPisDVwki0
XUp11ywD9CT9l12CWQKk5hgHxEJeD+HuMSbatGQJXuGZ8yu9B8x9GfVi6qIaqS7n
Jr4wDS6KcCG7y4jizNAkmuD3bPnQmC2YjGpfhE2UVUROIIeRnlgNEq2TAHulK+mJ
0XEVFkVJNJf0BexiqOKzT1lSHWJl+AD17tTe1hUL1bb7erT74hObZysYOcXLi0b3
4bE42YG5+ps7AepHpivx0D3FonjWF7lm+jOhe6gFkPkpwoGj6ZFu2bJNqJSeICQa
0GtYZ1c7to3wXJrGHIpk2osEWboMwXsAbW9D+ANkTocTpyfVO4YqZcrm4ftqc1rt
648RbQDJNAZGabTXGianDsT3+rXnQJprJkoRA4lmgHkYd4ZGstbkJmK1iBbQyNh6
uoMAqdnhZT8ZXTrxY8L1ntAOngTO5JbAtvhMPizMfuIlGIWyhxAueAbwnq+/qdZ1
ZWYuONywfRS7tlFKjKoW+n4b0utKuqU3A6OtofCbVrvGwp74nVtfm8KVTU7YE4Js
82xsLa4p2/4rvAnGasJ5PuIM+q9tghg1iZf7BAb3K8SRMD3uQ2r5LvNgwxSXgzYg
lmYstO+YUj0F1ew/6lwF01jTIz1Rj5YaCvKSmsxKFBvTyvWHk8wBzbRTLHNT+00U
8+meBw84g9zhIzLnTUo0D00wOFIFYl/OCEO9TRBmUxMIMarIcTgjMSzDdQdWwK/T
JSYbIQ7rC05E5vnBZO5rmaTRmwveoJ/PeDX9sCVegSFFzj1xzcQIXTJZ5nERQpqt
dmkD8JShr4qOykEXYI7HpMRlVgea/Sjdk/sWd88N5UoP8OcYY/Fss+LK1X6S5RK6
XYcG/d7SlPKm6N46dFmS9d/RsWpF/vRc1odOJQz5gtpD0HUs/iGJ6SajzxC2eD4n
OCkY/txOuJ9zWhjoQ61KSi13VWhc+i5fxq3YBf1TgrWYOv0kZf42cn+iY5rWxYY8
BXv82PQJhY8INtQdWO+3rBo/Z+0qllUnaid/6jQT66YvGlIjk/+r66HfChmAQ7FQ
r2H+HE0IoIbE9A3h33wY1+X7KGIqaoSwPIGaZtA/bCNalNQg7qpurAPcsullMN7F
pRnPQsmxqMC1V3LAhFnGQej/HJKAjFrue58Jnz8th8Tq1VToJA1bGaPmQ7zNf/dB
6sg4kLm8UcR3rTah2gjbMdenKmlTn31FlGd0IKiNKYSEQv96Glego8s73cALuyeU
l5nC1TRo+s090WuPa/4I1IxjNFzpwZfYXH7ceYe8nr1bGvc20y3e1T3ZjCnqORbf
coV5hqR79Ls51kdQe1X0rsA6uXDxAHwTW4d5bDEe2Xr6ilV1G95yLcAY2rgHX6XZ
UZA0fQX4t7hXm7B1vKYL0WIlI8W7x/i+yOoHB/w2ffX4pNElfg6d9/QXbanTaFO4
zMYtU+JVmNjn8f2AixvsjfsT1ptLKuyve/uQsghXqRSRtrHuhuHC6RrvAsIqi5Qq
5abyN/4AnHWfXvMZ+9r4OcExI/rB/M/Ztzj4ZYPu6yrO752NuD3rRRJNu8cDWL5N
uyqwOmw6oclIhXOFKS0UeUUp3MVX/A71Q7RaxtB9oL7zGEeHaolm12OUVZLWMY6q
sYiZg5afhGGLeshYfVg3JuIdJ2PgRvgCoN3xl1lFlvMtdtJ8wUDzcoEAo9mlzf7O
1a8WPBj24tolNCL+5yU7koH7OI9JjjBUZA1UBg0gRT398Yvb8mIINa0N8xZ8tHls
nJBHrWoEASiP4DqTWj+Q93wQNuW8f0xwfRe4j9PNE22XRRpB3v0BtuUzJnEJaMSq
ZeHI/8fNNl1sIevPnBcLW6uE0GAOnbjx6L2gxchT2s9H/8m2xbe362ODyg8RjQCh
vfyR7F286HUAEaXc1aFycWKFgt5e62WYcd9uT7StkKwR0TI5ZHlBQLGP+2RcRjNI
ordRmWLNybTJpPc48Yp/gXCRYah3leVO9eQdVhLIrDcP05f2fVwhpsLzootq4vrr
42K5Lyq5F2LleaNm+HmxmYExHOBhag/TPyzxPq8yuHCYlBiOwDBSlbhV5kvEWHT8
N8520gP8adfAz4aMEvBZzWo8YGHimfJOoQDvvdgQenaNvEsfVpzeYEPoKAVRunm7
vbmu4onRZb3iwgTtyxDm5xEkMt2bn4xm50WlxNtYAmZta7BB1JhBt66yJQdgVnyr
z9t2GTPCwp9ScP16mhJyIQRwtKQWoKN1aozjyFF+82x7DCsSFU0attaFeQYNOxhN
oy57QU4h+aX+DxCbJ5XL5xVLqMXG76zj1Kwmh8x3DQbRsacJwKeUK45tUXeQtvho
yn526YPYKPPezZ9n8sHY7hbUpQVjl1LdRHo5w5vdbOqUifsODQSa3cCvO2Avdm7J
M1uY6jh56jQvFiyRBsf1OoetFV3YgkvDzrvFlcaGuzeZVry7svgMeNbjVpRbR9pn
/YAlrByd4AOjD05v5lQyDh9YVbbQ95yIueo9o6QrG6/QG9QU5o3+Q03dfeIS/ZXa
V7HNSGSoHQynX4cuIG5OIirNPwjdb+l9dlV2rVVazSWKkzGDLJMLSBaigHthlVo1
82+/vu/EoXQXmRe1FhvYpEi/ZtrgXZWudlYhZgvMcfuJLWRUFw+L6fTOz8NlX/i6
P9LRmzrwoRqvWKcau9LJRnBrGftbn8BVVy2Tak6dxmrx9sTfGmJuLurU2FJZwss9
AzrvYNIpeaoKwjy+t25IihfoKuN23ZVYzseDrLH6xc7zyqTeGJHwKdr4OR5MI5Sl
f8QzcNGCxEvISLIC/I68mVHFRQpGVFlQW3KBwIXZzhZUaGW6b2fUcW2IVDegAH+k
zGWG76QK7JyKLsmYhCUKBF5VHTzdR5S+VU11mdkFnn4Id6U/H57AHhw14hT3gz9q
ZKqWaZ9weQ3ybpWQmwEZK8NiPwhEyyGW5U88XN+oaU4SigFCQ38H17BPwVbVn7WW
Pbuj51UuFvfucGvgijWhndNKQCK4GnnTDIE4lwVgG9Vdb9pTVyXfQCtTya3fvwgF
D8zTuxqswcu03XTyzD1AbZiO8aM/GmslJuxDrshTXx66Dme+2w/i61aWHTQc6plW
a1UijMLZy0hsJh5qth2J261ZfmJpTkha95fPmdc577mWfb0feMLTmqtV+GmbUaOk
VqoGMo+2kfIlfOw1i5y/c0sQ0GSfoJta685wMoQuXwxpIgYyiNvW82KytIvE2Wb8
zaZtRf74EJshE8K60xBpoIryUwk3Qd46vfcZZDkrLzImWHIVRRvYuWuFeh6DzU6w
xgLAKcu+Uz5AL3wAHNxGhW7ySN8/ss3jztMTO5nHRuGYQzBOAk1Q1XRo5NUVQKzc
HW4RM8iUgn35gpCOFoR26HFmCz/DwLmlCkra9v9KAwKy/dxjsLO5jIMqeNCQevSI
z+7Zz81kRUlh5Q4Ah4YQFqbGAz+5K6L2izw1Z//YPwoZS9pgs+WMmNF3poETknRk
DU1ebvH4wLJ2aUDyWq6QzMxVMfDAS4q9BOiVBP2TxECdk8wNg1tk/z7sw0c6Hz5J
Y148Cc3GqBQUnCOwH/al1/0343NT0Icpgmh+ByZ0fhHL6YfyXO6roWlXlGswvfMD
+CpZVsf2r/jOPXO4p9SL8gP+I+5QQXYtQ8d3FkNp+UdACOurA0dQr/cdE3GqhIgL
bX+0CvGBQocUndAGp2ki3LtDbrN6mrTG5Bcqz7Px9pbG1XmD4KQxEN7oLvG+ByFD
j3PYVbbv6v2/HAv1ZHDa+12ddSDlrL3xS3qsnyvfkakKCD8fA8PgTfDrC0+jjPgv
La45GpJmQcUlgVTNVNlNHxnk0h4yZnW21LW7VbE3sZO3e/uozToXmSFTXSXw3Vjk
jk3nBjVI/pylXDwXkwu4nVs9tvcxuTg+wz5Jzxx49merG/wKwlS7aqO+chZ2cY40
aiXQpy8dqme+BdxuijP/0LKcsRSTA6tQQg1fV8xTd/kQd+gT5FfDde/IhqwXr4SL
eu+Wby2CRjl9zV8JlCwmWFsjiRD9qQaXiaZgwBl3ocr3UIBkTQUCKIV0PsZA3Gu6
wwOLrkLIaduF7FnIXoX8BdTs++0RGhicDQZCr46G5jMI5B0rC+2VdeOvo5SWs7DY
Lso0pApZAbvaRF1Gj06dwksv8guOH/Ap/TaEJxhgsXqRB56UPWu0O3warS6bwzqF
wUmnFdhYi7WPEf9bjidXVOK89FdUjjM/tEwmKPruXzx24n4nzK9sjSQl7aaJ82n+
BsfBTv3gb+43+j0UKF8T1ep0oL9WZleSgq4w0R622TSn3GJ4hDm1NQigCs/FXQRr
RrZxACvpjQOz+EPiGTuZABRPIhuVkGt8lwrf9eRLdWr639xIVv/bxamwc5RtkgAp
070kl5odbRmJ2zN42Vnzm3x3lrXNO2VgjmeeIMlJd3bpeLPIDE/4FABk6Mbdf7uk
h8eNCaOlZMWbpHlij46A+9Xf1fo+cqmyWX/KyZACs1uL8P7G5IP+QLnG/b2JU1Jg
JbmxORfpMCC3/qGz1DZNVeHlDc2juzmIJq1bfiVq4L0lUafjwx0Bvpz2kZ/nRnaO
0OnvYqDpr2d5QR3dJWHGbm/gSs5zHggL5ixwM5g2uBJfYD5li6tIbt9cIdw33peG
6kO2J79XlKW2ebtPbSC2M5Gf1VDcXjCwrX6/CWlpxnx8+GqKF1I98QCt0P4NU8U2
ZADJFgHy4EKczRK+SMDYhiAZWJHKQGs4SUonIu9/irzR3Cho6MQuTFb57f7qcvDZ
tG3FhY2JrtpFsRGsW3d6mCHo0KL6mJQqABruCeogyx3cXJd4V3lSKl4b6HCuzlfv
Q1N5nQY532lWKkNeaBjH9/cO1g2qTfcmlFVdTwIwRUuRTqi8wDH6xiOG6rSeA+HB
lsfsL6XZmg+SIjQ846BQ0ESQTw6ehADnK8/9GpGuEb3GcdohDOXCUI/7gx2lr5Is
syrnmLxVwag0lJZCma8Svh5SGEKDnaTlUMmGIc4+KZAkPw4r0wX8G177QRUZCvjg
fyTJaA41GiStgIe1e7e608eaBjZot/kSyGKTmAklfBnB6BI0GNXIR0Juh2WAVbhe
cM2NEmgsIK2rubQYOvP3tB+V19XMv0t5KwGliBaAbPOZTF4Pk4fx0JJ2qOgz5Ym7
qxN2lUlW0XK1CggObq/MbOpsCo9BiwcFzIHmNtTGwShxDJZReI7B4MuvALPXQMJb
j3GkLvDoxGFVOucBxlzoCGGEFGG8SxNG2KJh1uKv1x9J5fI3STxvTcjQIpxXtg6z
ez+z9KEOZjXAf7ayMaKQ0RuIUMPwSkxg6JCzMgRWyr2IGiaDwpBIGy9p+wN50Y/d
qltuPY8i9xXZVfUrck+t6M33D/aHQg/ldFjN4dTxq9AXER4OKc9Bk2yN4k9KuQaO
7AAvWRbtimPmE4JzLA39NKXaPBESyh5DooLP+6u2yjTUdX5prtxG986uiDybk1Yc
IYIV34rS2FjT13hkSw+fBNAqyJvmo5sMCLdg1Q7Jbm2up779hwmMH8Ogr7m77AIQ
rzrAeqeeMzTKtnB7sV14SArs7tUcK96sisk3bwiRGyg6h2Edxx/Wl6RKxc+C34oC
1LjdZmwPAuHMlfi3TuqaYxRGii1gJdLDbHxm60Du6RxE4w039nSkZBWoLTRx1PoC
vygj27IIjoWsPeIToaflEFEN90Iex3c/dYxunOu/pkPeeiERGHBVYUM6w5PRS/hb
v3R/UodObkYSAenJZNWBCooDO51StdnCZmtEE2Zdvlc/RlFSK15N01yLAW8ravXu
6tjOTsbq/qeSPfZPWSMYYoIdeh4gZ5VTEi/yHmwuwkI6BkyIrosemjF0p1DkSAf2
T1/aJB0sA0cavAZrEaa2oL2eZ0GHuvhbz68fJHrdlkJDmWr1y37oTx3Tgf6eFPEU
xtFgWEqPaGmoxgvPlgtTHDIwg2Q76KlM0CSZO+dLkaBqWqw9bMgNdJLfkghi1Dza
eSC965F8ja23xnCs/V7ZrNAom6rly9CwRSUCIQYMx8/Y4AYiEEqhf8IC049Fzh5Z
prvTa1ZmsDpnuzoZmbprlQKCUIDOHN/JyCc9RHWqjTrnHpE+BNr1QCwQpmWHMoRX
ADKemAgNsj+OVtmVfaGkLfZrSiTbnXrL+jBX9j0aAJqd8NBD0rdw4Q32RVevknhZ
NxLYgiVBofUgDb+gWWr68NIjC67pic9t8H42Kp5lYwZ4WmS5Atz8Rf74OgoJc3Dw
qPE7OoeMWiE98cIH0RayVhASoIHgw1HmCQP8H4Ou+JeF03wb4Ycv0QSoWxkDkGs2
9bfP5NVhcIcdVcpgzmRJeI7auDUyQfcQSU4cxrLnEHWFrDeN5qRchN2UKN7ceET4
HRO5QvKgmyFWm4uCp6leUPLAxLeip6iCfYC3lW/wZAJzTsjTV3If1XLiXYRrQkqA
pz10QktM9k0umuKYWKiOgRrnPUCZjKWYBoKx64sxnF6MdVyyDZFe6TdWBgyacYH2
9ra0qsKtM/Wj9jkTXS3j/RBNaZ+O+nGUo20yG99rPdJ4K1gAfeadjSSk9+K2E/fL
euZxOe4KTZA7ZlFa3sMtN3l8YYLxakOU7Ih/JfDg2to6XOhru0DC1/2QxwaEnKGv
NeVVvsahG3eF0yc9qtSstydvY6YwNH9+f3roKjFdIyhGU4WCMUMa/cy5vOu6vptW
JcxoH8SCJL10HjX/2KO27fwaezSP4wuXAfNBma0HKOFUPToUCzIGHebfDSLOrrZZ
btPba63dBBfZqqecMXY9c8g/HmSDd3jb8LoE3ujpXTRa6NzCahunmlsA9eS58xCT
Bpgr9e1OZfeBC8xl2gMrj2TwiRKt1s0ms73yZ0wPnipnHb+6gWF1gYAcXtjo51wI
/V4UYl4jGCWCPN7Xy0Zq9hPoqas87sPL80H6iB4oroRG5MGQfwxUUX77k17nf5Qf
IyAL0qILS7MRk/akih1o7dWp1ZrBKcHVRPJr1g7+f+v9RvOcwmGAIZn59m6n/3I+
AKqDeGhP+Yu1bqV6HSUEX4giyKi9gyH8WWBeyYPCqSKqKOZe7LRuUXVrbcwA60Nx
1XEAujbm7xOS35RSdhjZ9/yZXYe3yV+CHS0MLP4a90Y0OpOgMMGMlS+Gm889fQve
pTb3x1XEHpTy6fqCokcY6tfdqtmkrTCaT1DTt+fScSnj14X5I5i6fsskHZFfOiy9
sVnPx6LYMVc0K2yw38ZVNjylRFJYUy+O+x9mQr28jfjJPyf2k42zSUqdjKJS30nS
vrdKDugyTTzGrt6zlA4T4csEKjjm4b4atklCDhDt9bfoncrFI7jAuXSvpaNGRTen
bY32KcVY/mhIvvnitSHqMvDeqyAdRLt740/54m3P+Gj8XaxqE8buEFEcvocMoqYI
+AgBO+aCnF/1a8IRP00nTqXMXE9kJYiG7liyVSIqnkNWKcXxFraAWjmx8J47Plqj
148nRHgZVgpAEbCDXTGKvKKEniL9/IusKmX1QLGIZAhy2WxtOfKQejeO7Wf1ZdMU
j9dB82PgUVvBP5dZP0h9JZUWsqmYmHgJ0fi1AzkfAPMjs0iWYp6LUdnCbK/z5EP2
rd7v/3iB0t443zYpVwu9JTiqvF/Iv456Emf4si+O4rXFkilEs+dTAlnSa2oBmpZg
CkmMODYTq2Q79oW3TFIObhM36rhkPdQf9jgjp90ZIEE4XAMFHx6lV3xNxgLvlYm8
U64YqdyecZsI4WmWbPBKo9OYyMg3DLK9dlk2jsBWMHDosSog/rwucDGHbGsJ0siX
ug/fEc0EF8Axst+VD2+DfdQIpJba5pVATafcuMWoKFXyUyiI7Y9ZTm4JZOm14vC4
Sh34PxYJTTxtO/Pl1DVViVBWeMWyaD1MBcduxZXW0edbN5Fto0q2GredYG4mNp9r
BgbvJZs0aT3xJP49iqHYZJQTWP37dS8vZ1mQQCKyekdOqYRpCt/g0VeNyTNx/mg0
H4iU15fTxRNp+E4VSyh00qawO5w/izckNGr7LB90q+4gjUmVgM0b9xGUohzccfba
f2uTE++LFQVYpnISJ3Q42tQI/oUEATGDEv0fpk0XIdXEkOtSJqXY2KAnkYonXlUl
4OtJUTOWUrqJUNJf/ZbT88k0XhCbc5zKGximJBFD70biNJbBCukjwPlYN3pvSzxc
IPJJGb5mUOghwj8alfqOYkmB3xAZ2z95zqIoKlgfEM9Mf4wmRB6aS0V2aeFpDK3R
Voak6hQplS78TU9T9I3wI14JGmgDdHBVkSp//ncb7d5elEpJJWCTujgvkdtdgUvO
K0DiaPpZTCbiGLDIpv3sP+4PQbqaWKcfLLSPE1GW0F9Urc3ZoCN7qUCBYS1DIQA8
hPlyhiMSsNZuVsO2lUv3zpbZgUi3I3eQvwmEjuEH1lW9zm8RNX8FqZ3u6aEjYgAd
+hirl7K55aL1TjPMo9FXp95fVEoVE1xPeGOVGz+oZOYHdlc+jCZhvlpVWp8EC+YX
Jn1xb9WO1zbd9lMlSIyL1EaKaYKtPFW70sJ7QK/K2w32PHgnVjGL1yYpxN3hQYK2
wK4EN/VUgSkbzVR9UKv54FGWVYM3UmzbEJIOboFRZvxhkg9SdIIbMdGuRn21j27R
dEd1/hVx4k0mW1+w3tQY+El6sN2XWES3LwsvVux6iNvX+mQkOYXz+3184vtLku+9
ULy6iunyUOqxhwdsNz/KP24WqqX/dyNo+rRDbWfSQTP4lCWB/dw3kSHdSgVPpgue
/662X+Y/xnK0hpuj963oj8Tk8styHDK9028Bb0FT452Wiue3Lbxep6bJbY2YLEfE
e6c1XnoNFHakhOFhKt/Ss3OUmTXaMjyqCw8SUpRZLQ6SO19hHHlMMJjJr2Ey2V02
GTBNM+L/CbyDQByGdvsXd3C9AhgZFUov0wRFWH/sjQBTLmWbAkxb+uhct3grmhZS
+O4KABampNEPkR6L6WZif2EuM2JSCCO42Mvcen2bB0FF6ZTXumTqKr8dXzO8VgOj
zt0CqrCKVz1v1773pk7nJ1TgJEFaih3KHkuQgqHFq0GiP+LZxxpoY/Gocpdjm8hX
09zypbsh2srxLOMMTRCgb9f9C10dobRnMdqSNk4gQVMVaYU1MgSwkvQzsQCoXTdp
VEy8pi728oU8To0LKu9kF/7J78S8SCzSvyqJvxbkFRQQSCCgDzCl3sFit88lQwR/
NviMNHByCQA9Mwxo2ZeMwqxy3IDrhG79orDM8dnWoTuXDtbbpPAPlKUgkwtk98By
SIDs2qAjbY7Le7f9UHlEDrktH7SITaO2zcJhFcJsr/tZRoA0QdesQqViULKy3pGC
7NiYejCRC2XdufcvioS7QZcpM5zU2Wno4GUtdQVkDg32w3/kQI9no8WaMa9aKUxf
zRy470IC+nwbkwKHKLj4x1HdGtyICB41z2rNhFKuJOreCkPMnKpI/QPVAUIoruaK
1e0pznaiWIz/p9xY00xZmTL+3FbHQ3WvyO/RUHohIVDAGNdDVL+40d1/1kezEgEq
IKzBh0mUY1qBzL3Pg1UL5Q+McTogOCin1GDDa2nufyoMXpztpDjG+nusvwPEkIuC
Dm0QM4XjqWDVPk/M4JjxxPZC+aBOsf156qJQnLpnWcC8ZOVTji6zEwXSWQoj9dZP
/fZyBK7++1FsoF5/9mDYZ1k0z4AmgLxlEsMlFwfAmDsw76d+Q3DVSoSK49Az10iO
e/PXwHb+OsWl7LJJ6XnIzdsjxFv4JnX09Q2JOrzUijX9BbH4pzuzGWCaAmOaPiiB
nqROn4DhZYo2hgSVuSfIgt52GCJbJgWL35SwhAUFsZTfFKEyg7kwFup2LGdXw73+
QJ9gtMoHrdOCncCUD3Bioyo4V5Y6cLnkhD+68ObGWE8pwuvHLTdmHQMjV7pmVi3M
5kTYzW7ut6CuK8bMgacBaKqhbn7WVmAJYwC/5YtqBXNuQYIEKRU0+b2RY209VHjG
5zqOp33Yqq7GG3mTOJ6BXjUiJX+9+/5W0LfirdMhAvJeVige6mMDoGEnKkxxHVq0
y9r+NPFnMNjh+hfho09/4OeoZa3ggTaV0ed8xEswwq26dluMhetvwQrGSt6AmR5i
JfFR+bMg7Fdb0PpjqHv1bq6YVFsjJwt3sNPYKDdWKRZaq9Wgcvsc3lVxkzKKTIm3
zkJ0KZbUipTxIOMdbxfh6V8LhD++ST2P0wV7Ofy3QJwgxxJIy2PloqMHLZRwcGlL
uDbhQI8trjIQqntr5Cz+J4GlpGIbPddSc3+2MTvkFfxggcAZ69GirJH8Gj9gJahi
6UdI1XZnvsEooF5fc1IieBVnCc2oVyDjupOPwr+gBo0+ufdxloo6GOIHlvgbNbr8
kzALyvcWkUNSaszEw+kkYeWT89CXIJUhwBJq2c+whebDZntTdn8rAQfNDxJb3Iqe
Lafq/VBVlcXvF44RMXx4+PPcVtx2I/MITf1okHMLA9MDi357Uf46ga4slnoUoOzT
7XtwsBymGUvXh/CgL9Et29sL/t762sbzdJMpxzFgBYlpr+PBIpESNmFJl23W6zV6
DcAmwN8LGE0rpzOq6JLI7Hgl4rQezTU/LBkKJA79t0IEeZMoNnjFjUozOKcGkxPP
DM2PWcWj02ERmr6vIH11o3Ou+jyKydtIwd89L/6NIRXG8emzlffOAtiYLi2QSmJR
diWlX1GvIW1dP/mTbZFXdxfxW8eHxO4t73Mh/yn+ijL3/eamQo06r7sYrGlGWuJv
4QAie0DTZDE/GGoETVDP4o3xjh6rDVnbAJVE3Tc9MUxKE5RQonVzp4cdGbsc0KUt
QETHfrvaRQY+MiOspWNzhCHkajuFgIZiprxccLsJlyi31N8nrmSEhgOEzLJ76/PF
wLBmGDCb+7905w63eWFXyppKZpE4jIkVrF2mrGMFiVnmmXaBsYNBr+YX8EgAiKuz
y1w72HBIHcJIK/ekhW6rgevT6bHPsfnpt06/JkZKOkSqan+fBGtgIPFNylzjny8A
WDD7H/HP2lzTyPVlAykOwpkhKsLByEjtMEwHGURTAdim47C1yLVajdTuOWx26l8W
U4HNQrh3FgdCfv7TmSZWfa8971FXcMinVztGkEn5rzEMwLEYVvndTVrgUl3b07Hn
BbvZa2wUstulenrQgSovDJByggcfPXAUu3SZ7ZnyqDGJp/yrbDaBgK3DqwzieflA
Tfa4I3sgkfzUPAO7ZJynUq6eEsM2fmJmVW8dVZbCn/DQdzCiv8OmRkKnR30ebVut
EG/ntTRR3zdqfd5Kaj5Q7oM1rWmI4Nnc9iTeCNWcpxCorwHAJVArZ9DxZ4bvsRqJ
AVzKZXSMbTGvgYb1RTJkldteXdPFGeb7RtI6z6/ePhLvfZHABrSLrwP12LtM2Cy2
WkDRNDZDsqTUrmmcgvby94IZq5cLauSpdE/nxSGVue3YeSLQBCAJc+Bg4PLtT55d
MWsStbuAIqhUEC9IJnU59bIs+KVMKKje6j0v9oHRJA6ZDHUeIo3LFAztM4SDp4zz
XuGoA3IB+8E52FHKqOrSmaB2l+ANH7z6awA3/qWDuihnuGeH9sSMLo889eF9dfqd
SQBA/zQ1mTGVg/SGrua8xhANmWKJX4RJkvoYjEp+Cd/0DEp5iyZSoUvFFGSDtHiJ
U/JHTXOxibiccEl2DJSMHWE2bpFP4QAh4GXmCiKn/5i+nUDCU7SqQLiotvQgePiD
TeDkgOk2g38tlhHmimxBRa2Y3oGUyXqguhFTB2Qs+Q6sfkbL9tvIJZUCJcJRkic9
9GJPKpwu0Gjq0tKk4B0xZcJLR4p+Fn9pH28fN8Wwhpj+C1X1Ilv+oSDWYc1YvC0M
CSvC4zdDwT34PeETNRTBLuWytSZ9bygmgT/t1bCzwmY+PQxbwjwcgunfltC7qS8z
nKVfcqXrb+GzDiH6+tCoSKv34aoCdineN9IIS3gJVFvyw8f1K7I9guniBFTxs1n+
JWlAGOp6GHZlYM8UwPn/kSwhdwyykyo9+zdZFl18jWvctjXh/oqn3h5ekuCzUJtj
WYIsfZS4r+LT7TW5i2Igrv3MRlzFUjgBspRlu8xCAtf4FdVQ7BJraPZOujCV7ghf
cA6fXsTfESLa2d5C4E8b4tj87p9g5VpudrhLKj8hS6u04jh+FW80j0lhd/36irYj
yuKtZCLuLElZZqqVC/XGE29FK3VdrkcX0C6FSlMH5fj1km3KcwLIiOeRxMlN5Qas
y+AcVLQtTn7qvo3OJeZwrfMshLbL22limFh91aQ9V3m0uIIXuy+UqYxVXLUpm7JS
MfQNNEss7YtovlnV6j5yymS70r8j8iOMDW665gMLPFf9nY4Tot/BEOITWjNhgubm
8sFKoXrHBE9un1mm3xJJYt3AEeunZzqszHyGeiWjOlMZgg0hBdOgXKX22NGeY4v7
1oI2E4M8h/ujpg4SenbJ8KJ0MzEwxqYrSdqbo5QeelBbSlikCPmBJoSfueobWN41
bBEsQbEG14a6xKa4jD7VmQ6tPwMbsSS/4UTLA9JTYMxonn50p/hxfmskzI/vwqzA
NYFh+/3qBccHPuJydeX73yIJHt54qhUmqmP8BpUwJORpoyDnrGXAFBlLAkySaXVd
lXCoXuVly5gCRyaQnv8RCn3DQOIv4hFIDIV1nJRsRMtBxkTPKPAneT5KB1NOKIIP
+T36e7aftK3JUJp3qF5lhhWZzX+nR6fLHp9sRPhAg42gPk1r2ggFFxDNRs6m/J4q
OECSJgWCQBjWrurzsXNT8oykd1k8ICsFogM1BL9gWUijLHeQRZWW+T52u2m4FeIA
05OCeC8/Gzgb9y/uGP+IBQBQ/bWB35XVnh1ex5etldfKfv/atAzODaHthUvGutJ3
7DkGJkw4Cgjwm751hFj04/YaQKONWYRv+VwOCHVPb3txVbw843wDZugArv1qldoa
yXeCzX39ZpRjRfmC+DHKZdhDHkg8r7TZuwmDnMvq8xIa20TtNMpuC80U8Bq2JdIb
RLUTYgEhY9VKtgZvXER36gi8eT6nS/SdBDnHw4VIDS8FkgwdF5Y/Q3j/lNdzbGfv
PZVjHQJAOgPEvDC1EQCj/6vWuWHy1s36LiS5yubAI1dHajUQ5nqHf16OdsIoMCHp
ctBIhSy2+qZKBRr4Ny2L12LTaMlVHGcw8TkIyDbdYdJlp4cPU2t+sdgTq6zjtm+j
PCjva0ca8co9O1+03i9lVYNqhf5r/DEAF9GcLj++tGZE7/VTWgdmSkSn5fhyEA2a
1v6lIqLF6eU0RudnO79b9DSm9qj5r/Gs92BJ23VacRc1RBNOO2Mibl9zpudQ3j6v
I1dNbaPV9OTFSvr9WcN/qCkWK0S0tbbkENA19x5Q7Ixp0hCECpKie/rr2iWXI+CJ
HXqlwHOyfDWqJJygYkIqiwlsG4TRM6CLUETEHnk0jaV6xGsZYqoJji7OnLGYJJQP
gnJI8RllYMNl5NAq/E2F9jzRB6ZxVH2Q91wSk+OdlVmHNtupm/tBkCjLhuVb4Ksi
m8vdilQtjMoh9wwmqtIcTsmXt3DYpyvUZEda5RHGvm8eoU3A+2gStrvYQ73Jw4/8
u7Bi5bdUqp+0ZRY6e7TBWpuLDCX6mE+SR1fzgBAdxlE2o61A47dXYvo2/WfYSTsA
YIZX962+LzVk9x4p1M/dh/bJcMurgfzIRRmE/0iRBmygieRisRpyv5HLlH5F8HfT
/pN8XiD1NY4Ut8o0tqcZoyrB09Vs8NOHdukytKHssyortHnbBYk5Gr7SSf81MJds
auH0bDcgVo+8hAXmCIo5hlLFG97qck2xNXAck7jL2ekdQqOvorFVKcfI14smVu6g
wtQBhZomu4sYnsa9vwhQBIw/NVygyQ4mykfVSXAzPdog2YnEGy17r4PKLuvMytvh
Qqb+Gv31G+b42UtyHjiauQOPxAg8BadkHry5GA8c+lWUOit5ALUiUzSgBVYQiIEI
TGWiy6R86K7nQSbr9zZj3jEBkwcg8lzSskPI28wgk92wnTvX6xlwE/edY7mU3GYG
2jymPVMXVfQ6asaCv5h2qWeUwFmDn7HPLYHB81u9mTtxRm0XAhTjd61wkoCJ8aAO
0ddz74zFjYTYW7zFVi3MSAsXwUzpr5YZdEIPq/uauxoxBYHOW9nerDpsFJbZ7SLz
zWMlExVoOF5crOwYKs6vZKo0b6SxgZ7Axb4XJzYkQJkSW7tRTGmNRRDvLFPnXImC
wS9RzvgDiKG1h87zGx+nw4WsPitJTaC7ayj4E4OUPPo6Iag6MNv3JnpoJ/DDspeR
rH6Szvik8M5GKb7XKMZ3gJZMUNHaHNu0m6fX4rTX8o8Hoo3emb9oJ4KbkO/2p9ob
rXBraawQuQ4yriUJ82OzWW7GaemLKqXiEH/g0uhYcUFZM17CwLJCxbW5sNJxvfKD
I/4vIAB6tMUUjGOdKzNHkwXkoMOToYvAJjBwSgy1H/jJOo+Ecj2VjKRd2P4hKgfb
kf+38kUSleJbga9GTt2JLrZNkUptqP0Wd8SEWlRgwrLIG/srmJ8pk8O9fTRVEzZu
bk9rXP1Wq2pDhzlYumdZEjR2PZv6BX/nUM6tusALdtS1a9nsAHQ2nsNOr6ewUIes
4GgeGRVqyOhW2MTxO0CWdxvGMnsQRh4bgo7DteeYuZpjj/ooUddhs0nKgKelF5O4
EadkYEVwRTuOEYiFbWoI7d0GgvL3umc9OrAyCyITFW2TU4uhsA0lsqv6QA7FhM7L
EBNvqwNttj2sjSL4GHppqj45n3ZMazsZ1SAqjYE28O9GG42+IJUXyhwn9j6MCS1f
zwp7ysufM6VxdDYidVQueHtMX3LA9qbWHd2iq6XKrzuRbzlqzRzIEB430OgxH/J2
dlthoUaMnUqgNdFDV1yZNjU8T4lkDn0HQ6S5NttydpaFMOntbtCPTBlUwEfz69uO
Wq2+IjkAn7n1SeEztGmskqob6nxV+BZNvMnRpDZsNaxBsWpZWYwtozg5lgfNRRjm
qmqB7tVCwwu/Eghs8+URgnD1QYa+JhCpXc56+VM02cSdWPpAD6fBgv/+dKkK59d9
ljjHnQBIT0SNTMJlm+S6cYT2+IYKXmQC3PhbKSbDrpMm9cl6CNVP2Rh6tahDbIKo
EHK+L3jT+18aNtEdXD7WLdDCHMSYgYBBgk5UH9DX2o5lEOY8wZIEVuFaVhfKCX1r
Oo5h+NRVrq3SsQ9B3asNBi0yxXaU1YDWZw6DXa5z63sgdFyCbxqQYBRcytHOe41+
1LEgOst5iQrd5zGCFs/3/n7UgMfunBqtl0hvSadkRILBobaxocG8STOqj29I9sSL
1PF36v03nq+OGoK3WCvSt8uZqMo3X7wDQaxjqbzKFKQjmALPSlVonoF2xkUMB6T8
Dy4Sh1LYGeHrvp96jrc0EcZeNip3zwi6cHAJmGbrn61HfVidC2+ujB+HOwUvMnGl
TxfLwJ2Dc1Ffe22TYkjVHI5DDaeoSNITkB+kDGcuUN5Mm5GDjspDfMSpafaT6nj7
MvBTodvKVai1kMlGwu1N+GRUxed9Dkjps0NYGB3bKfV/mlMFAQd5FljhNEht7MV7
zMxPcAtLBgfTnLhVo2EKYs+bJqyWj2uKbG/DBxH+IgbD3flF8kMDv1D/VC/IOfI/
vJwg5gyV+TdFr8twRvvANmBcgG7UBpLEIWld8zeqxnp7LPGgkmkgI8WDYJJZ2CmB
HdaCjEgOQjGqkxJml1/XBGVm5OUFtoW7v+ykwDLRTp/FuA3n7TjiuR/baUih5kvx
fvoVpdRel6yfOhHZaq5nLnxlXyP6Siuf+aEM5N8/BQivdEeaYjXR+vNQLX111Bf+
QrI0YpRJXheBhW+MLWXphD2QBhhDfqHrn6jwuYMy7FjHBP+c/aCzTcssaSKJP9vR
YJH/FUDWybNNo6NeNkhiolvE474vAQc2zmBEqhvNMiDlm+4cf4O7kmIh2b4D62Qo
DL6EVnTVzjDnVChHiNV59mGCfURqjNvEYG7lRqaKyw2ocm/evUMf9nY5Ul+XnBMK
h9Pe0928Vtm36tB8e5txjyPQUcHgEh7nh8Dbys4Lb4qhjFUT6Nro3/CVbyKMQmTm
cXiJVlA64CbAB5jz19Ug4dwzLQp7S4xf2Ov5eCOtjdx6stdnFCdCIVRY2FY4bHe6
X49gfxXhR9YlcQfVxb3zegIJWTEaqgfELxd8mLQyT26jH4PBzcceMZdXUWw4QzWw
sB90Hkbwujsz39avM8CwNPppf0w3wZWTego92m1NbggVWrVph13JxrbYJPJbp88m
iyh0cVM6tAE2u8Y73bq6s6GYPALOszQnVaRwhiyaaQOoZ64JjU+72EtZg6bcsz4+
+R/iYYL1ciCb911MxSaTxk4JdAkqT8wjHykSugROoK7eXwUEyzE6Nch5KMNBp7jW
UB8vcKuzKr9rzgtGQV56Y9je/i+XzYNdhJ4odtjbmkUlqtlSoZyAn5XCF1oEirzS
PtcilYApB70QRcWVOdptkzJVS/CNFzx95IeWBihZ5pN5c501wBrtapgQhsDpr8LK
JtbLTss6iWEgTrIqWfu2I3KE79k5d3NvR5MCL1yzpFmfILmpus6CusqxKaRMC/F8
Di0Q+rStcVNFNmjKi1WOFFltUQhZHHCnzb+bmYxfI+Y8aatC1FGeC/5Ww0UH+Geo
1kUej3lrxgGBBSZAVidAd+p8ouV7AABDLACoepGeVFpG9zv5oeTqWPj5jFC5Dv7k
uAL7jCurskvKZcLIZdprSoYVbWvlBSP6kt377kY76Ih9eC2ONXTwQiIbhSHYQ4Yt
RdOzuDN0G7ArmQAKX1PJfmG227gs/se8fFdqiP7aQx5VTdGULVabokKgrhMsQb2c
7nlEApUfuCtSKnXqWtAHesd3Lr14KwOgY/FBEScfxIV7INkeyUzISNrJFybpIuyS
xlAtMoBBNokQSipFQ0lFHqOe8ZQm+iAOLTM54jvJIEFXEInGuqsEqVmTNb2jZvbS
koXrSkj9QnJOJ2jOvNkF8KNT51CEZGLzxHmu2trkGeS52e2d4hwQcmkJrvs54qYF
kKKuv8/S3mL4vatXqXtoftGcQIzwJ/ZN3rbsmLzfiEtQI/eMAS6TB7W6bDlgXA4Q
6apyXY04n5LYHqIa6pPd+gqjOqVwea4vACLY0JnRTDiftcoFfHLAVTQgULGBmuBN
rpVpomG/LCfs5/wqpEHmlvhOwXgsKk6lxHp9d1F4XI5fnT9PBBBP5asvycWCESNz
EnwjkFqmZMlHxEeHz8ex8d4oWV07DuPTqF1usBU7+bm+SMvl2irHi6hEwFXnl9me
DIFU84FOMEQFkppwg2jGfpDG8qUUjYcCAxu7PTqMyTGqnxnVCTjm9cgxYVEnqxEa
VnEq1pAYJNAb1/HX8Uf6XYQRvU2ngfAmwoNQLmo+UwGCLy1uiKGKfMf4iXn7+OFV
1+hNkeWUzPC37rN+h5DF5KeAS/dRp1eHxyvmBEmxA77HBAsp98q9urahV7k9W3Tn
VsF5I0OtgFOXBaKZkDDZQlW6oA7IHO+qjd6XxFF98y0u+jGHQPmZmZQAaNrIJjQF
MBOUAshf8k/h4gPik4mfEZTSrmzB3qCJGVwwIhncrmZzW2m+gKNOn+Grv8D6DXgj
LAYPORU6APRWKHlpOREe+SdbC225i1t8J4i4i+JPuth9o9gYDnnp3RHyUU44niLp
QV2iFBtZbT8tENGUdlKChkIigtdVQzBT5GF1lZGOFtxPBXWgKT4XIb1r2qMozsV4
rqoAWMziKnZH8PUl1cT3koqdgFNNkDvoLYxZMRS+MLyfUQ/3QNdQfFUxU2brGIbi
Ggh/CzTrst5Vz/hQ96QY8wNmQ9HF5f7+f9+sUAnI/+fycv5E7/zQhKSrc6FnUsOF
QtFO6FFXsSSn4PvdbPKL/gWNqa0MNJPYL+X66/lsB5q8ZqUpzuVc0mIaXrRj2Nhy
Em0xP17yUr5QdP8aaAFEPlT1+9U9arKwnzOTdRZFrsD1LWhx1D8Uqd+1Oulst8oE
LjiLCAzW9hPFNayZ8KEPnhuULfmr4zi9KmCvBHxYgCvIvYYBLhnhFZj9Wm6yy8dj
BrMykn856bWUzQhTgdI/KF2at1LPjp6xFOGYIv+oVNN2cpXz0VKqXsHXYQJNk7He
p1gGTWXHyKER6LdqQAh95sIExP2oC8qYeorAhzeiEIQo7t1hm2u5VvW6kM0S6WIz
pa8dPfvZmmm14PXunOm7lceTFs1yMnxtPpqpEZAB+mnWdq7dRvUfqVx6h/GZc3XJ
qtgjJ6oBI2pTfKdrdWEEorzKlAnUqtnRJZ6DsleCyjPESAvNFektclAbm77S2+Nj
gB4OKaaE9XQTaye4JW3TLrK3v4KlevWxHx+Jmzx8xL4hX2JdivuZMw+evR+yflR3
p7lqXcCJ0uuoQG6EjzC9Z06HE1X+sAr6airOQ+robQa4BKEy7QKpRGXCa6ERxZBm
oguP1KmHc/XvQpDzipNWiN9XUVBOJMm6RXMJHJEc5cCENWa7fFbIUyA7SX0hjOF7
I6wm9k8SqnZbDH7BOi3NmjtU2luG/7rUdGgXSZ7lgartAqnPbNvwa1FwMqwckW8o
YC90hBroCtN/3ddHU1ioTMVv3CE6af/4YO+8z20l2esigMGE1MNNxN6U7bHylB5W
IPERMCaiJu80oK1f8JxOpggt6OEPIe8HLoq+o7mnH8t7Oj35cC1Ji5cQ1/+qJABH
2tOjs1c9Q4/BJx76ak93ryvEOOY6fe9m6KOnHj8faX60CZdSdmUn4CtU31ryS2Gu
H+d8G56ewGSg4xiWP2UAxysn/HnOB+uFY/8XRLUvDl3PulLQyFFsexNAbtf/PTRV
kog196MasIID6uPiOBkfbTnF6fOM5+Aojji1tKaLVUjtIJYL8KCnt6inHwhM57Ls
tP2AILWk5oJch4pM1HcFpqRtne/lWJN/uDz9WsEwgL4kT7FT6Qhpv88hBuaLISRx
IDPXzOmHWM1ELQOCH0CW+454QdmtyrDcnRVKM1nvbjHABbPOYgPRdpJD9O6wgVVT
Fu4FNf8isD/tk/1aPBb13m1rz0AYpPxWNKa8IB4MJmaklk3z7Fy0kfRiRy/nVHS8
YtjxZtWqb0+JP3DPovgINbawcz1DrvMsIBCVuUNjwGCUgfoSD09qolgx3icEoRy+
ePXTMkHYBQhZpoedg63FeYH2XwlmRD1nQ7QvtQETk3bAm59oHmPLP8MjU+GISQj3
a/OUoibxEyrYWwLu7eZRGMwfN3TMh5Nh5RTxMTGJ25WuAEk01R6HwKUNcAwBx+5P
UGXM0eM05woudZPgBQnTz0XIxR9r6X9rplzPIitj7CgjyR2i7OyYndwzYZgIV0Og
R3stM6WL+2BcZRNpVAs4T67KrU3uQTnw7T5CNGhf3EIpaqVvhjC8yw9Qqe2LDjhf
nBZfYrY5h7S3TCd/d08Wz5OPTt7vIlyfIZIGliR42IncMMa1m0Loz2Iev3Nj0Xe1
ZXeEoO0U/C3gGgiCn/SSWZU9vB6qcWBycusRCmO1wxrDhR8jkXk7GdJEwLRFdRu0
ObEDwm+EoQHmLXihz7EtWCxai6QypKb0UBxOh5qugDPysMneRuVHFhlWACFMN20U
WgEjw9+RHrsV1FwLtgyGqjuU9v/gCdnJyxh8vUJipJhgIp7GYBuXHWl72W5SNoQ5
HZ0hnBEXDpeYBePq72BZk5ZCLK97qSkZpB1QbMIximaHfrDYDfkpaFpF/Hu0MbLd
YGO30TP905EMBMsOUm+2rXsM4ifaODqp+aQwm8xinkx8Yiq4NePG7cUQXbqvkHT2
ZSmi3M/gzE1ugbQS5FSkulv7NtOm5HdW60o9Lqe+99f/kysw1VnYXC/MSQX0ff6i
IWiXQZqcsLn9aAszuk8Ob3xraz6nrOFdmsMDX9rQ+bKHd3pjD6AdxqMIJ/SkzDEV
yxaZlWPG1REFI4LYI/HZ3KmMqS7T4qJvcMs0o9wmB2K6+VUgv2upEv4v3PpD4xD0
77gsvj9aVpZMn6VZ3Zb+O4ukobqbaCjcHC3kprTeuRBgYNRsmTwIlZn9rEjhyR0C
00hZ0DZbib8tq22QMDJDUb+ykbKDckoJ/3RQVu3JnHY5WY8DM0xrjkBob5jcde5n
r/s4LPQAXLDdQtBSqwODqEtFuWuu3fHvaPJuG6/s2GW4twytbCNCZ1ZcSem2/WvM
xy0qdvOW4fESSo1T4dGp73EKVFu0Ah9syCKOO1j02GQ6AK5JxQT51awcQVvXieN+
553jk568acTVV5KBc1Qwcxn/zvxEDwRczOGFdKlgYz5rLHo5Ufschu1M+fxGF/QS
oBgkpvglBvEtI5xTlqb1oBXD9eV4WGPx5odOCBscQLs3cOPUBerz654g7Bs6hvi6
pySmUHbzEhODeHn50/5vz93t3IzV+Lx/lZ9rW5AX17/QiKby80HG5eJ41e07QDf+
OO5s7Czw8gi+zvGWuqv/LutI6gRWgZ1VEx20iv+yDZOz/VNbSuq0EQOfD3ZE1Oio
SmNQ8d51Va1kua/hICuaYhh3fxWeWqT2LWlyM9GsrWobFLpD/8jttn1v9AsfPr6o
MhPwSdO+UkY4+XD+z+BDHCBXiPu5o9402W8/56riXTF/zqmI/7lK3xNLT47da8Ph
76sk2UFB+ckHXH5xqoSfCxyQwYDpeVFQ/yGmiKEmGW9tgMBzyw/bniQlVj6j3Wnj
mIOWjvpmGphpfi7AFTA22StTQL4lxs3rr8gjTy8GRSbbDnC8nI1BcRCSUU9LIe+l
2BMEViZ46KvThGhUalsGqlR+9kfWz5ZOab3wMOSr17iqWmtMs21dwy/bMdUaAIDK
mq4P8XUwyJ2DtvvDslIWKw/5mW7CFVkrec0WVjOVEU1TDAHgYFdYYNOUH23ODylR
IL1dRG/S6gLbWS3Lo3sQ/w9giZzCryV9Vb2x3WHof/MZcuqxxyPn3fOY++h2svj4
m3zt6EmqpUWuzuIG4Z0DiAWE9jPtAQDEzFb7Ve4XWkSKs5TxDE1OJRbqm4FFglE7
ntm6zJKmCKgGzr8RcXsHiGykA7zHc0SWmyy6g4BIg+FLiZOrL3HX3LE7Zu87Q0KT
WvZxdikjmsihwfLgoEIEsJ4B6Pi9xWF96EUI5C3AEJ0F0a3Sh6XWPA1WTnU5a5MA
k5BoMEDD0/Ulsf2oUtxCtuyY1rDR8pn5sM/92BjMD8MN39CFLMEuKlfSYJ04kbUm
aVrxc6fYdrJE3NDlqhV3OVYlPzlgrnoS0egHQdktzz8Ir2ZDsct+cKG8Lwo4tTPy
45+Coznogtm2pc+rCmCroyOWsMwVpOQsKldSZ6JZ0YcCrwM5Dj44+yP5A93RcOyu
bejj+f2V9IhhtYVfnOg75Ei6JRF8tg8x/1AN49HSxvXbkeYJlHk7L1byY3eVldcm
wXM3mRgrdbI34xncvW2fGzoQjBbth9G0JhauEbUb2/vZNnoQgalfHtfGHmJLIoJT
aWLdv6GC/nNpE8mrwioJCndJtAIvLP/3ReLRm2XQSqBbt4f0W6452Jyf+YpW5ulO
p0s5Ypg7xoWzbwWHrK3rTKGto7CpdjiYFjmPCrydXMcjDRW1ekMBZTmSDjI50//F
vTrAUb+Y8Mz7sW0tsuDKcx/gKfYPrYo7XJ+AFZAbvNqK1OkMg0ZVMmKsuLew7odB
3Ec0vl02Um9ELz4mMm0YNvoNcLPh+vPcYzecNY0/lhQxhYQLcz3gaJIwjIoosU+k
6zQtpzHMVxSdSho+CYMNmhn69Cx/uNXTm7eHOucHxxJ/5uOkucD0NvSL9KbupyOB
u3RPbWD5W3YK+7394/kL6KiehM61Wd14UdoGX8sq/6U0Z70Zgtn8+IzbIws7HSIa
VhjqTOOhpn7FeEF8tnGLN8//lc3s+9iYmLRBlgvDcmowmCj9/7KiAHdDIQGVvjEH
Z0zRMKJ5h48lz4Elk2yc4cnQuWVmumnOB9A5TZ42oZSgbswKxTD4YEIs2WK/Q5IP
0xrXHf3/RNWTDZTpuovmgal6LOAwQlJ2eF5gQYKBlpAnA34YPuVBp6ENaQB8NHsI
BZcVJ1aajtvESGktcGhB8N2sXsKsHCX0NApOHLe329cgjSeKWmLYa9VSNt/M+Rrf
WAcHq+u+fq5eMKgeWwLoKkMCXJJScQklKgW59jKOLlXvcyezcap1HW2yT1RNML17
FPBx8g6LLurqs+nUVRSuH7niXwmXM2S3e1oUKC2ljBSViVSMYlrcJtVmHcMfuJaq
aYmZYY5YXRMy2UBBP90XKJppWYzSkfNuJn1fOxJWiDvfvSsegKsr5lV56cE+ZGnC
c+oEDwpwWzOkvJyE4qX5y0SdveMtc+76nf+ajKEEMZ3tMn2JlVzo67VH8Y24QhCC
gJrS0lAe7o/gtLME+BWvFIjWqni8m8SsVkcEwdB9NzoObfrl0uM8Iyn/URjCcZ4R
ewJg2O9R9v7Dz6mQ4DrcdtAwRUA5bT6Qdtu2egcx5W6IHIxvHH5D3jshSFCKksYp
WKPSH09cZTtL2Y5418NzEYRFHcYpdVFNMUmf40Idz0cPIgDGyiUTBVo5dvEEAI0F
WcEL7E41Dy2ch7Wi+Qoi/RuzU6jo4d07z3wC/w1s8ftpSvS2TSTRYtvKoPQcE2OS
vbE1Kr9X+8bUvjJ4gR1utdiewK8DKYvDSA9QWD8wy7vL9t8FbN0h4d9DlxcsfMf9
Zu1CBc0EvBXozLbycW+lozccK8cANiTjiq9UhZymhmmj/4HatZEyW57PUTVYs22k
Jwk4FQk0VC+9TsZBlxI/lhyqr6tuHBK6ME+CUIob3WxsHGepdg1EIjctMlXx76tn
lkY8CSc2+CuP/gW+wYLBWcxsFj9XEMCdsxy3t2VfjPmoktnwWTNE2o93IdoJ1YfW
14NLyFgHGxxGykHF1z8NHxfYY8vCftuQWFSmYuTj04/JAw+40A3+x9CbFw+EcBRY
J7nT85Pe7hKd/aEuU0pYAkTb8D/UGmdd7n2djOb3ONn7N/wTH+m5w2cJjjxb+2BB
8WmZBx7F8hgjai8XybCG7YShaYIbUqmQgmxdEHKW8fuwQQDv4Y+m3/FV8oogqmBW
PpalBXdJob5qfFAX47nvzMBjwb9Zb/Ab4yiNd3It2rRLmuBpd+wdg0cYFOTcqv7h
TTRYI/Mb4+QMMuo7MuyNTLsqX++cHY3xPjyg3SRBIIMSRjZbHL+RkU8ASRdwC6AN
oBeZFAZiOks7oml5VgDgxz126xdif6DWQBWG5QEWBJfaiq+s5uTdwSx9AfTCwInz
sheFq6uOJ4sfNX70KZJEXmZmBstTXOS99cmBimDADrUI5OFo4nqCX3/Aj6NA5Nuv
YOWUgwvQ/oX5gNcp5bQGrMEcE98CLgMGB4z3P5xNl9ap/fIqUdUgiChyO+al9brC
uBRKVXEgDsn6FzY+r+wTrJ7zbnQgV9VvXxHYojYK5aw8YiJp9zP/WFkuli+SJ3UC
pAtYm5byqepKnoMbj0qsp+aY/vFv6koqGJnu4eY2VYFq4y6WRHLeMltYoDXZjwXC
MloWhHXnh0KmpXEdtTqUueKNa2dyAlqZFn1Pck4Hg8itq0E7C6YaHzaeGU5vQe3b
WIEp6mJ4Zjq6Cn22xR96IL9N5cYc45aGfU6L512IQ2PB9QVv+cuEdzSaxQ8xy/KZ
e6hhZgGYrMVVXOt1PMCNDyLcKnqhK97y3eOZk2lAPHKorCujLMuX/vN41i6DAZ8j
Etr4bq0wgVloh9mwx43q4BxTBRPDMAC4rsfMJN8StZWiOgy/5k+Sx+9JPlsLRbct
pDbutrtPus425TsmOvygTs+9zbPk8E/J89zTzYbyZK287WQTXtukMwQf0lioVujH
9qs2h+vwW99gesNUEEqASf1OEn97Yo3JliIKCnm/s+hUhZqUUDLCEPsaa4Xa4ue7
YVgv7ezM2/VRYLefhi/ZPLG+v69lYMTP0zvsogLqvLuEM6WFDldnEY7eLEK2H5yV
8DO0NsnlTkTSAlUbQ6VHsTruy95qRhyjLTiITPQHbqolDiWkevTlZ4a2Nr05MFRa
CHsPTB+XCIpY/na5GUrwnM3vCVbiZdLOTTOftRelDR8Spk/5IiK/ip6lJ6+iit19
nEQ+1RUfUNzr7lnwbEFS72sixqBxBc1r+Ie/Em1e8qIs+ycnXwFXt778SxzDuyyT
s0olAgwvJPdw78uSbkvQJloWR3fO5BxqfmkOdyOgfjxLXaMP3mKfvShvJIsoDADJ
g2//hqa5EeYUQfDrYerR1pomfx6Usxu/Pvew9TmRU0L3FWmo6T7cn4Olw92cXeiw
OFNIbpmC1XUbLMmznE/VYhf/XDUSvdr7hQtNJcDaeyVYsMWrJlWBU8iLqX6VoGU1
jZPguNhTsJDHFYLfOhYD/r0Z1LJcqWZJlRyC5XgS9xw3AtTC7O0gKt1bxbJiuGXW
Ly+jF2c/zK9PepPjm7noZtjXz8PixzLvzepC3gg3t3PJ5nsrtVGatYM1tvpSt8H1
EG+aLOg6MnP+na4fjOWTRHMa8fVGg6wZpX5Q2faJkIl9cVi8eGxAtGAee406LpWm
MVgl5l5gQzk72HaOIx9HPJow9iwxxxEIs5T5QRpaPAmfUZfJ+16B7U0Lgy5ZFQn+
bREPtl3IpcTKX7CD3lF05AJWmTiSYfr34Sm1CGKjUj11N4MnW+p08/A1RQKKLaQL
7ibBmkmypjNn6+O2JPzJ7hSAUJckAjsF+Es1/vcJ89uwsotpjM1gn9VGHP/WS2sK
eAC5d4d63Vwc2YN/+tQxxq+I5JUQOt2A9T0KUkNezVZ/wkO2PnPruv6DKviXDYWc
shwCjOdbEWZCFIy5ikLcBFuKjzgg8YK4qUihCf1YNusdbYce36Tz6FDtX2vH/dv+
91yvfzkk415TJLXu3UtCBCEv2pvYlFGbYgWbwC98UIEXUhzN2aM5Gi3iSSlDMaql
pIn5ZI2msEAJ3nXlnxtu+4oxVMzr8m0TdzjGGPloLQEXMhDhy2JoAp0Bb9qjry6g
vfz33l998JXLj9lID85+roS3O+NmjcuiBIm0fESb1WzAPwqYV6miBzNLzUjIZLKL
8aaE15FKK92SmwTT4AbliOzm7MNRvWz09c4RoIOY7v5BPYl9bMc9pekUCJ/YLZOa
HGIUp8rg2jDOBn20Nha9MxGM+RAMoLsSHKn8tw3mjoeFNEzodAOad1tbaQqWwOMy
opyTCARxWd1O4qMnQQHjKI7fVTY2yxYLy0LtILTBJFcShy5+gomTJF/RVIFq0Cfw
SCoZN133JHbzChj3DsJLNpwLm4BI8w1ZmGkjnxFQctFwyRtex6w1q8pOZsh87StP
l+zwbBgYGeozgA49ozKM2DFud4HINNP+dE9HKdVsiQgmjwmEzCtVNXV57NeutFyU
KQrxn3NXcU93LeZUoYQ2MXgwbbrKhXxbjFZNATTF1AiH1y9Ff9Qa++2F50sMf/0J
6CBzQDqGiDZ2vgBeWyJ65qdYcFCy9HiF5Wdic8yJyLYQEmRHnp09aC7P1jftnFmR
cFOZiNVVbVw+8PUR9PMl/WtkJNe3viZhaj7uX20c1nbocTo4fqLwoNhzszb3W0fk
a19JTDvPJLie1b17FyQb+j3M/RQbn91BUlnc1SroB3/K5Uaf8D3NFNO5LcS3tLmP
J4ryEUTccPdtC6aEHouigZjifHiZ7gArMQ7A2uEXgM93r8plcxFL1x5LuJJw52YC
r6Hu8ihEpYfO6uHYTerX5PUXsVM20ycTmClwgD5QLBGy8r9EW9M0RMhaMnMLu/3H
fog+c9UAd1dNVgjm3rOjyEqGUhHI+7KwA+1Unb3oYz0QcaJcLYXvY5vcQMtDjyZJ
Rs6T+2Os+66VHYJ2fKdrbCfHi4ujkSJ8uQxnSPwoM5ehkdTqAYjGNPNFOZSHwWWE
7++ccBFtT5US2ljaDcq7CM/T1WGAc862IFPJbjt9sVRUEYcISfX8ynBJtXKueVYK
YB9NVvG4N+WjjKK6vsHjjbUtxZO4bKtw/kc9HE9vZhL2Voi1kqhEqjXNfQpD0VG2
d/zOnMmsMJ2pY7iWt4yNduq4F9WyrM8ZPgvwul34DvhkdbvlUx/8X3DBZpV+971p
+hyWlqd56R1e0wdHGpP2qJWu5ACcmgAfLQmkqED365yXnqXSiddE7L3nDdBVznum
CEyu91N2f10aOG0RZh134mTtyYYPqu2RDwZnFebkWPIQQl2l9MJrTdRHEbP74Y5V
9aS/lLhVmwi41WG86oCe9C1lu8cAKRiKT36qg0sq22m/9+pzURxhKu3hD3rLBWnW
8Cn9T3rhx4+/oz4VfaQj+V8/dE3rLPygjhUeHPSC5N/wbZvDbezWRCePQi5GqLTZ
0N9x7ZcRoxfoboB7KQuU0uSCs/5CPvlgVMYNYUd26SAHbx3pULEW3RbN0FTeI6SB
Lg1zKJXz81uUD3C1DSh1zMTLK4GO0gMQdMWt/Zf7fBT/XrNH8yc9mEYrakIWLnZ5
2dEDIw6oOxokGIY3XDekZqhG3WC+vzK4yMQaBET7eLyyihPrX/DatRjLPVOI+LDu
Ot0jcQanlSlJLL11fder0v9BXjGYjlttD+yUP0HDIlkU8+SCFjr7NhoPngAVzUcm
LqYASmhmjRg+5GiXFL2/hJw0cJLO4AzxO6E3fASvYB4FyU4zZBvxUA62yH7Ckj0s
+6WVSGzD50u22OAnKTiBDfvb7x7K47FKR/n/WkGSHSzN/oBgJErSw9X6XqSQIQU7
2UL4//IrBDybXnSPA+GAdOuxfi0EYc/sLim39YNTfaTpkhfONAXk1XqDlcVgYriJ
e4X7Lu1AMrxqluij9zM4zgLhlEeq6gchkD4EwZM08s77lQkKTCjzMMizGQKHX49m
buO2dqwKxibT9noMVPOP7j+j/uniplwRBdNpowmItb6aqSCbGefyBI4wJM+gTaT3
zORkihgVuFbtmyz6dHWvfTe2HniPO/8stA+HbsMfG0F2GkyA7nNjXDDL+uofL9Gp
FrNA1XUzNrU9eBSjemdv39TXq+u4/gPn9DbU3Vc2aBLUE9sFFDAiOJaxWrXPWhLz
JxrmE9pW9dJuxpSYefbopzDwlAPb2rtqx1YmQCcyzR0luLfyOZeZKG1qQL/wvUBV
is+qWFV//7VxoFNAJ5n2xIrQJSH5a5nzGxyhP3ANinFbM55IQltR4xEbTIStDFjh
2qoSAUi2yjLtD6Fft5e3rjworAuwQlkdjThQwWASJp7IWjPO4ifOi5XXzK5TQ4Au
kq7cTmtHOSnuRyrmKjP2ioUQ+fQHaF05GHI60VwIrY5pi9rr6oypL/lmU3Srpyqm
0InEqPmgEU/aD/ZwjnGTifEFV8VTZwnGGktv5c3NUyEvQ0kinQHaA+BswTTiFPvC
pjGMUNtOeqMnZ5QMcLvj6IJUPqflM16P7xNVIi88HTYn2J+/afbtde4L0hIn+GUQ
Uc/ntlUFsWxHV2vaceZAzEhl6Yx1yYoBeBrG2WDef/n3LG2osfetAsu6jg9zBKls
mffaAKW0G2ffP9qfZIM1ftcFm5KD1NB/5wBhEeBS70jwvLtCoZIIkdmML+eUL4DQ
weUhh/y/WlwQ3y9+O0FYgBWQEE/ZufTgBYNCPgI205L6Dk+c6PpjBLe2HL0BNcOm
od7U5uPe61J2crfu4ASKeU8lHDZ8DXMXQOSYk5xjiwJf9JTQ05YMuJlrSAP7xJ3P
byddB5+4nPnpUQlN3pqOG86VSpuewz6U89YHhasxjUTgekVK76kgXJb2aCnE4pVH
Y6PcUGXfH7NDViyUx7RrMnon57QFlg1sSi4p3GTs84X+Qchvt8MzbQI8amEhEq6D
xdJCQSJ61LKEFGjjHP7PPJBrpjSrJGRH0nBlAfGp5mtAZvqjGSiGfLZ3v54V4io/
fM3FJkE7jr6PjEkeY5CcBTlHog4VE3frt0G1x5/IOrIVTnWXWK3dWMSU35UPGYBZ
X6s4RSd5R3/UNZymMvK3lxX4HNZbr4+1OVGaAy1lUvQd1+rz/GrAblVX4R/5Y+p9
jug0wiKxQQOvQBmMlgE93JQOQWHPMcWj3E/+oB0JWd2cPLR3kdxAotwtfXPqjkFY
m+P32zzk0PJGiOFVAr8+SPHlrpIOWjDgC0JnBuxGhK2Pfl/CWP6oEdh60wPIsvqu
2GVOMEMsTyCwkKGOiZ4RYvMFgCV8TjTouHE3m5UoMdMoQaw/+V+c8pWgnaek3Xiu
P/BxlX/CVdDMmpHaQkd221ZgZpPQ3YAqvJ6KBdOFucs/OGBd66Xq8VFioJDorZd0
S4+IFtW/KiTli1deZ2lP2cTBmHfoVuUknuY3hxdzwo9xalTNci9iY7amzASrd7lw
e7AtymiLy+uJO0eGksSOJxH/kyfGDxVs681/HHZiCo+ctFPbTlCY2WyrUbzB+BZo
eEstigfF6P513Obo+bMUWp3LktCWhO70KnV/Zk/3S6mgDbCSK3V6ssRzxhqMn+Sl
57qBUYLBnfe0uGvubKvXgrKjqTecAG9gjLLi/xcZTNCNUTMgNdZ8uiWHT5KHQXK6
ZvSvGAYTXdw/6V2ujV8EV4FtshM3uovlR3M+VoyEZw0DNeVVOOCJAliuKUJZA843
sUjKdys4AXapcd3O4DzIyh3LNblU2DUZXMpLaRROdk07KA2Xb6F7Dxmkl2GlsUrz
OnnCON0H27h5FezDsE6eglv6vMDO1AKUJF8Ij9MIO6hyhPMleR7x2VuU43M9wHsm
Vvbqi2nBBYNapNmf32lltlgr4B3HilCjZPEelve6iQRhanxXQ1Bl68m3mRB8LMkJ
0lAvHpVBAxbABo6YqoDCXcWXvKcE4XH0WG6II8aBcwe1mwC51Dq3mm54lbwPa4lX
kH/t8M8YafzKdTURfSbBTiRNNyaW9epv7O3r2+05Ps4aRdQnTBQR37OuvFNzYrPw
RaElSay60pSxj5CGtbFNESSP66FQS7zjvboiNpMo00urvJmyiWKhx5A3t21R6Q+H
425avPzX8NLZpUF/r3bw6jcRgf2bpRYOzy3tKkFV4AXwGQiq6sga4CyhE91kRthz
hpwBLw8r/XzqigxheMNrtCLmbGJI9N2ABubIya3JTVJt6h4uY0x3jyJ/cOw+vEe9
e8KjGH5Yso0P1px0LiPPzA4+dA5k5Xb8PHEAb5DRKBcYDu0N8IHaFcPeNyNZwpAL
PWDUOwsQCh1Y5WUBcgaRDdutNSpjdcQZvubrdqo8HGtzrNisRJhboVgCGIkxGWfd
ndWTQjTVS2sy3DoUam0SBxSoKXc94HlK+vrXzht9umILEArk8U0r8vVMh/Ww1us8
Dd7cL3lHgOZdrRS1olmD/zhZ1p3I81ZLiU2WyRE7i0j+C/Q/7YedoAS2yjfrWCNX
5JvDr6//BqCKCNqksa+H79oSulJXXWS+Pn5g5RFjHbnIrGauinssnX6DeKTRR+6k
ZOqpQeF/JrmRybGWVezUr+6asNwd5Zs8UK2r8bJbMecp4ftHbqI6sgK2Z3VUWR0u
GYucWFkJBZa7TbVVDRUTJsvyAlrwyMO48W6q5VXoPV4moT1B5Q4SZY0/MqLoBvgo
pewS8evRo++KdT9XhxHcFoQJq2W8/4LegYclrOzl4az+j1GZKMnujnuQvP6klcQv
iU94SaHQQPcIFJmcaMsZhA2iCe0+kCLf4mYtVeC/zXyNvcqMY+oXHA1Eb1dcAAq8
gRBi6gS4KPdnlSC3EN38HfvNHhRdCI35oYTpKcWh4rA8MKDwVl5LNNVZ4mZZ9Fnb
8ZgxWlPZZWb4ARkGcAEErjNqiCAsgk4lwQZiULbtajbW9D1CP1z8livNB0w7B85q
pXuW5FOd710ni5eLnkswpN7vUup5HOmKrpAXuymJDm8xIoXQyz4dPbNjCXu1skKa
7tdUI8t1SIlNzLii8fejfl4xechmE2o039YdrH/T+j/mj0MQZO10PXj1HVNklONN
KfXfimtSwkjjNJKZIITNUVGN7b644B1eBLQX5ofmWYrvzBbgQ5da/DfpFwPVKhdB
UlIYflQNaMrVCVTC6USawCLUxNgCr52cpaLEwgPxzJT8FNJPoyhKd+qBLc0sjBsH
gmMkTbtAUo/xNw4tN3ivWrXc2jnFpm3LZRsSmKEe8DU15siz+JthFzUJ6+a38r3D
KwybEXGrUEj1HnQL81ok/LOTsi+Inexv6E9coSbeDoC5kQ+bScXZilwpVdB1qKth
6W7d2fgY2y5Xn1F4G4Pbe7mZGj6NybCdoew1UfHehjUrxispgsdK0PS0K0vrKnwQ
i4vwfPX8BoG7bvSG+DPEGGu3zo5nfDM2ZQnVpn6bILsevHVZwBqYymbFcFdLHAXP
9MHYszviH3ZaiSyltkBqhuE9JsDbx6bi9Fe7ok9GO1t2amxnjb4pmSNXtB0m/Rpt
G2AJf64/6663zS8SJ90mhKj9UhsMDxobHQ2xldOCOLZO6q7/gfa+gcN6t6OiWlNx
8QtMFr1p2q6Y1903VGAe7dSyZ7uohwKKZXvxlrpaOTkxFO1R6JvKGvLYSRmh9pfk
Jf5Y9Q0LZ1ytL6RrfZyPxSy6t44u2CHTZL/oMrUKPwce+4QXXjmj2VA+hKDMNKPk
eZr6hfZiuApEy9pOIi+jhwp9TXajeOuW9FooeHPjEnJKCmbqJEZEMhvBZTs3me6n
enXogmYGR3dfzQuHvSX47029Qvgr1sjzR9O8DukwkdxnW+zSDZcVDt39vRtggPdI
oOgVlTD2uWfmjnp/hkaX74Hn+MSfHJUVs+RtuJK4j2Ma0EB/EgetWwMZRlLC1XYu
BUN5Wj6qk4m57/Emw/NMBcvMjnOXXLSmg5Jjs+h4eRdqEpbHwWwzkiJoKceU2uTQ
OjECYt/njNw0SgM54Nt0H9l0Pek/C2QEyKWPHnLXyWJurmM3tNbIoxcC8VLQXFx1
uX9QdMe+FO8z5X0kzTFo27ZqTkoea1QS9w4G2IGaeAWS4jTLDzAw44rfcs41Mw68
Dv0shMOk4I0LUp/8FeaqIf0iBpMbUJ+YyJSxZaSxFzFWFqQLweKXFuft55pN4o9C
8BwSg7o/4wtmdXH5nkTsbl+IFV6FRqbpOsiq+smTxUZ31EXVy17027raEQm/NGlW
BAkNQQ3YNXFG7h8C5/rpaC96WoAKSihSM1Bxg87sGXfPeCPklDDoHcOqxgdCXvHI
frhvKx46Ph+MvoPex5WQpv86WsAW+0rbZ93ngTIaDMx9mW7S6Oc/By34srraTD1W
LZiWhGlo21BX3joNbP8mmsqKhiZEZklYnNbd4R/Mpw/sK+dev1Vd5mCR3laEv2+4
8lxvrE3IkT3XIEcl0vC9Wau2W29TN5Tvdwo/ZmB3wkegLQnD3vcK7be4rckIfpyQ
8s3xHi9iN3tyqFrUH/KagIDkRxaCAXePhyAekHD3H0E5XEj4O6fMwnOgUOhX04XV
bHNOMhxzgtRFxcc34fYanK48Kbmn1n6hopPrMb1+nl04/RqU1bGUDliWfazQDxIX
aGwT5QP2V/ldySyEUivv0S2o+FTc7VEU2DQGso4HOXmbo8G1kE9+RVlkvAtFTeMB
HMzhs//6lQB6+vn1ojndJy+K4djiLef8St8r1NqXP39cnAj/OEVE8GIRw01podI4
NvNXrp85C8isCLjoc193Zetk0zSx5EXD52WevkhW0jaMcL8CpSpcQYdxtiTeb8eD
erFrPjAu5RKKCgz7Zg+pGVa+KGsNw3uSdBYsw/OdqzIfsDfzIHQ89vcQpAYlroEA
lbFqqOeZL/9L18ckENhoWjPCRq1mBgyiAThbp2PVlZhRTnF4L3IBcr9QeyR3OTP6
XQ1UogFzpRTB60e41V2a0b96/xpoC5tyIY4miB4+UD5Rv4GjB7WxxeS0uJULI0di
mLfVOvQRuF6LjgA1BDdlVOqTIegJZ0UKic9IPyxOgufr6rLF+V2LstSuImEYPrRP
SQnRK5Wic9RCWQqe+MhRY51ROPF3Kikx1Ps5/jij4CfQagumtXiYYaHueaM5NDoA
1kYqPPekPEZB7fC9To8Fy5TWPrU2vBvpFB/XYhyPgdFNj6hujT7L3yM9lo2MjWmI
XrEhEQPnkz+6ir6RDdsOIUq06l7UjTPPjyL6FVSXO7eDLDixkSs41+yr4/1bC1o6
1RD7OLcvff3wN1LV/5hRlkyL48IIAYiZ2Y10WAgJL4qf/aWBA746Hz7GfQQ6WIxj
WlJEI7alfEDi27LFZHLJaCg8uf86IdOZdQnKkeB7uKNmgLDeQYuG26fW+IQV5qD2
KKBtoQUoruBvYDO8I5szaEHtNn6iYWryvtHKAtbMNJItZCR3xNZYHOikYkxFG0px
Av1kGL6PudlmH3iRaE1UM1xN8VJpL39hxbXROmS/+4fTHyjFIHuGfeXGq64ZMfRP
iPa1YCiJCakqblLsN3ninRlHpQaQgQPdI2xeGXTfan6UFnev41W0ggSU9e60e6N+
TZ7YlL/w/Jdlo8FZEdz2i1NNrRMWG/7FfOd+b0i+MxlVt1z4TpCsf2fOgqHb+TZz
jRd08s2NDoAnux9elhQLMn3UydNxCzelbPHVHrP7B7rr77lOKcmu0YojQfc0qGgb
qMRkBXE6qy5Ms7tB44oC0r8TfZbCMOF9ifLHPGAPAy4SFVUYtKV2OyzaCOmp2kiH
6fl2RUGtsQjtAym5l4csn1OAbpSj93L4r/L+H3okif/+dYZWVcMPU726+rf+bPYh
r6EY8LDkuRVCUclddKRfSF5/6xM6oRn8BCUN0F6+WF8Lgm+FL1+fkNhMGhIwBceY
TWE9bLH4TA7UKk4Ya74162Cg16gwLX1CIJScgTQH8qQsaPQJt6mwJorgBX3aeMt5
SqpLn5BRY05jSMAh9IRGs8fopP63YqmWvEYr/tDYKh3mGm8xRrLk/O9T+uqO3GFV
qnbtsNryySkdXZhZo1FnQyxUj6o0Frw7zHErxxMTlCv57jmwNyc1FX1ruJYzbNor
H7xosexezoT3uj4rEGvYetJb2Yf7B0ZLGLWv/s0NsLNqs8dlRkRLziZeKw0ns2Ps
2FAhK544u/QLv5rrt3Lw+RQPjT96+5tbzRTWhudCoxImeoX39anPp56b0Gy+Fv27
sckw51rEYUWtaGqdeVzxegb+dxldNvdiT/o7ZejyGGE79v6ShSiN3QcTDqSLpJ/4
MAN6laxvgMUaEr1fvojQTMKJOHLYIDOaTl2Sqc6rO7pTZFrRGaeSDUxs1spiAzy4
3+sfdJUNxxWmFtp6gLgUatZRhx38he9GFiP2zpwJaLw663fnGZUGOsxsl1Wy38jJ
B00CoW2NyKM2uDt9iUM7BxbfCUCiDAWXG0gU1jQLXze038YwZ5js44ButaXIlrQP
HpoUoNuOkRziwAOvlw2TlWeWR6B+Jh/pgEH7FuOlm4StdPB5gsinSKPchFUyCEV4
9TEVkgAzK9taIAWKWAr24NjozoqTqe4d5KUSlvMs8xRANWh4JJVMI0XUhKntbz35
aSQgkWdU0gHRcHPZI29hezpRfjLlja9MKzcqSKZzUemLFt7ZcQuUOkw0vU+44Qs1
X9JlFgVOwtgaveVdzn/FTpOSkLHHx96CqyNMf8V8IayuMW8cswCaJajEPZsF1siG
Q8wLjcRx5AjMpAOgNjZVJ6zU4pM+wH59KdddyKOxDjmH/KeZNhi3ys5WVuoUKUlh
HTpUpotUyREOTtG/OEi8soDH8xnezYhJNYw3cw0+TFM0CxpCCEJa5wBprLCXPY9d
mZKVZ8NtoLfhkyHRm7iKKt+1t+CKNwC3s62MEUQOlDYD/7wVa70tThLaojruqsLh
wmdkRgtdGpH/2YQHwV6dwEZTKi1qr1/lTia4hIKq5M+/ds66/1BmWUtpRIKDZZ2q
dJ/3QeYaXzlfPzGYEsFsu8K9HAkUhuSHI1lf+lTA8GRWpTR37OWI/1WKpKwj8jci
74qv6Upm42LDbXVq28HKXh5+T04pvLNQZYIpdkkwIdaZ3gU4PhTxX4E0y044zZwV
H+/AtCz+6a7VI7e0zUuhH0bcKZG2DqHIZygNLi6GsuBv8nDhF35+ssEy2l5xMy1H
bwkFxIx6bIKMaonsXt3GNOYQkRN8/LtCEXYlQGHKnozrTYjmm9G/az+Lgpg5/W9j
toB1ccXU8MFvg9zNFP6l+XUWKgjWPg46glY3e+sywt+2Q7TOTEDt8VUzYjmtk4yj
kdvt4q0SYZ2o8nlbPLXMyysSMPZn1EhSwHPA4rGJFxCBm2I+Rd5jxIR74YFkc7JA
LkyZZ80IFPy2iK3SZkh6qJcEgde5AqvfNAnSbuZm/Ks5tzW7iUMviOXVM3loRV8o
LU9nNxL6iIXKySv0YYHSeK1OtiEu6kWxGkLbxZN9vXuC+00MvWD85HbGRjhMuUCZ
/HYXlXER/B/PF5tVRwY5Oq4jNRb6Wb1sTaykxgOm8iG1i178U9mJ+Sy1Dxy5EwAj
mKSNKeFS2AVft9qo6+VygcMTBViB6iF1XH7+OoVWpU986GvQ04BHfDklPhpaxoKm
qs1UqWsRld+7DI6CQbL5WqGLiYeRAgfRd03BxW1rCwRgTpYO/PRJhSNRvXWgXHik
U4BUweF1grTNa9Hi5l2H4R2v0hS7YUZFHJqJDhC6lbvJMewaaWgyfk/GKVhLePrF
cQw9KNJBGh1QQgpBx3cBNVIVv2es1kvuS764qMICVBuRH9sLWkl4k3VYwSmezVww
0aXADktVxKwwaAQZ7GSqhkVvcuGYwapv4yDTQ5b0r8BZvn2FUppveqYzJDT9F0cR
RJde/XIoU/eAlEowibOULQoy4QWZWjm3+5p/Ga0uQz+1XJqYrLu9KuKlg4GDITh2
bbVRxsZEUb6AY40O5r9GyYNXAy4O0eLTwCCOLKwc8x+XwDoMO+IsaMlf9E8ezD++
ojOI9SkhGzk+pyZCm60lyhH8iKkbipcFbskfTYffxnyrSl58jqIHG/4XBzNO4+9z
JklwWql52Vb0qWBSbD71d/MlcaNjivId7+R59c+6+n5ucCni4UBFvJUumCL5Jeyf
pIxRSEAwyrM2d/IvffK6sqL+Yg5jyTAEdWggsh//2gC8BTg8t/Jdag3DzSIZbpa2
jZ/BBQXGmXFwn4KzV2lRK8SfP3/lOD3tU6xLt7/OIs6vVuqN21nW3sMIDH+xLLCM
JTmN0k5YE0CQjN1ess4vlyaZmBF89U1FNCvF1J2/AmYMS9RyTIfLeREXIslaeAv5
gr4449zdSjTK2QXTTmZfHQYuynblmf1oKgkMwpsBv3tdEZd6CBHj7btK+nZr8Anf
kG8MMI0k0SnGY3baKIfAUwUweEzXeWZnDWFy+5de1n0he7a32c+U0Taw+RDZAeFC
kLOHNYZmSwCyr8acSRj56ulVfaUav2oVCe7lm8nSqet1AZAfW20fAel+kODfmKVq
4BR5L035KJhsZ79FOtVEHna8ipwRB3gWlUqHtj5n68Bz9T6bmfPDPWw4HVKUiX4z
5W5/Ft5RXgFO4je5ng3xNR/J36+QIOSTtnli26rmjLDrQDRx+hrmAeVw9J/GQKHa
C1MI9cDfMTCW1Kzmhw0fxIVi5MyzKueP3OZwt9g4vYr1oJcu9t7LyVyThBG1bTmd
9Y8mC0mwoMFmGDRmuGbVcgROVUfXMOb9KTPHriPPmGdaFc7Ko43NVJlKRLZRk5Jz
Mo55e2sPelBcREfxD4VmD7zhP7VGgghusdtMsfrtm9aWyzTQxjR38ltKMLp+Lr+H
EET/tusPdNoOQWGQEAhz7cOqHljcYxUB9Rrm6lulPb63u0ZVdvgyvGYd9VvC4kTT
AFL4esYX/+fABJaaG3aNYBqoH3+KE79SOZ6i6SoNFc+52MbZ3ud2um2I5gyv0kQd
pZhIDZgC+I+eaKTjqroeKDmh07vv4OyERXSqjr4F/HPy4baU796WQowTa5GAy0VL
fbgR43+kcKjy5TzTlP4QwuZ2zigpeT/x1NVx8V0aqxGWWNSeTukSOl8UEScCwVtR
cE4I/YXz3o4S6F6SauQZ18SYJs6j2/BGk+m2OycKpvs9raQAyD+NE6SvtYoCTboq
mGDkll+NRJ9G50qh3Q5fN1n4kbmVmaSPpEiupSYKfkStTRVOQwJ/5f8qsuTH2C12
DOWnx2PZKHSDrLCBnT2O19AJ1gh5wyqMF9UVVipm+1d92HD6tG0bg0VYQUegh7G2
Zfbs1T4O+dLndyrlYdOGM8U2D0a/Yy0MKynRRr4oEhrb+sWMWAyOS6rbMuwRmYQY
Z6+adnmB7WJ2v94nEB49bt4C6kxsm6maws2xc6ModScfNQlFmCJnaabausMJLc4o
5TY/IdUFTjdvtiQbKKIum2cdkuWCj4ugfk21dj9q0hHJJ6aPGLP5nlqO0hoJyBsL
cakm4M4ro+NMibt/pjAOOs/XbM+lWgpMmSuaXcdIAZ9K5NjenteXG24MR8uAVBnq
Zgi0C60idzME4n2iwhL97Fke1MIKNsTlD5rr0xRcFK7F1FVMPQtqb0NQ72P1WPEB
yV1pC5z55w/Xb+zdvD4U/XmNzT4fK3mbc8D/yKv8CsRKG6i1SrGMbG24aJj5UbZW
72fcrhe9m/BkcMOKWrMJJuAy9oEjQf3x93bJsEMYqUKiDLZOwVOk0gCDsNoqbjka
bClP1301/kYLSF4HSDsuehPmEmvBgUJrkmUFf/9CvhI2Ip3lQRhxmpJymhdUU5do
I3s4Gamlz6Dzo/dwOw1d012dZGfVPQmBmPo6tWG1HmUW/XATnkcLw8yGIJksU3Uy
DzynYM9O3u02XIZSAQrfO0V+LMBbnj3V7QuCP3dBmNm++MdycjFkTx+Unjtg84s1
E4JdvhZ1bIWD+zM3XvBGI3+ay8RuTKZxVLRiqyfruZ5BdpmZO3A7Ob0julKuuEqR
M/lhYolrfwaC9jqkvxQfLuq1kYTPzCCyJrOBnyaEJ1hToYZ1HhGKBzv01zFzZoLM
7llKcDg82sXZ2QEZ1x40BRLtEcUM2GbTKeXqK7ahvBHKE0HjkDtLEHrlxfixTtTe
+9HlpN8OadegOi5+T7jtkLQyJ0CbCAqAhRn20TtBNbajfESs8jhJaCRA91wScVDv
zJTDj1zKlmIs0XdO96u/wJU+fsyVgf4o4mlvIEvyrtZ1l3dehsDazyGrRE2af+fa
c007F6xZTPTW7KD8xoDJtknmYyFtjR8KW3gIwwmFpKxWulkeyHBco+gmtqrVZVIt
bTPCgkG1W8Ts3QoHnBX62Xc6plmd9bSyM3tK1UeQzTqjuL9H8IjaG3N7QfZ8wniW
yBuhtEcbXPJx4up1+jAC731afDG/tQ70FataoHTtjLvaWV0g21AZkrFGrD8NxotF
hvDZOoomvVObznhOZJU3fkSoRuooK/wC9+dz6USSHH2B1uBJ9bOlW/qTN8LikIUX
sWyKa9si6jeIer39tkQVV6YY3fCeff4USS6h7Ie1fhFJTUsejivow2crgiSmIOPf
JR6KuLrs9zgU7wfyLJXc7dkEn0EMu0PcEwApEfPL9q4pbCN2qee8ok/y25KWLaaQ
r4hm79v5PC1riiU22slrLpl0JXwcThni2Sm3B+We/W4GE67cIaTVyyoA1kO4kauc
SF13TGs5R3+Wbby9DGrBjbzjTg1rYxxj/90hNzyhKLslMdQ0O80Qsoz287WdaieN
kedpxsSwfWnE9/0Yjmfh3l2WbtlwaDiVcJS5m8BO0OQpkruaQ+ZeDr2aru5VqUGK
6L0ybzYt6Gcy7KpLgvi/jJLTTXQEmHxYQ4WJwLZ60N47PqPC/a7OrN2MDhRf3KN7
R0E4VB3eIypx/BV0I8KbogbLUK4FjDVoQTgncp5pL9gqAcEod1yW9KbTn9Fr7AoM
sqwRe4bAGWj6uRsfsQGf73KjLgLiOHkWWjXLbTerKNodDDyggfR8eYH/JMQBLRxh
oZ+FqojsFsxc0g+Dv9hmjED+OnyyIGJ4w0RsnIIe5OlqBS6aSj9VTdrbveW+nfVh
trkXE66Urv/9UwOcnd4A/p205yhK+uJSVW5Orvby6MhXjbFa5hYO01Vy9mnMPFWG
gLWYQBIck2UhC26+uXjhESN3ZILRvjRXOdmwUH76cvjvEY8lHDefgVmNuezrPq3w
74FvOlA3idr00RvGsOrsuGX/O1owU3C2WBl2iAG6vumA8RTaHQxMXD4VswTp/PvY
4IYJIwlA9zkCUxkWDVq6VJWYFmSMq20L2n1PtiN6vPYyileQsbxa5AGM+yZGiFTN
QuB65wjRlOxDv0gQFa1EiHcsFh4+95bfEGYNSeJiFEkqdgWX4LgMgeQ89/odkRHn
BUoYwq5HvyuZyrxCbUBReSFOaaDj1PdcI8ptORjWHKtXLeG7BuInCLGsKQlfu1/g
vAk6lMqXnDu3PrrRks4wL6RVa9CXk7WqWTWVKK1GM8hE7vM+bwtowqF9HQdZbhit
LkZFVc7c7YEFewmaK3jG2guc8rfy4adz3CvsUUQqZH2S18YAlxbzLfrcG2cfDDMV
mS4U8govbxqWF3eIoLSSc5JGbuWP8v9xcSm7RQGmZuxtdfr/l3dIRy9UuqpsWzDd
hY7GX3HD9RQ+Niz1tOYXgoDjqjGLpVIfBOVSeyNfEP9oAhV2YEi5nRBprOOOrmPp
t8oCmtY6Yz+C6k2yhtuzrpFcI+5ABd1WOuv8HfTNuhqDIBP4CaVOIjkzC7QD4VX/
pbSoCj74cARDxVEDTbxTfjUenZzQ08ZaDv6iF8Iay4Gm2nwXX9BNi7aPhRnr/ZLa
7EBgD6P+3EyZortsqz0v2rLp/YFolILLraTvSEQptdVEQRYt4xsKuz+A2TWO1Rjf
rPLML7+xxu7fNIZBADUoE3XooNjcTmY3sISpBb/eQ6HviWM/0BAJxzgSUZqyPklj
tb+HCLs6H9TDCHh4xko+xsRVFAGFsjgDDuoA9/FzYV2R0JliGuv7RJj9Zd+CG7Dt
G6jX/3Mbou7zJR7H1uxAZ9roYCfiEGzH0Hmxkam9tC4Z7kXgj9uO2MNbBGLbiOdZ
MZ8faK+N+2/WNLpUleiSvoivJd2b1SDk07Iw6K/qSttDXqv3D/NEMdb1kB6u5idh
4aneAVs6zSvfiygICRGigMFrnHaRc/bo4xhC6VzZ0p4aJkaUtjxq8/pcjhcMrqdj
alQ4knBA5FNF/h6+ZU1EZvncfZ/OoxWwGwVOkMVy5BZp4/gdta1/6YMcPGVDvnVS
6dIERdxYy3nzup5uvT9MaOZTMwxp34ciw+/UKQ+OKMPIeSz+Dt6i2Vhgm8T+wDZb
41tcKRG2kTZI+Og3T4og1OsAPfYovoaZpBeDWFJEalhLA8PDXWwxThkXLMBDBwhV
eCUcPL0FTetLMHS7YW+22SGrFOiX1Le5zPwZuCHrNoD78sAB0sddcCqAD/3nxuaB
XUrlpW7E9l/9zdxd8/Z8ZjazirVrReNNUg5NG9fhXzfJwtZpehzZpGcolvTFZjgA
DEjVfiwlVMjLs+Ppz5Xk18WqLoPsigXTI8ShZP5a//G1mU46imeh4ymHp4rimj9F
z7i1BpgH0jenjWo/65rwThKwnHjDBVVIHi428ymftAEXsdX/X4K8wjWVPHpNVnSY
IbtiCDamKWT/qHJwEjXPUebr+RxzeYBmZjQR8eG0WwjkIIH4ZSvCy8ugCZlsayop
BvGwXfUVvIxVcFaYX4rumyyfNyG3JCgO6YGlZhppjFaDpmKMQQxXtfiXBw60n0Gx
6lCUW/VBxTHtDX8r0V3a1Gl/Ybv8W06ErK4MW9uSng9NRXc4FTU16LOu9uKJa9sq
GYlvajNdonRYFaVA4Ns+nChRV534uiWFK1ktro1LTOTQ5zDuCHKqXFOXbXleAhHR
qFwtkZ7XX+TolA2yfFTZTqMRm7U1IWUvj8oPa7RqMv956fX3Dqi/m/J++5aaB6mc
aQfWHqG1/Rf0CLD6CpW2Hi14cHWvJoU2DvojpjJ1F5Yv7+UjBcoyuxocvTG+U/KB
TrGCp8fwCt3FpyyJ63o+x6RmrMNRlcixiM+ZsVyD1dh1NlJaTT0ammwfiGtgO8Cc
IsGjN5sxV97vXsJFlqA7Y6AcihykY/ohq5LiFvPC2eyErmj0ZQ6HEULfbZQj1EaF
DcFKZDfw2Gb+mbQssnZvm58w6htCsQicbvoLgG5d0xjWU0LRNupbFbG9F1uOPMj5
A+7ciVTuLLZnA8Mz5kKDBDOH1Y2WjdxbrnD8/vPNInkNDQzw0uBU2eIlh0zIoJ6A
97VzFUSw/Bm+epcsdkb8GR+AUJdgyCo2OhPWNQjiDdgPzl3ThJpTC4UrcTOZsxYX
97X8sPX5Eu+hgKVwwfOl5g4gzwXzKS0fiJOsSwRZJh8T7R/Es2RPwft1QEYJpyOp
gmxzoPLlPmzsNol2ix85VDD0oBaSlYGWPb9oqhhLexYcGHGP4gB8VotFnaF2NhXB
X3Jp6v75uIKciB0sHGISkvDfP9fUKgN0K/vnZJxKfPT7Y/uuJknomKC8IuT5iyei
ajvgf2+kTAaJK+dI+cdhSN5UMPhPllJ+abhekFkmn+dp7T6xo0BaU6pJUQre+/oD
H7klS8dgPiGUwXDqnC0ComOHXNy6u8xZKg4bod0XbOtzYw/Z7Hlh927P+XM7hGvH
BvM2Fbx+Fynx1eiLZHZh2fzZJKJ2uimWQmCQgcjOVMAdjvD8TK1mYYhj/mFSLa8n
CKuPLvbpojWajIhuUiBa8HYMG9nS57bvPY3GQHHcCGHgIRgxwIq0O+9BMT9CPVCJ
dcvjiX/t+ON9wlox+ofj1IIPbrcHWH38AuQ/CPGTi+qhevmINtxcBC0Yn4Xx4pX0
qEwY2FGkI0jn+fy5CP8I28Qq26C+uWIn5uUDWP1dDiDK9Uyr1iVcp9PjLT6kjY9S
fx1JwfswuGv9UcATsfciyrSMxUNBMWxlOu8n8i5j6+1D860DyP55BhzqgPrmVpPy
7kutpxoO2aK+PbrijQnJx3p2SGENiTCLf/dp5KkvJKncs26QRmId0Gmbbd6zX3+i
Er8Deqpqgh3Lz/sJkljSRnAXEWvf6QqGQ45na3zCO00ZN2T0qPHEqOU8bd2fh59D
/PGO0RlWGDCFZ3A9anCuIMW/+NpE6teDvDtNnBMEJGKS+bdQ2KmZm2fTpXYjWSXb
fKihD5majp383b/zkQDNJrpGfugKAZw0XOUJPB/4qqLZZ+bFAHm3WBbg7dWcmFlS
pkjXvHrOpXTY+ReKBVv4yLjXsg5O5RKHaB9tr6ud7yzdVw8d1/vLz7bGXB12u9ie
WjmBIBfPTPU7prR6soxyRwmhIj3KRtjqdnIdK8YjIdKYNaKzec54zAdil4/46F3D
CW6mBFzr3W5J6YN/Nv8iBB0+jRIEo3E5p4n1qZ0MDlZNRIr5HYbZba9M0vguhGrL
98pqPgu3XkOkO1VcUMzTXGTpWiSLyqoiPJD2HaoT5l9Lu+ehFaY9y+iH4khmHhZG
8N2QA4UW1rqvVQe5AiBCIoPTeuybKtZPHTBDL29shy0VGSRtug8lveAuUAYbgAj1
8lMy5tC5QXhgtWpYLXte5LElQGCk4chzS2XZCIVww29/jr+/LErWCIjesLqvMJZc
6xcEx84b1/sbY4y83h5n17rij96227rHn3C9LAhpiV6wPv/ym/yX3S0NJ5969KWT
VGDqd9H//yp9hK74smeru2i28zJuH4r1ekZ2EYN00F7NCG5LGd95yvwGIsMqqkEY
hNTIiOQJDxHrY7A5Rtw8J+0kqKKFhCRbzwO167ve6XA8D54z9V5CawYIAIfowdxT
D/JXo+gIb5xdWZvB+V9SyWI2NhZJu9sOjB+dwLG8hTHULOiA8aso/qnMgWfl+ICk
F5R9EFiMSEpXPvKJWS2Mee4sRrOIMjv2DqkDlVZwS0v71/r8EIiwA3AmRkJ4vxoO
7ytHddN030Su8e5L/XysT5a6T67GoAqwjLXq7eH8ZEBVu6P/Gw/x4d7yTIUr/wyI
ApQ3UDIYm845E15ZQ/DXte/xh1mbrKAcTPlqlso5By0qn4lOxjpO2emWiDZC6M8c
8zCEgdjH7p6+gLzbMx+HInEPQFR+HgDuNqL0b8bTDfO+10xpvKhwzT1qYLmNkjIH
pXmvqekVr+pvsmGMaU73dKoOWLnHFqn0Pd/bJRw+wwecnbIiIk3m1Gfqtw9VA8GJ
k7lfngHy9UkwCep32TwhY9Hwo9t6hpDm5ItryvAakpXvsb/oCF+FOWaLUA1N8cAB
pVYlYz29VlZO7xUUGNNmBxhBEoOqZ7I5x+1Mt07goZACva8Nz8wHEVFGVFFVl6wg
AVLm4DI8TLMqFja96b/OZWT131VCGl/4tp+NqTy5WEzaTDseexlkmoUIVN2/dIAy
NzFed0ho7rQxLggDo5ShmKPKvSAe0/7YGHByElikh90XVHjVMbUykDV+E+WPyboJ
RgX6xiGG0SxIb6wfnRhJhW37CroES/aqNjZ+5QJvkSTnC2koLJSguHyxvYer5tvz
kGQ8WAE7Bxmct8WIzALmfAanSYssbby8CvEqHo1fjErSb+/cYLOOI+qN1wcccyXj
3w3HJVPEVjOOv3021UqPaRFIsjAEEJ2H9Xk92nNhjyUBa0T8Dm1Z5RdtTzYDHeDe
Dl8+iDcUpi5k7uOx2fGaKCfcjUZwQtGd3AfmmkFhjZiNyd8Hnw2/Ci6C8yDMNUYZ
hOjy46suaiJ++KsSvXbtB4RqUpm72jIJCnef5Rt06eOc1vl2GiKabeXFCM/KfoNU
BkVipNKXNQk+xq6XKy275+EMqRVE/C49VnncsrZr/VcEp7ELu4+YKlPnL4x/urqf
1a5U9zpNkVtsW8Gmr+rbgzfrCVVULLe28/OWmDg8jIdCiGA+4d453LGRA0UupCkY
r8oPbPBlBgA81+6vlgstyhFK2X+vV055VP/N97SHA7o62HoChAdfOCZCuzdmitH9
6DpmEOOUwBtdfhWsTGLE88Jdiz5tVOz7/zipbbnwfzLBjgofL4Z3g1xHuQ1L+oiP
FvUW8CzEZ1OjBjRXeHdNIXz8BR/mBKhUhF7yNBff837bzcD+h3Ca0cisHvym+6ty
wklCGWfSiJVaoQtWLg1a/XHqHl17XGZ1KxwFXwpxvtA3iDLHp9DLysDUuHo8ZZ1N
bcw7lRvj2Yrd/JyW7yoNcwzxID6/qtJknE4vsP3/YjJ/sXRPMUAFlVtzcESecCaD
zDeqVLYyDgoDUN8aDsyOrmthGJ6fDEZ428RCZ86MQd24M/Eno7sRVLCXw5QrMV/F
Q7+qpmIEOk7JveRT9koFFBV3l5Oj77OTBxXJYpkWfo5ZlbrI4Ai8eafuvCcwzB9X
wT7WivrtcKqueAQYrnz4F2rw39ivZgQID/XsiH68KU/bnWniZVa1rl/U1gXBVXWb
zTvRyq6aDON+afF9B7r+PhTskNWGIbM/Win6IuB6zlmOCb9wQDXvW7BBX6IsroGv
+UivfbHZorkTFtHhD9hZJu7lsFfSQjdO2teuzM7hQN+ov+5gKkehputbgRyy4zai
E5kjwZ2xDrziPMluIu5xO8/4yhVEA/s+z+fKMqUrWMu7lrO73CZJBkMpGN1X3JUR
ihkrKb1P6k1rdmrFqmYFr1Fe3NEz9I7z9nNBJZch6mbsUirGcrSfc+vKVLu3h1xT
nLA99xEzJpSqnva05ICOHlk+h3iXvIxwWPeACsXPKWtwl4hA4lUpkbvNPwTVwD9p
P1ltOdxLrsTbS42BV8pov189gjmm8v6UOO+4sqxwEtSsnoLd5m2t7Nk8ezi1Mem3
IJxYTo4JaCjnqnVsNbh1iDDNIipSjgS8azaG24of6EXtHVThGWbGKDIPWxwZBZ8N
DPOtT6uUmEF89arbKz24187bZ7p1MQFExAN3YKh7ccHHpU1ZRXDgB6+La83z1P1X
HrE9SeeJAlAyapYuFVY25k6fQL4DVqhWj68/qFQr7dxXbhWPJxBN+TDBuhYzJ9zS
s2ktNB17wLHClotib5wcwqD4n6fMFfPwMENMMO9kNKmY7e8QsQ+78NxNPVbxaEwn
a1WPSoRxPlvMMTTJ6yxG0jA7o2k8MoLC4mZSclQcIh+2YsK/HwGWDOcrPEDZxS+a
6DbyUxm7/ugrnfNlGgmRyFnJ6VR1zt2eQwPD9y5pkRUx43H9hW7YJU+vGGEnvBFR
yJDYbM+miGcvTtP8YAtziOR/7sbEraAHA2+HzLehlcnGEY6YRSvsflbaspLm3E34
LJfSZCk7GZjIsFapABXqC1Q0CO4b96NMQnwtB/e/TjvNLveJf9DBk5GoNOQNhpMf
E2tl/ZUA5QwwnvOEjhpQfmETCun9g4S5rromEanQJN6fu2tawA9xj+Sz47XUwTSt
GwLYUJBlDanXeUR0LOVEZe92H164fero55G2Wu78zHF+Cp8FomdLPZsHE98+pFE4
viHGlXnKuNLvSeDO2i9XyVJ5X7BQrvNsA3Whch2scIHEDdQsNS4rB57H6SleJnHf
6JeDivbKXvaCz2F2A6lTRtrrCkNjqARVmqHxUuE2RKXZ0FyfW+E5KIppyHXrMUMb
J6taRzO5w3SGHV9WwZsJ8CnFQKy1ro4FUUWO6e3HG/tcPxo0FJhlYqN9/qLuVTN9
yqnrkHMFixmpW8SYv34YCRI/RfGM5LC0PXa4pDjKPCaXwnvOMlSe/T4Kn/PTV5tw
iTkluLp2t7VOu0Sc9XaYrtL9P/qc+dvWYu+CLf31++WXZHTSGggDGFml5L4OjFbd
436ESD6ztiC63U1o1cy5hF31xb54jRpzL3jxxUSmLKZjrFXceLhF4sCxOXpgwj2z
Z8aNEoGuKq15kfjugsgWyksZwgJ5jnLnOIrfh396sP9RU5Aui8ZEeIF8mYc8lqsM
k4pgI9pmHDIzgBK+Ef14oT/ewtAEYYozHQWcpWFmWptKTOm9snDj+hzUL+dfmaqG
oQmxO0JsZf7QM3cBHHdAaSRoHNnisOkbESLxOSgzyf+Ohp4wrRIXsE7+81DVXjwz
iyPg47lrsLlcb7vSs9dKzKcAxPxG1y+vxXfSXWKUPxGByn/X5c8Btt8eS2U85VEH
1tcA0JO7JItLYEryLH1csa4PvqYbR+oo4pd5582oEt7gl5hM3mdzae+qx7jRtVQW
ghf4rw5AZ1yD3RJLksax1X5h73+SXSbfLJ2kUFAweHWdSjULq+uXMPyCaHcEeTdH
bWC0wEOJLR0Wi7/jrHHQ5Mzz7BxfM/gnjYGVNJGbzlv2LLM1FplniOMdiw39R8H5
kbSK8l08GuY0okg/cVUtIQyFW4TseRHHgkfWRg1nIylgRLkIuLG5BN1SSFLXN8wz
LITC4sGwuF5wLl/0qoBaj92nWXDmN+w0QWaBbVem5mjCRq9iKRM2ikn8M8XzptHY
75aRrVMjklqhAGMGjO1PPaP5QgyubiLYCTcte9KMNIT791SPF36zXq7+vrsJzOv7
c6fYQptCwmvpB4l4Rmu5OK7sybIdgSOMrekrhSV4bG+nSBpVXtrcuDGD3wnXi/mW
ht1S7LGaMEkaoGso5bWt97FrzaHfkvwrxhYDlmHQR8LO7/q4EkOX00gn0DisU54J
QLBweRHmEQ9S18nJX1Tl51iIGc/A/F1bHJo5eI1TST15U/3IdvVakiY/Cgj7uvUQ
cacRs+ldJXKyzcAkAesR0KK/2JNVptLNS4OqDktpaV7Mbr/2vUzBhaeVmxanDJHy
BgdEcyDke+PsQbauI4vuUrnwHPXqWUzBAVigiGxfgVgjzG6F+ZKieDCGEgcADjOc
oyosG33ZzxNzWYwTf3AgAHzylgSh65TIma0HfOl1XMkt+/TdDIuBrgQO4+DDS0ty
DZbqr2BpiCwZe8rUSWCJ0jSSpUccEgDX809rC/SS3HzJN1xpIB+zgzEdFZaY0JIJ
nkdZnzMNOj9OmXh5tEbwQwkkZVsCO8bpr9WDfG6vqD5ud+bP5J7rXZrJtVGQcv7+
dKLdKa+DpTEFsP6m0/WtDG3/QKGieVyk4G8dgxkQIbtNqvQonxLpeTtA0f7D2Z/N
/088yQRDk166DJ2p8derVcjqhJAcfeDdldi5Zu3FQT61fZ9HEOeTk/c6+3oj01gE
mNOVcJe9BeErmk19wBNBtJvHT3Qr1hgdwwqGafwJb7KuotMFGx59LGm6CpWoq6tk
xmwZff1ekrCBf26H9wt+B85e062yy++XDhxetXYWvJxXAWDjF1zjyAjTRLRrG83i
jZ7m9VLV+1RvtItgAakSiDVSiKE46E51rRHVGBnnhnty1VrPY91FiXrr8tapfxbK
MJPxPRIrVGcfNX3l8yO2N+rmODXEtsXNItP352abE4q4OzuJ+YlhclgASjbirwvG
j79AAUk6rVTj5sN8HeXfsXmuOKLsLV6ld16WqExN3AE74ZmPD6m5SvcOtd6cJQPC
sQPuA0yWMcVpW5LHFzP3YOCJTgFajV+Y7c2pv1xCe+6mRJMTwhARnArlSknEAZia
3mX7MA5brHA4T08ARySyABb3BPNv6wiXF7h+vwbIxlhzvN9HRzH+S9S4gkxpjrOf
0h2bHbS9oknBe7TE7HjqivtILUocclwnjSKBEhKSci99VN/GX1KEY38Jmq37O3/Z
clmY6/bakdLIsynDirAyXJiNqMGENNJKaaAoBQZrsrmGpRdw/N5usvouDqGo9z67
0p1MuofM4TaDk4sRTVmiaVTBo0PTNju8Dyxjqol3OYDyAh4aVpVQd4uyuXa0pjzL
l6cuc/YV40z7dW99rOaG0NmkymnN8D9rqEaFlNopLhMsJtvlbT93MriQQqTgxV0i
txGfssTE+ATstT28DTXpYqJL3QIjRhie+8hc0ck6hDuJi06xp7WsUz/of8KlfEAP
3M6z2pEC7Jgo9zMG8cNwDRuSsT4kx1PekEn2VN1WmS6e5pUUKRVEtJA65392NElN
xKfd3i8O3Aq+nExOT+/v3OYWV/QW5EMizEGZds+tiDgLZRyV6d16vtw10l6xl87z
Eag//NZvi/fjr+OWcFdpdR3gap79nGbaUpfJKpk6VGeCL2p5XtFnxnkOuBwQR7Us
pilS5gI6UH+xo/4DGyD3ggrYCUwEgOO4sVtrbyumrPbqtnnBDWC/9jn/sRKv3r5k
n01brmoSmWDdnD5cq/bmOUEGd0zxA/GdtdRNvyqDVeUvUpTuZJdC7aWi+kisXEtj
1///bblXconIjkPzIuOhZig0KiTM4JHKgclrwhO/u8S7gkkBUiVgD45QYRbzpR/Y
bkU251GbBocC/y+43t0ecF7AS0XsmvHAocR7VHcca5JF+vMrfCdFU3sTJD9Is4ZT
2FIM0S3AsSP9oTI0cD10skck5fRFL62uOyGk0AH3Qs5zrM8tscumxkT9UCUtXHJW
W2tZBdtzUgePEIEP9XaXz5OftFkKZ7JNmOucGgRDKydWQd7gicJaANixKmJ/0nfl
eGokQBN5n00PQacMLTmd2/Ey3KIWntj05jjG1KQY/SMTWqaGwaP9qNGlQgKVdLCZ
tXTD6bry+2hqz3l42u16f8vAcAlpSFiV7S+fP5QEP4+H1r7GxC0vey8OY5A4lb5Z
3plv/FRke3AzSc1XNo/Y9AnSWctK8B//f6sETaWIHa31AH+28OszV4E464tWebAc
d6dmZeYSk7jMIPD1VcaZag3SbEQjp7Xj1yH5N07r5RNysIxB6D3gYRKSleksQzfB
UBEaYD7rMcvch5nhcqtmX640+jzlavAttUrh9CPMwpNQCUAl7abR6TWWJwjbA+Cb
KSGeS0g2Qve+HHKl/ChcBaluQcma2idjo8DahcwqEJdW3gOAj2073CnvZKS/F0HZ
YMBMupzjHeEAVwl/pIUIHEfyKL02JgxrUmJCLOTZtYOmlzp7du+29g72RgtfU5IZ
YkWqMBlqMV8pQWiVpCjvZd0yr/RNVkqZe1T0WUoZZsc2u60xhD793Qb7aOTjDdoT
I39tK5GgwCUHyUf4DfNSQuIY1REVp0aymz7yAa/EHJOtO6Z6HlX6suTNzGad2RpK
C4nS5Y3TnU86oV12Wz3r3RRCxyNtQbcyR+a8SRTgOp/zjLvxjohOZkPxzSvIb74a
Oawkoc8IznMlgmg6y1EwGo/GIfCZzPY4321WyctVszLiD0zONgKM9M2yhgYbp3RR
ySxdC+2+nnkRvhYnq69nkWS/B/qSM5QayVwCrs8BfGLheeqJpTJ3R16bZOm9ka3N
yYKz6gmuJGQbGGypQcFgL5QdPbbcmm32pXKHzBI1Myzodu21UkI1OKcPKbkrGMLP
6r7QR/RcJ+4+Z0D9HtqSpMn5WYM/+R5UHlIdyDYB6EdZiXASu6Rlu5rc2S7u9cZj
AfZjCwwU1JZnvvC0jYmY9DKTjQGbpymokWI49wvQahIs2/B25aQFxSsek7BT/773
lD7+3NcLnqM1+zQ1WgoHSP9JXTWq6AIEJC81+9JU7LXd83NeI2F8N1Gx7LrHTQKs
jPaoeP+wwQ08tNUMlU/veLPYUF+u7lSjckkwdYdsF/ApFAbBJkBN3SCQ7lfLYqs6
BHoNaGdmlQZhPe4cikAahJGS8zGw6l+HOyqq7D0f4NJHBBOh7rPhI6Y83E3JMyBS
Z4qq54WDLl15OnUTKakXfUH8YDEfM7cB9n1GKykjLlky1KLfk8kCo8Bptv7FhRuu
67gc0mtlKb94gKWE/Hhv7LW/DO40SoGaLYBN0OIL9MEaaZA2t6UJgFsiaAM7j2Oe
u23/Qn92BwrsX8+O2fgV9Xz1octVtJUTvccnVKvmaP9HkVjKfBYmchc76veAhaGO
itKnm92lI1GLT53SRa0I7BxLVVt4JoYtjWFiU6ylDArAgPjEWQ6Pn7qJZVaAx6kK
IZrnh8WCqsj0p81YsF7Rtlh04/yfMQcBZy3r5/nKckR4Adkji8vckj99xozQvb0w
NMYKp7vvEM/ZSqxzhofZIVfmCZRQsUTefERfsvX/BYMNrC1j9GddqZUD6kBd3gdC
Id6IJHZfJuNMnjjqqlrkuQ/szh6AjRu1/U+LSQNpv4n1niuRu3CoaOA0zkHElHNr
7mmAuzCMj39MPAoVyQcAkXvMem0NJXx0I2o9HtjO30k/WlkTMkyInxCxy4G7o9jS
LfjEuQm140Drxr3qUW5IP1s26dYcCcOX0VUCLbxYBkPLpQA1Ju24PuDXYKGExzxz
rfonSYAklFTqTtvnbfoW82tvpUPc8k1N5BjhWlB0Kl2zgoS8/kUElEimOJPdFqXk
Y4MkZ1y4gJnXcXtIKrEiikrV9wFREdoTOzIR87zOg1R8dOBEIkYU/zt3aDtjK9g4
4df4zSt7GI64N6+fUZ5kaGDmzJT9yMa1Jzce2aiiDPdZaLP2rVNUm9dacTLxyDP1
1PKesI2ixQs4qSce4ZsiolESgAAVErJAonGZ6Z+ndEn94HqxHtmicQj5uJSkojHu
eAGhmBzBqRakciRx1eTgh60/KfOq7SF0eQyu/HX/e5Za1wkdQ9Z/H6JHPpaRASyp
bAo6jD0auasi4XWhDIaNoXvS6bIkmQDwPlqIgi+WQN0QPtCYJ4/fgpysXAVlKd3O
kz30f2SnJb9FIixxRP6doCRjlvgdcROEsRSq9pdzhhvG+55uHjyowAKKZI6vM6V3
U0JQzaDXDGFyVigxmHu6KeUoDA+7pgLiODay5SoiA+GNnupZjZVjaCfz0HU0ojIX
5Bu3MWTyBcZyeIuYmjZIQQ2P25/o2B9YQdKCnZ73P7hsxL7d/AJXHpAo0B9G1H19
UfolroTxuO+Wi7ZAoYEu1sBuRIMuJaxRBQdZfk4P3u3njC99m+rNAsZE8ZMkYruu
B1oRJiiLMSwNQacqRTClGSO0HUR5fNonAnx3trPVP2BRsz6b8GDlzrjxqTZhbX+a
V4dffsb8B+seA3A19AsHiqO/hTeNZf809mJvg/SxzsGxioZYRlXeVPKP6GKnFx03
2TrbzlGTF+yJBfj7+5AuxeKXAnvvQT0/fqS/LGqh1skVpN8/7c4l1jKFU/0Cc7Ab
rD4Bc1PpMrUNoyuzoqws8qBUEOM8KaV8xAVfM72a2Z1YOiG7glLY1RNKp01dXHiM
ZBiB0P0sXMRbs3WND+tPE3loehC6dHmsvLJp2h225IGaiIMddU00W5AJE1ftpZgE
QlQN7WFp48TIcxXAjokeHaaJh3ADbZtsIVXG+mfbNrNNLnT6BMLldJFhoaV9OZ1I
5k3AVa1KOPhgGvnqUNJtajbDcJ9IkfW9wttyYg4mNI1FFwSdtaRSNO2mzMR2oIdQ
LpNj3kYkHftlB0GkD9WvP+vaQKj5x7Rsq2wcE28C4Q6BFcjzKmimcH7G+q2qdPVQ
rFSnNJ0Bhji64Th+2aVIdwyl8zpAn/y/vxQpsCjXfz2njkRhql34qk4fhYoCSXE6
IQxr6BrH/1E/j6IRQHnTHNdstORYdAABYsDfn2yDdPDBOvg7J29+rlwi9k/HUTxz
/m2omV8aGPtFFSHDIyBvGGRDDm3NG0XwzZR3WYfuAEgCAb3ro4z4Y3/ws9Ueos+l
A1k95xKPG3RJFm7dhqkathZneu8BJF5nN6ItyES/s/Lx+T4KrgJIg/QhT06LkKGE
q+OAQXypnyne/sA5Odvsdr+VbbOKxG6wo3jgu4sonQXeHbSoMdhxyOOEV1AGOz6Y
XpQrgogMwzF/RRB1AD61BdW9zh6ZKP29PVhMgExU3+9RfWLULN46TygRCrBSUaaF
fR+GcoI2ahDqyefSsvZnDMmUe++3JmdA/NClAPthXUfDxLHXJ1xcn/opvL9a/obJ
H6gilVuID7OB2Ghf81Ivk9XL48LaCULO/aCUvxUTuVoP5n05o2YcgcDaCBjfn0xc
BqTwCqVnPGQQkp/cYqcpzCjEA6mcx6ilh3+3+G5geJR4VTC1JegWjtibwIAfikL4
bOOeVG+NvjtdcXCbPWWfANcPgawARhXEvBpP/WLVwqQ3XNe8GfQemWouuxPFBJd3
3mKwvA5jzP3LNHZ/kzgUxxiRvZj8Q3B11NL5PajDIn0hrX/CnIn/t0DIccy/YDRZ
HlqXk3B+hR6rfKAz9c9utf6KEogDKgdh6gOHMe/vFxH55d5HLrl9dcdt0XZ0TKwx
atfhg2tgEE6PpIke2HFjY6hfg+3aFEQhUdqr0G8rgcuVW0ZSyXi+feIg12hJXu6D
Isg1FRRRM25o5P9kOXxTw1o4ahxjlxRyt6ZtW68MMldbqk0N1iAQGkayb8RyZW47
fv7OgGGP4eA49EDvuDJhyhMer0/uP7ZcFMtXxWFDwmS1hiW1XslnXjqaFsVchVIi
WuFNcuUkSfj1xTKN4FZQVOEiFMlQG2MDOFOLFmOt4WPcWu8WYL7bIUTPCkDltzSM
Jwbkg+1+jMMrIy+LFt7nQsRdFMA28X1fHjquKprKQezl+Bf7bmxm1vXOqRjcyGyL
iM1yNQrEix5KAPs1w+Fd8wgwhRg0ZTWZF3zh4bTwtmfSeDH4Gi4UHKGVAA+72TdO
pe5+IqYv69FbQQAFY71tRpKojFcjrPn1FMmmzBCnFwF+x4gW55YfcdPyq0ZGKZ9w
mTJS13m+MtVttNuHVPL9MaPl1S2bQWaKzVqWIEk+0Oe+jkzC8Qu4jJ+SKtWYvjXo
x9LIsdH1Fw0CddyY+F96kNGqgqukdZ9kZlNg/GqYPQ8I03jT5CeTZ5itJP9d07Yk
qlEG7bNS0441gAaAImBUh9m3qz7yVjZ8ib8ChETmHG2l6MqkIppzh9dzw42b3612
0dsxU0RTsm9Tq3nRFl+Yf7tlfxK1L+BF/oDJ85Aoyr7HirvGUToBxX8CAhzOCNn5
L6hbaOhn4brepGU7lRt7UW/8YWo2awpdkWMUWrer9vPqtDZrN7I1BtxnMysoZalD
eJtJrc2s3EevkLmI65SEED/2vps+46bT6o1dJXnm0EJSLM1Gn3qQlDNrJOS2PaH4
dJl3P6XIhh9kRHk5M5Xd+5dGJbv12ke/gOSRgWFd24NjuYHcEAXjq/RSVgchDPXy
4z2Zu1+1Kxq1jW75BUiZ4i4tcZPyjLxOllGEUoE1erXkuA/3bXNf2EheU0h8eTLt
ULV6485peuGDaCgIuWr6xWHzFBTjV2L3r1Me4wHAnl9sCJXfBPRbyF2TG1Yr8mSK
gkcub5oq2iViB0lE0QMZ57la+DuhObh3N+pBkRsqSK10WOIN5urgzx2ATFd0eCmw
FJXyV2KdkfISuf9X3nh1vP6F3p3wwEFQyH4zbWkS2qm6w2PZp8DeOE81cKw8+3vO
fHdm979YZVcgfztz6u5NwAmo1N6rZ601xsBj8YTUOcoTAlagDXCs587fMkJKh3rK
1d+ojh+eN8nRKrOtSeXYsvfBC9ZFMnjE3HjWjZ900vrIzuA6rZ6nf4cbTnW99Doe
OzVPckbkyPpa1+f11qNDqClxVOgsPyzIFuyYXhoKXReNQeZXlsB3Xek/oxBAFuQX
Yp8ICjXDq5yFvhj+q3L/a+tenM8hPvAXGEpP0vgcu22o4XoNuf0sf3X8vtpm6MSk
593lC9IQt//ijTCBX/62k91soE6ORqFsgizDTGd/zUDdcKDmZ14OQzN/tFZZeDT8
BV6pXGsqdQgPL+Nd3gKPFygeiJ+B6LuE6BBNheOuheC1WeT55RXRhp4DqdHgp7Mi
TCBvSM8NSCXAJzazAAQUaZ3ALHABAg9KAIi5YI3gC2VYb97ldJYzmyrjo39Iwaox
fkt1c76kuJJJxCLKMGBb0xDIa+D7KrJ/7BoUqSmLtoqCePKWYzvdQgexhujW2VSU
iUGntaR4E+45DcJUnOLcnaA/kLTCp1rzxhtbstX3TQ8gTtEFV+pwnAltN+sA2Icq
QWJlTW1RsAs9wM2/yz7uyuXa9uE+3UgiRCBo+Tunp/3bMc/CGx/MiPfjsotaxXo1
cwAObS1vmmR/N3EgGOIr7UAK8awMoMEo512wkgdKjt0KmHOox9eLB4MgnL6hn1zA
N29ze8ox4L/DyOMJat2H8SHDWpkMtL8XlT1TRO5MqfTZsFYTjhXWZdz7T0rX3iaS
2PBfHGuuCVx7Ug4r/SrVOV3RHRU/FwAh0wQB7ymWohBSrZw3f7rPEBDfLqm+7bVa
6e+ZcGGwiMIvyBUG0bIgrXau5GKzzyJYzjsiKUmxNyPPjbzKwUXrurTp+MLfcMao
mRDpEVPZ6zwm4Z2kUu5T7fJpTs+rMXp6rl5U0PSlipG4v7c9lohNTIT7Wwt+ZaJt
u5ggRz2HJbre7TRCfJ/eePT77QeA74LxH+CHe17sJ0ElN3Td+zjSz8MQ65ciH2xN
7kvS5DuxLaWqIpJ13+c/iyyIgi/sc49D2y1JPQ5Pdm/EGyIsbhqQOC3FWzrgq2IE
M9WM6qW5sRLeAlOX6PTg88LwWMbQbi9QwQSee6e06NhuTa+rsGUmlh8DGNMY3E9d
LvgMsHBlAX0ZxRcsW9b7s1jpjGZr/yKFdCDddLl/7HEjz2e6MWSwDjL76l8L2nae
OGAOfZSPIHbA5sRYIX6baRd+fhYtEo6JtQFTUk7WGCffY0dJODlc7kzwno8Tseja
GoWPlrnOnM4STnpw+kSrgSSgn2bizSQQ6qyWUOvolZI3xHXLWpFLdY6zGsgdpMh2
8GXSiKtx8Jxm5Za2k0oGU3nytM6atItJ+bcatY/IKtb+P3oWgTQUPlUJsGe9gljH
zO6YY76TbWoI+DXEhkX+te/XCk1Mw/tGHqNcjeIqsbOHXuYz0rFtBTZ1IUojtEJ7
43J88u7uACN3pqD0cuzcCIJsaHfGSheJUASolxWwqXTP/BviJUIj6Awtl+fU6MZA
Z+8L45mgfAvEjfzOv1kZprLaLs4OuZZ0rHxPECpjxDRwllSa4+vTaVE3rYGloIcw
dQFqw7DcMEZ9UnOKtcSkPF4o5Hfd5s0MI5tmUWUeJ9NY25/3CjDNOd9E562Wt/EW
Z31ail8L0n9eTJ3XxyxciBMmRXkVv30gR61Y9zBloiL62KVZO58Y8SWWhpaSxUOt
RYBE9CIN2n6C1W+kVIILDgVcUri2GMootI4O5RdpEVbgoD1RZh1++cQP+f0NTMQ2
pe/6jqOyQCpa4bOj0enG7evWMhAn9a9RSnNifm0nqHXm0EuCPli+Yx0NpTr74vu6
Xgh7gpTC1SCi+wSbEUf0q1PqJUL6DGcuURW3P9KH2lck2YTuMjboevbm4B8iQDl0
5x/q5izEgqfQNNbyVxvnlWHcnAv0zzQfC1nZRR5ITYR/tVHiwR80kKLbzGC+BLNY
4NgFfZqUuRjyVWt1s6fLW65IP31mPEyFsiKnHgUnZAAu3HGtdCz7Ha1M4F9YlNA/
g9VKHA4eDh+rDXAl3aIYbuhLgyNRbeCqOjp9+1SDwqDtr6VKjowOlQE0AzRdAEzK
YN/WUYykOSC8Lt9ycy+ciq9hbloKJ3SRE3vUX2+iOL7x+3bwOwjebAQGYsMjnW7c
uPvVysnoai/FEWGkIXUHykj/pJIpKXpTh7UP7s3q8xhoh0tVfORFuq2o5AI+zQSQ
mysNpxBgH+mNosD/T2T0JclewHpFmoa3xirtWX0Fi1EoQ5DcddRlPyn5J/tOQ7Jj
A5ZFPxriEwD9kiy3OErlMpzCmFvdcfla//dw+LVHqb0Dj2REY+JA2Yixrs0I553q
NbUCC8nGQYG+XONtSKvJmS5RVEqZ1cd5w7DQWMY9WDtwRh8l/XYcaz3l6c3etYOP
fGHpcR4oaXDCcGxBT2OswaII9hqhhLnKIpuaPfprZFIJw68lBfGz40T92H8A71tT
napT8uJpXOzC+gjKLlFQGrhxe9ajp53aagVNLFb0/ifaTjxlnuCWxXtUR1X3WI7R
wWJ17KahW+6wQJ4goRkKzQM2dkLlEQqfqO0AkaZAv/ovHUhQmYA7uL8NoPDkxvFR
s6kzDpnx9Wln5cXZaHrpCwkJ0IE/4gk3BmjugNF28IXt5Sc52yoR8g0XAhX3YbGZ
oGb1Ib8zgLYfNH5x3ACxWtcEdiqPBBa2rMVZa5xEBB4WoDtRCxu0GOcFKxNmWONb
m7fK5BxUvaOKul4xtpC5Kk1O1Ra2dRTcPIsNNO+nl4IGllM+3+wGueAK2PHrSSd6
cLDHRrJ/Cpev6fTmNsTsKIO9q5OF04REei2zhDWzFVMWOqAEu3PyVimvWipr0YDY
7VRH7Q3uDGFKOiQU3sZhSd/V0B7/TqoIfoZkHdrGc+ioR8YBhW+7o8viUDOrIqNP
xZZqZvscjYji4ojaPfxj4d3GoszOXw50QXD5fTBybnSr06I8loFRhFO6JIdcW0Oq
ZPpm27E3Pa1MVorKQ/UtbIb9qLkhebhYK3d1jZ9LhU2sHleLKRhpq0hPtVMS3/fp
JwDqR1eVykWb9PSOUBHlymwqOF2XYBc3ULhyBb/xiyKoLorTJP2ApoJnMfTfmXop
GJPQQRqjOawpUK2IstOZ2joKn2emD0nWd42TPp165t0qYWJfw5/uwWmXFSyA1P94
1xPqz2A6aRR6SGSSyaOA71Yuu25KFR4KM87QhIO5VmFAQi5Wyo+8rYMjqb7zW5M8
W5hvkpSOZ1XbXsHcx+bR+RpU4KGtZsA0CZ7O1zG7FbGa04qP/wLYI/gAbUjKjpV3
s19IgLJBWcZ51wNeK7hizLMrEY3ewxOG/SriqbpIRwN5611Pz/kqkD2t7Q/AUBtS
LouhzIAAdmV8XXZpwyEWs+p+sqN+P9v7BVdmbyiokZ+kTiYVFTGU02frATHUrbZz
BVGasBkXPqdciqO5obVKgXZJUcjTKJ/sSCODhZ+Jr/bvcQhwv7+9r1ZSpL9vcsFN
lZ1Q5lPffL5tmQt2bzKXIdN+lwJnJEvUsvvgQkIZTOktbEvZ5uMFHIMqM6QsxIgv
ge0vXQk8Fv+oM0nEP8jOw+tT/imT6AilFMkcuA7ssW6J9VhlN68r7Mu50VWYaTWK
6S7mslmahe7qKd2MuyJQ+1S3hOeuh7HJZcu/62nF9o+aPGdfvl8xbz76wgm7njrW
gU5g7n1sxBrlOph4J6EZ2Jnk6StyIY2QIZm0DJ8jCfmcjAzA98PO2RzmUaSs/9Qb
M+Q7+MiCPHxji1w9B2HGr6Yn35xcwm3pVLlnpUTrhiKiddfiO+gX4sw3xaWA2izU
X1bK8EA+dSye8+kIOMKTNibcEpBwjlJKT2Js95FuGCdm5M9VJqR4im/I/1OoMHY5
407elKFXJHFEcLYIRhmGJdgMYZPWHDEn3/pn+zUjBP+a99KKaAm41n60YaMLKWuh
o2vdh/9IG4XZVZaEHUlLHudyBB8AwK3st41HgSCTVHBjyJ2kdraLphuKRTof7eYV
iyi9ESEN47ULn8jr9mkZRwpq8SOLT8Y1laaAoD+V5oBD5Nm/KdY1Gjm1ZF+23lzV
r6Nh5CMnShToH770zzVIRx/9UIHUQlGZ277F8bZVCpDLuDJFrl9XHzJ+9qqaoBYJ
qWtCH0yzU0/DAYOLyPz03A7kkFKjvfMkDBtyE8pPK/bbfbX3PN16mogo1KgIwGdi
NPdC1NCHVb+CGM+Yq8AhePPr/ecrphhZeFlm7dpJyc/AfYfkhbl8xca6MTq76mgv
ExqKiNOEbLhkeUOMgs3a6eiIL5k8VxDX/x4nWvFAP1XfoSmwbtJcRZPibwpVnojG
DIfMkhpbhtrPvF/BViyEalwx+5l/4L+R8NTlpLn8hWzoh3Nel11mitB/W+6Ujw8f
LmdfMFUcqWrPfNAenL6G5h+0mJBs4jhPGJqPEa9KHn6wrFqDDCe4GJ5rS14CD23D
R3UGeccHY5ovAa/iER0B+S3VT9XyqJmndEfx0zujvAOKm0Tx1+7Q56LvBj0tO4zo
8HQsct9na8hLbYL9yAIVsGU7j4ZEslCUNm+tCFtq7TaV7Iw2QO7ZIjnAY2EO4Y2Q
vu05rQ9u7fVGdbM9gYFFaJEzOxRZTdwEpLb+Ux5bjcfYv5bZtXaAE/8se4rtyh3t
Qp3l3otNSkjk9mOHfLIAmprN7U+6RwaqT1m3S8n6hQW1dW34F/7j907z6jpvm52S
BeJo3Eo9GwEzeEOqZOhtgTe3eVhoentQAkhZDO/ABo1x9b5p3/N1ge5VtymuCSLy
aW6y0JTy8GgkadJhH7Vw9Xs9YKVkZ64Ser5pzLvC8Ob2NE+TywoPprCC1IXKusoi
0+RYA+sJjPxIZMZnHyemtNRo3z3sTJ0M1GxlhyGWFFuvjbJx4ANWBQ8I1bTjz1Fr
ckRz38HNfAUxrsPbYpEhlI2oua+gwFuikQzJqg1b0rbhoyPTWfsSuDlDBpgRl7CV
/HEEtP+TAlCT3fjKXVzcpnVy7Uuq6TGSgREYEZRbhzSEdIWWBgnc0JWxEjKp6Z2a
tKImHMpgXO7TnL6SrB3/s3iL7NWiIz7rX3kTpzQeR+FTOpUlrdfoCGX9UaSyka/K
h6iIj3IX5tqfO7lRevIfkh6UyzTW0WMFhx4vYpcBIv41iPr1hP8Gyh31xYHSAyV5
gg4Qob0ET/rx41aPcJJuXbIfkQeFdhjgUC3muTgC89tZTNj5DK0n/2WKlcBehvcj
hbYOboVEH5bRGEMNQCtf+oBXjJLwy/coLX/7VgrlJQ4LqrsP4zcEUaVq0oJxeZ5+
hpeERT9MTAK585vL7I+To3xASY5OJX9AlGnxhR7uhg7J7KmpLLwaQSxaNM0Yj5Hw
yRHOoUvxhQvLo07U+TCfQUvuo8svo2k4E5sY5LjzmZJ2BGkXVaFVCLxdnfFfTB7I
sOUVu04tiqUMF1JT/I5qTMvE0EKgBqZTdCHdO04FbMbCYErz5oiLyccRpfTzgmQd
QmbGAi/w/isbAtZkUEHTh+OH8v0tg0lNRNRGbdxwOD888UuYnONl2P8Ot6LCjnnh
EDUwWJJRXFiaUPNtp8OiUR9hhkdV3SrOo8HqZ33c+90fl896qSVjf24QYBQkTtlk
ZIIbf3aEy6Za8DZVN+7tu9s05iHCZFkecZkPlWG5htYVkjweU1EnMWlDjthBIhUh
8aLif4Hh5gbHyJCJvlSmz3jS2nviPLu+xJXC6hQoFlDjZc8ElmEEwuBnE3OiK0i2
kEITGNJv4c+5022TkvMYwoezjSOmiphMty2o2h0hYQnqJXTt7tAT7fSlzeg+ZvoG
v/BDGxcoPRcF+cxC5lS5yW30fzOckzPfSbq5NayhUoyW0uU+HRHY5zFwNrBueMTs
88d3nK9xBEPNMxxt77zFT3pzCGK6Z936t+91RV5TgjgplxrmfG6tCjo/ejkSfgHt
bKtJ1VClwQvbo3oCst3KIMtNIh+VxiFRyrSLCzfGaHOmZ2Ps1iWcJ+D6ccRtbzQS
QPulwB2fjwn22hMujKW8Je1Yx/TC4Z7vT/FTkFFXNrTDFdfoqFeNNhJpx3HlJfup
OJ6rxSCWujtptNRMs7QzpExLmxyXFeAd00s+8cQr8lv+mFTyKSHxcwE9Iuz5WZy9
NTbDZWavfI8oebU2SBfnPFg85+QJwJjTATpUrYA2jGvwi2vku9U3QVgrOcITpAj9
W7NFqGnHYh/p1xHjjpWcsD/jqMiO47eClMDU4BdX1YBl5BqSSjF/gAx7SLYAWVdm
boSfoGIY58dGctauH4jrNoxFP4tMgTLi1j27gWEZzpE9qEmV3WKBIWeas/6jme6B
Na5ATgT3x3wo+clbozAklvvpHu3VuUjRicmhfY6NwD9uQCUm/XSlrZahoywF2q5P
gBAYAb0IU7MOcT/rowipLhdMab8tbopiGqZjs1jSffDBdS5+exzMhwT9wMlB3Tmj
5wV4bJNdPU1sTGpVZ6VdadI18Ri3rZWae5R1NK4TnSHVooS4Q4RBpIoM5cHjy1Sr
fbtS1NVhCY8oc/DSx//oEgnk6fSwTrKWRDmaIzcfVq3ZjTe0JdDx8LkoexLtmwYj
jVvOMhLlDA3trACCkime2Z7DaZ7b2RdDuP3crNn1aZ3EIlBlR3FBaOKwOIjKpUtc
vWLH0WNO9OgVO7L0NOZ27WJ5mys7dIDgaY5J/njnTAmir6AvSjEjpZCE99SWusht
ZwF/+qvwvMt+TXkkDVbEh3FliqLnUJyGqCG5GUmff3iHnQqAT5n42aiI3W9oau5f
OupVkaz82vEojkoJ5mcsDDmaJaPX/B4AjcYmNtKOFVi53wcxQC9tzaCRYFI2bJu0
J6v5d0npCA/ICj2IlV8lpA0ZXGOebVX9eRbXl+d5KgqahlrSo/FT1/MJeEDN9Xms
ztKDeXQPbNGU7rLVEqMVm59JBVp6Ty25ps8MXSUqKcIfsreOApiOb81AU0oxqKLf
6t4Maly4Ijo50dQaJ1OxuMJb7zaSAow5kIVoNb6dcIoTom+1qoTsrn4inIg1bZvI
XqVeLdG8HxOHIn6Pj/Q15nyPpxEUV2XgeUh/p0zavvteFQArE8GKcilRPpZrf8aq
WdRm511eAxsaw/TjJCU8+dwzoKwIrbkYTj3RR0mAkYvwFt5aLZ1JCd8iCQr93ErT
QIkfBAaQEJjELhxzmc26wX3bxWIpJGyEbKbEBI+CYzwrnutSfNMcNPle5BAE9P3E
uMWVbEC8bWq1WBq3rwf9CXUv+o59uoVkw68EvKw7d7jTVvSPFPdYnosSTHfmpU+v
cvPeD8EqjS9dXVNVWEo1B66qywlgITbYoLtMTFn3OrOGjbY+OPmCjYRzT1LqISHk
mmA27zfbm/wdZvmSxsuLZmW80hRoECNmaWcu7Yt5YxZfPh/zHbww1vMkq8vRlV/H
cymEM66zKSD3C5Hs4eCbo8B9EP26TItlwOMU6jOV6Xp+oqM1IGygGYpZ8zVkWE47
kXMw3FsgSWadcRXHFu1ZSx2s9twE34mouJKdzBbDaU+FjkRaiHGC52inGc+siAqC
sqysrTa3qZBeSCUN6muVWwVGSDksBMfFjfK1qU3jSp2mxsNXcqouD0izluj2S+L1
WeQjegHFfoP2xekBY4AcHKVFQ3jipow4ZdjAqvHwifjFgpOcl/PpNqe4EuTFcc+/
EQ1rYNynbxNjQYP0NH9FILZUJgs3Gey/hodLg6PqI+mpCzeb2WXA1CEq1uWH6pdV
pLx7VuC5d5dV8HvRLqb0w0RvxbgPd1hsibVOkBOVNMMILSku7NrYCavm8uJ56QeT
azbAZuPsf5VTI9EYZm3EpkVlg3JSEGVpgDRgiiXPnrJ983na4Dm8wcnGMh0GLrdB
1Mkd1HDRpYIrbhBTIz2Q9XwdWrCGrEp22QV838okQvpIBu0FplURl/mspfLuwAmf
2+OvjIpAlo/dlL/Tj9A8w65mKZOMyREgXmz5Yo96EtxACUYuVMuY4sE8+fe+EUxA
LWG56C6s+13pzoh/TSXgGlPRSZzrvXSLn77tYv9YOiYUPJUAc1iVEpQd6yc2GhAE
csgp+iXdSJb3gH4S77b42LHw8JVAdSDvM6iBzWJUGTa8xdJ+wcTPNsOo3bVzT+eY
IlduBxU306WP8i2qTGkmpNseh7pcrE2grZ93ESai/95hsgT4Pn2U8b5BWsM0O+2n
1S7nQjUnWSJHJZh70RAxBj+GVYb5AQ1pAFDOP3bJVVaeAOMjzmxVC0vXG2t6LxnF
D/o1hHut5w3mus8ClRgSWCE2wmZosnPFUzQiEA5CBlouxA/XHQpzGZSgazZuu0dX
FyyJL+ZXhsouMZNtFw3CWPY8uEX4ugI6CVtM+j5A393M3qrAhqGi3zTFtBPFKQWD
8i8sQrbgKWKr5eyzMcguLAP4D7nw+Bso6ziI8zM0l1fDBR/MszH+RStFBr/7D0Vu
UUnIJcICHT16kdjwIkquK6ICSdNzZmNtubhVNgVsLqugUofTPCZeXKgJ2EEetTIj
6NnkJWQ9GOWUOjyTeX12W7flnKVTr5UbQgpl9uMJG/1FmsH7uY6S7tLgg+sboi54
J6cfpyQjlgPKQwMJU5Ro7cjsoqYsGFfVW7rPkqRjxIEnIJzil1c/a6PuQoLKv5qS
K1nJKVD9kkR+Nj1YmG08Nk9ZWq3kKKBCclGBBcyiMB13NG30i6cxlwMZDdzHfxvb
aFejZkER4EltgC2sba4ryR66hzGWqNghuI2Q22LdJdb4BC6gVVe+GS/eD6M7WZQu
W9IQdbxSFDH0+TBNN09HUT16ChoBP1G+XXrVjeDuGsQ7cMz0exbbITaL88HlLLMT
rw8ENruWCpDr/w/xIGNoyqTZTx/Nlv+dTEDGLXnel3QiD04CJzzK3jSnyHWC5Lsz
1fAWa/OZEoLU3aEnEO4+c+b/MndJLOdxDYgQeIf0a1xHkTl9Uq0YTWigNGXyPC45
WKIhRwigTiv2WcVHbPUgwggCDWCcU0D1ovoUHv9mf71LjF6NEPZo4AyVJdot29FR
YuHPnoh6hIVwhrmo9HlpEEShNJdTXWASjlQEr/UHXTuo4uUZWQ67S+DnQJ79l1cr
jSsN6rXwSyXsmIGWESjmq6eHKXGE8R2keXD0drGLoxIiTx6WRbB+ddw8fqSCk4EP
Tlf0CSkOY2j1PkNURSSuBQaHRMDPZQi1IGXRe1ZL0DPwPL9DXBtMZ1f4rO7zgmuz
Cz7469jUCw4HLtDP8kSYiqoSV8iN7Z2sZAwmjZyYTUnlLDibQo0M27Fcr7jgWcNI
pzjZ0ndN6E9IObRvwF7wvZO6MvIfhqacgeh4Pm20OoBoJ9pPPR0oaQeMZ2x4HC9r
5wsfh4kYZsPIWiXHtFId1QcWsFfYPiA1kwGNi+kct5SmSjLjjQmSGVWAvv7WqUqa
1gDGBtgovKS2rO1TbhwtfBv4n6IUzEK0sLSNjiCqrE7avuLl2PnWqRU+lz8QsJGL
V774koD2SKiytmJDIAciRGZkfnKtsWNjf5dzQR0UUQj3r3nJdEfQ4IJwUMuWTdfY
xPYB5lPcjgTU9erqBQEzd3chBzlQxdEm8+USYzY4OGYlqVHTY6sL/RN6c1I/+AqO
woJ1IZJo6QSpxqOBvrj4cKUrISomAQ4wgqRx6R579VM9T3WMR+z5V1ovKW0V7MDo
9aLJzuDy4CQewFqCB+hDQEyNSLBTsTOrbZolJbNQDpuyAqMy+1V1MzFsrV5F4Ek/
Dfh2Qo7hSUYupGgaQz9QlUOSsBFMbQ2apbF89V2ZDKuGMp8dxndKGdu6LRexIQIF
JtnsBwgnCqGgKTH1nvA2BJmhCpAzQAGHxcDJ3BtnVkMFAHIw00KuluXebBG7QsdA
XKV5NqqJGTg9b3lkbRxAh5boUz0d055azuGmT12ZggUKyDIxIoven3n5n/C/j4I9
0rdOI5Dpzi/hxpR9K0tpeYJoG/hrWOdyQJPYAy8hRpLFsFGUfCNURedvP+ZxZnW5
wrCbrkXkZg8ndrri8SjaU8NuPMLf/3ZFYbtGBHnJ/XHeHPuOaCHNt7Cc5Rfk9Bpe
6SjoPAtu/+M4Y4yLaivAkOD5bIs3fnpmZXlAkGMYRgMKgmtl6mJ0OQFkpBR7ALcv
74msKZOaihoLj3/pvNeE46MwWhNLTREYmMydxFlctj7/VlJaelZ37ogq7ZyO7Qqu
rv+N5JI6q7dz4wMlBWjsTmdVqbgJuL2bgGbV+iOSfPH/oqwuZmHerz2IFkIRYhpg
iNElljnAYnnrbXMdXpn+0wGFc/9FbK6OPtdtSDCqA0gbvuA7Y/CJotHc4+zwnsWm
4lyw7F3FrbnMOHfYUyFOJDWQdI/y074NzIjPO6N9JQ0KU2rpTqfT1eiw2UlRJMEB
xHg06xCgl1JF8DQhLdbRSgDr42nwPDubdnmXUVyZJIQ2ZaQ2ueVQ5aaklGQW9MZF
0wyu0nFFsQ39oOu1veWWx6zq5QPPpFJMIzlxiGNiOTX6WKDlrG+0hca8r0Ir1PWR
IsOgdEkQ2ncOP16Dg5UqdyF1UYu1SmXnBJ05DVh0Dc7DT+A38vX//C25oFuSHcWq
vhnOuB6Au2XiFnAvIQz1LuTRqNr1ZWCmRtsEybMun66JsFv3N30X/XZ1G1Da5w73
TKveJHK16gJKyOsmRZUa0LfWDpJUJaXBNUWyEvYH6XN0v8Nalba+/7go6SiACsYC
60lUgoj9A2eQBKTWjWMz9KLW27ZPDM8meM5FaKrioUFzPMNS/mQaXzaoi47XFdMS
OmnEMWe9d3WgjcsWziq+r1zHUXjiMfmWAzpG4szUUzQM+/Ts9YklSwwthf6p8XbV
Ybx/yQpbNQ/Z4VM95mp8O2UJRs/fxfkbK1IPSwbh1k4RiN/PPRRQyJ0cDpMtjzk3
QMgcPb8o9L2YqQUiYV1zqKDBhY0qSyh930YrtKpDtR//oFScBH/jbwu8GJdXhDPr
zMmxVFrXXPdeVdIswPWW3TurF/p+svPMpkOcmhskuSOlXtJB4/p+P/vF+ZpkL8ny
KAMZvF6tUYCM7dg3ZCDbrGS4L9rBR1/Dhk6/UfWTkyp1WMax5b14gx41Shwy1nRC
HJBcD3pqd+LiXTZb6bpWlXlnBekPUwBfmsEEqufWzUCv2Lw2QQh6Luf3CgcT4K8P
2sAHm6jHlaA32v5ZR1qUWiE77DhoZowIF+G7x8E8xr6Yz/HxCMWOv1giVEp9ylC1
N98NQQFSgqr8v2Qty3RLGbnKtwGeIh2b/P2nvsC1RsQUFH0RrAZXTBot+5buWKh1
JYQib39RyHEX2eTkAKOOVBhyLI4/d35+lOOlRi1TDwb45wtupTY7x0zqvgZqtPy9
AHt5/TaTosjl6EtDfrafvmD8sfnykTejNxCf5bSGDfLwAFDr+tpWrDQK47xv1jAg
VdGx7E/S8HELNRMHWN90I9cwKS4zd/f1B/ffKy0SShBY2gcwSnLLzFFUrAAJswXg
rdwhI/hM2UXLYMgZ0EP08J+DDuxaDTvvS61wsEU608nDzbOr3UxbGhdxazBbbj4g
A3HB0eC9ZDOEpZ+ANxy/tKoK7J7JqGd+Sh0q7pLg2+RLG6osVKUpSG6B0FcdbixZ
q/n6zpncywoBNlVll03NtG6UuQExzHXYxxzmYSV9SWtiqO+ztIpWjvO7o1qlZxyl
MZivpdJYOH6dot17vxwP+zwMEQGZ3nUTWNb6xuJExnisiO9ntI3jSAESP3n+WHhT
NOst5R7QBbe1On432SU+On0P95ZBS4FV3m1N0W9RbFfmPAo/QcKWcCS+AQaVEzDi
olrAosfKZGHhHR7NIA8rPeUsMqWnstlnpwjm7KO5Ygtjnwde57JOUrNNUgHnPM4O
EofVfly8ueq+pAO5Lg3tTheJ3jjUwlAWqpiGSk4LBFNNKpRRR9K6fp1ucu8dljoM
TBhMRjaeTTtXD07vduFE/tz6LPcmtm3RT+bnClKAY0i+gQjUeCaBULfz4/g4+IiE
6NOaH+mBcWGYwWcmyd+Yp3UhFpIpMKfpgJnbCHeziwRFX/3ubTj/Ka1VRVSzZ+EW
SNFA/MkQ7okzo3S6NlLT6KN0iG0zYd7CRdxxwSiheI6hU5BjCYRCcqH4/7crLDzd
KpOfLbcujvRxFfqzL+SihES6F6tIj6IBpyXNabvIwLlufxoFGNpuoycm3Phxj0RB
uQTffKL33C3SBvN9RmjVFxI2RPBP5mtpah5JvcWmfx34Qe+a5zjiaZAdI0yvYZye
Q19Y1s9dA6zhbsgrDqK2coxcyWB+UqUzCdiV+KmiJF497cWQddZ0QPcvfmnYfqdo
OyLWkYszlgMzbWNv1YuPZ6DxycevjnZSc23tXq6qk8E1pHXAmqkubsz2pcrEI1IT
weVPjhWuKQjVF3xv9Bb322qvo97rkr8VIItNNSbORbzCXGwqHRxE/B3XcEi487LF
o0b31KRfwBdiOqiKul2ItoEeGkN8vPzyS6nhbDXW5vM+vxgyhUSMCKk2/vWjJjL0
fApx1bC1h/ED1e2ESFThJkCvDRpwijszG4jUoAk4fmh0K50Mg+rJzKaWOHYzlmJA
hOrg0ZhwgQd5LVBbs7fJ1wS47fU/Q+tnPcNT3wiCyF8CKpUVKqiB3EN1tUR03qxo
xrTRsy06tZ5lBGhnInGudR9BASMj0UMyppv6AMDcO8ofzIPJfwhVGAUYDp9h/p/E
Wbep5AkwLrnMBvenx72bxlqjBqjaVbVPyiUm9vxcgQmrFWCLcSidcvFuVJtY8GsK
84bYEmx+96z5Eo5xnC8jJbdw1mu/loCFPKOtveW+eZlvMbc6sdeZMbsEK+oEa+Bk
FGFwm6UPUaX28f/MdEgW2YnMG7Grg6/YumC7uC0RliLRPK/6VTbszSiChpZUIAlE
YQ5/YIXJzVmaZoXL0on8CvBruu3BODDt75wZ5bkceqjEbLZH+6q1ppNA3++jcH1T
uDNXF2DKxyv/djDW7LHs9IP+dLkOitgGCkeqlRV0PJzWozjL6ssvJfScXnK27LPo
anJ4JyaQXvFd53b6zcdAvlBKQchv8XsKUQ9KtmHeGEFPyhZZH4AZdJWxkM4uGKVM
NYrdn7nRhaF4YmC0LRyA0l02z6FBeR6FBbhQs8GZGtWDTxcAqiS7fZZ6TtT4zFtQ
u94B+tuBwMn/+QNgOjwocvwQB5QcVO/04e92+CdnLXSRUTViOaaswEnqJbvX+fnc
uijBjIKBQJJsp07XkhoZ602HrGPHt9pbgDDLBlROgV4/2aTAD9SIhmUe58Nu82h/
SWsb4oQJ/Rk8HKMdO0nfescRZlqagFIuAeICU6ikB7YAkROlwl8QteKSgQvhsZf5
QtX2JCtkk317foP1K6AmigB2Xv3bHPnJtpj4B8qMexra2v2gm0QFFZzUg3V7/FTz
GEg2k1xHXu2gSINyKC0/R2edutTZa4flvSpGYBNtve5dHcKTHRrv3gtmgGanEPAk
okpvZNmaPSQ8x0qngrXxPTq0balWlfmsppxmtyaLlmf54sFfx/iJj9yDRYkS7LL5
+4K0DLxGcTTKnqQHOW8ZgZb4zX9NA2O7XxoUE8Z/xL6MrLj5WcxfpIrSi9LbyESP
kwWa4F5DBCZgpxx+FO7S5Y8YzGM77OQcyEb8ATkdVEyGUNK02CcejJ9wa4Ja9plt
J3NEEpJt3/zzB5TnrPQfSZeAthuIFT/hlPZuaVKVY0K4473+BTlLXyhLRVofBmAu
6+k3Os02eBIbD3ZzS4aCXb+Fdl4/hkKTUpGJaw9A/EX/+geoab4839mvtr4LOJeH
vUSuXYqNDu4FqUeok9GBgwF9ALArinrCdYsg4tRtAMEOeCYLaOHI01iyDhBWBX5U
T+5d9Zusvlf6l9roazQ6eleglHCGUAAYeN1GTVKNwv/uvJaDQb1jz21F/LaWo4fA
BcK6HwDC9CL5wgAcQq7ynDFatmYOHdmKLoSzT+6GrIvH16tUXVzba5ieDfLja46+
RmZwNVHQtMhg+oeLGptt0cwmBJBKy0S9eajDznR1NUOAXLCV1AXIp4rytDvUGyzO
C8fB6QODeDhleOLkBLAY9nL/i/SqSVoBpvTMJZu287JxvkSNEn/V7eEw2T8k2tK/
LcXNAN7dCQ73SR5dmwYKIK79RE0ujkGiA+O9ijy2jeqsI9DbInSnw2OD6ZZO7bbW
DVb3cGL8AAEN+DaxBNtIzMTZhHRq+UTzwde/9vkaC/fkFJU8lc9BvMJBtGAG4qOM
N3Bu79tPJ3yrNFneIl9gDWlDaaixRf6HNTfi3+UqsiHk+5lZvIIsIS5CefV1uy2F
4RtiV2xdX8aSl3fE7KnWZ5RYIz4CALO56qAHM6CjMV3wJgp+Zs6M0DMf/Q/EmZ7V
yj74+Pdd85uA66pHSQj7jvGFGQaX0NC9ay4mPVgD3hTREPo/0K5vOoSf4EvbvDAs
JFugSMRls1zy6qMVgcwLOrdt31at6YPf2u9PXUQdRwX8kPlyCOJPj5eGhCAUq3uL
DFG4Sj0nZECejzPm6bKfNsOwjCMN6MtIOcG8sjCaQN9c/WnC228kJ4J66pjcmwGB
5mJwKThLO1a/2OU8UnmWepz1Iql65JyHAo8MZssZzvqGA7QdcvHfOK9xWwJ01v+y
AfAGvpA5PNmWcHdPt1VqBIwQjZmgVUCni09ibfMLmmZIiVdRYfhibCUbbDoHSsd+
7yOLab3cfkBhPrG2GVVdehOyJUB3VzQ4mQAmklWhFC1tG3cibPSMP7VsNzrlaeBB
Eay+WnWD//tSalknY7JxYSVUs1vjMN/FEi7/TOBE9m5HrDN2VZMgQnbL2OwaRrgA
JZXv+v0r0u7XNGJLNLr6tticXPYATNAszEmKQa9P6YY3tPmkQEKaw+UCvUfz+qOJ
fJY6XHV1d4MnOPe1C0XipaJhdZ86pwFjXJyyUwpsnuCY3HOBBLfxT+zixBMvT2eL
opUae6Ppqt9e1V8hNQZDorrVuGitdoyFRQPiIEqtaxupVgO9s0FkpZDbPkiDBesQ
PC59czBRVqmPHw8Z/skfuJzPhSQZc/QuvTfc5yYFf/U0qVgNFpG2IriI9TWfiuwz
Faa/02FHDwlrVEzyrEQbmT27RIE4t3X7993jH9TMDAzuEBh2KAJ+YYyXbwlF8gLR
d6eVsFHfTBJ/S0tLrrTgFUxBNtYg5B2k1QI3bD5dhZtTT471oWcT/CUqnhxu9LR9
Em+15LMwPp5GI+6tMshN0OGM1k8CGxgsbVZINNeI2MixmFM/3TogB6uD0HQg1J6/
Y5JBjPpd9csP1Pmd9Tmx7wITP9wszsGkmEOp67ELC6k8+hgRm7MDqsnTmzqIUTeJ
/8oF94Ge/if60ankCwS/xrWyI6QBZB4rn1HmA19Beq4NhrTgVnBgbku3r4jO5cFf
xqWjbdaG5wjSsAMhw44BO77E6CjieNy0OvJ4vhLhK/uGYf5ygp4sa5IBPJaw9qEI
QoR3k46RiqSQKF9LJ29+wGwuEc2T9nezhzRCQWuWlZY18AtJfPRqu/AwNyE+NxNQ
JqFs5nQSsrhD2xS6WPEgneBr/m8evmeYQ02FN7dhgos93u/jKSi2J6q3xb5ExuG+
PGfp6HJO03yz5oEW0hsYsvQir8VEINACZQqt0pvszGcCBq1/Dt1ZvdZbe/aso9lU
2ofbi3E+TGLfbh7ZER4W+brbLnkWrO5ipUUPw6nP087kPGSP9+NS/ImwAF+U7JIH
b/Py8F9d4CPlKFxUGaHT1vzYLcBhMK3/X1BHnXw1DkdOJZ3fHXA5WE2LZyN30sGK
FLYAGV6GZKHxTLl+kY2+Kyz/2GCbn/v0JV6pAgyeshqliXmIRRLRlzKaqNXaiABH
cWu0jASft3v2N80D1cLbcxpOT2rsp2pTOy9DWIUDfBIHxuEFJ10XAJiz/skvagja
Cp+BLbfnH1hfMePYZIokUCDAdNDdBgI5dSxizkh7s/SQHe5epRranppy2kcuL9mJ
0ZZA152mwNzEBjn3eLWklaDwHD0NsZLHoqTw7tugvc7wFKKzXLz+v0eo2EA4qLzD
o/qBRIo0PDnzHkPA4tbNFE2h6EriozMjU0bkCbYrCZj9G+AeiSBayWQByxz130le
WWCMSPUX47UUL9VVddKeqw6gUIh5aDzEXS4ArG8LcvF/li2ukDVIxZKaTlfARwat
sHrBeyFFfIvhDD6SabWt/Q5YOQxI1p8UFFQ60o0BJ/mKHkHUMNuzFaPBBmU/jD5L
VP1pANieha+McOebxSdd9/DBjB6sNtmmgIwQH7S8LmRtfaYh8EdRtEEI2pLS10jO
Dot9sSn4evxIKyh+Wb4vMgn1FZaPXjNJPnaGbk2xUu1aVYHYCN9yfhOvUfhIBwXU
Vgfs9upq59lp9G8Jed1XHGxjl4xvgUo857jXDkEoGbmc7qhzudCQOFHgcFiiW4Sq
M5kVJxO8+tbhjDDUEW6zqn3dFpqyqvOLzq5ITRO+JLTDlgTRW2ypFT1TG0Lgdyuu
19sNpDZ8k63+0fGOEQ/qvwm4PYgNYi+UV9yTdisCIWmvD68qSSImF6Ko6x8FqLTw
/kPfdtSBLSU9oegh9/QwilGIGpBqAxV+Dz7qwVDyVO72NIYXYKuyyRPkSfMk+2+N
DxdBPUiO6cqEtYp9MvDZ3wFSqROYYo9KHm9yy3pgfGHr3tfokmSgMXGJA0HXX6pW
ygxkhEMcTW5KXbYSj8XVhKKgzPNdyNITV4N+872GG6Ly7a+30CmU1+ccig2YmJ8R
75RTfGM4lhUlEc6csbgr/FddP35MI6iUuNBkOemp9lCAnvbNDCCQUs1Lsrq+rlFQ
oGV069CyBkKYbz/7gnb3FWAHM1LOoza6tRmZw+5Oon00/E0DgBRr+mBUZvGWAI1K
NGhiHtHStCb2m9hkKXdk0l8cXD85d4qq9HEFN0DH5ZKhD0z/yZAQCaCnOvRdxlCF
pc50nl6ga+aedIx1zYvjusVkb6P6tVAVuGB4ML12qacO/HdqwNESsSU5FdCu5bFV
Fkt9fUif6z7Niewctpi8AZICtCdirVhOcyoqxJ8Qc0XLv42uHt77B52XUbBkQ6pL
iG2Wf0qxtDcYdRWsmrVEU26EXA33Zof8BVcmgnFTFLAUFFcwW53iNbn3YsIOrPF4
uHeF93beSYub/KAeeM9Sw7ABxssnR2KhHBhU164ym+26zPyFHe9T+k4L3Ne5Xz0T
E84dVJqXXBkYOA3+pwFtchx5t0oNHinkJv+I75TCf9vb6wbRj11NnR6JfcKjmtv8
AMbQG8bZHIgKN/C43G1RD7aYWwkXWqjiOvWxRPsfXAPpU4fMon9uXHlacq2tDZLE
7YxRPx5VuxbyZdC/6hzQF4WocEmdbgDLCDDNapLGLFJAwuQQfRBVCkYR3nVwoG56
KMTGTGGSfMwqSE5ivkuK9seHDFYAUQ0MSqQQaRTgNXEgJLjHpNmy6I+v5868PvwT
Q64m4a6Oe3XqAIXbw1oLZv9GhU0Ge1b/6R4qoUofRORw4IyPJv9g6pTMb4MEMtbZ
xrdJECPFWYQbLHPKUSXG7aiWIX9IxoUmH9qFMU7gB9qjkD4SHI1G2TMLIZIX6FcV
HNpuJylcZWOk0SG9z1RWiU6R8X309RpGuHYiDIeKK3jJODcz8SjZwOGTwRb0vuDX
8bzmheLtGlIDOrs7jEiIucbHRoEJG7H/omoJyk3KYnJaYwJ5GgMuSa6E+wyStsuq
8I6hPMli8NfVyU9M5yI4XvY6LTUzmFPQWZLZrCH7hf12jO+0IxIZHcCmOfdOAhCA
3aeVHrHbBIzUhSinid1XvDLnQeN49mQ5dzBbAsWo5cXegn0jUPYvMJKCjGhoA3rZ
P8wj+rVUSN8ERNMpYZqgWfplkZirA/lhYkQjgu+FZllDwR8EhVyCV6wcCAn0U5KH
/OluatejOH+uBeJmO9ZE893fRQfnbtJ1OFeyloivP6MKrJ3OteFDWW8+kviyEcKM
T7HHINi5K2pn2ZSyIHJin4XBqzSzdYGYncA2bVBMi5zzCzCC5A0HrJ3oAIJfJMlt
Itin8DlcpcXw905fXD+O99vH/waZ0MMCnBGUQk8wWqJCnScnSdLBv792NuXkoZLJ
lvhQKqRCI21PWM3Ehy1Q75iK02I3/RWbRSNZcEhBxrhArxQSBXA2ww7l/VPz/+0e
tCfldgtbB+bD5peuxt2SxivMOM7VNL77zJx4yggCpvkjoSEoVGc0/WgV5Er2squa
KSt7cdiAwkpPn5+YxCRW1PW+v6rM6YuxT5bw9wQlQ9uaVI90A80U3JfiKRP/h9nA
WUtUZ6mc0SR6WHHuHXIe1Xs+CyQ+jtH1/7ZmYvEugS+HHfnNzOjSzD5bAcMVVJb4
hpnIKavW/2fvXFbCto9Mgwb3q3MvAgMTqVVMe6LxbezF46zNLrLT9yPwmmj6nbNj
n8cKvYPQFy7T59+TOQ6VBrqteUozwqDPHhV09X/+X3Ivg4JDdcwYT1Otkr8rf3ZX
TbK1+LtMwN1p7YwqsImXBKUkoTtmaDVuf9PsA8eiJ/pitAEgDGr5V7kSZUEjJ2UI
YYHeBSZW+TAfVWe1pwW5JdnQq7onePHKRgHIrC3IwhIXpZC+dEL3KO3xtgkxmvsP
nGpd6biOHqUGFNMbUayxBeUJrR4UVbXLoG7j5S9LycvSZ7dv7A+FaXH3Wf6Yx2XU
3HP12wpsougZvJqbSq/5XI99j917gauK5380766sutRcSkFwpPMUTuixnO7brj16
jcJKGVko2hSkYyZrHZQHN4WNoNRvz97gC5bfeBuDKKSOeFuvuMz7liDpeg7Wdlhn
exiNpKDxd1zPk5kNoNE+qh4N6Uoy6DbpBkvualGG7qM26AoXumes/68+DqP07gn7
FDpMFYkEp9LcWYMR/f4b8yDYy3PPkVxr/ZROO2nwDCA/rfxocUMr3O8vmfqS51m6
8opOnSci/bxaHAceNQpaf+FAtHIEN8A5fx98VXSgQvwV1fFuSVc3fsXp2n0gZxD4
SrQyZ03jbY8q2djVmbWW3zkwzXCyoWSgkNk3Y8Keby87J/oZrOeqwqJY6jD73roB
lw92qdhRaFNmKFwnI+4Cpi14e4mk9huKGbMz+dtqs/1PdcI3xamSllZ18YN0oJyU
90TJZRZmLb0+rmEYYS9GjygOTPm7bfTUqbzNDVWV0nOcnV1THuenW5b5MIvkb0QB
2CZWlP66J5omIxB9Ppv9uQiBH6o+1XV70weEcktlXqMaqAYl7kLd3hHXgtQWTJB7
mjV8ZWGHhHaZOSHGKKLDP7D06+QCMYVbSkplPfwlUygUJmfWVtrGIwcmcWji6tlr
ciKlnj0GaABiX9cPOnI0apdAbbiTwowd7ITWEI4A34Z9EyAWmUWojpFgY+pdpC0g
2A/E6VnJsXIzTbhAEfTpB35trfLiLrR07GYecrtGDBj5FWdSYHluprH13JXJALIf
UOP+UpZ5tpbfWPo283FzFws5E6JiZs3FyRhRFFDWbgqeizraO2vScW2/c2YxKqP8
zd5Bwxd6S6KJmct7M4s9Vn56cbBUljYGhk+Ods4JTQMRTow9htqkTbxMHxSOGeKH
VMyg2QPlwt3dM255Fuy55xl0jOdIaANUFaLX2z5PEtPn162drzv71KqhUKrBCZJL
vZzZNdLbSZkzqf/9SeIgLZaRxQ5hNSttiRDNbZRgZ7UmfyhAcxGmvmQiTAn20hkR
qOpW8EiimtQPbuMr2ZIf/hozmIQxDi5V4es+vwA+jchWH227ApihLu384jCMh2dl
mCUTf/ofGMb10p4fu23I4aQQhJ0E5mgak/3so/SXv1vcroL9AV+c6Xm+EE5b+2/Q
CtSiXkznKF0mhx4Smv+LIxP1V8DysPzt0t1FuvfeMIjI9vwP8kZELWpLxPJ8Ep3q
gTfyIlGsxjYLO5DZZdRUicETH89Tr/I7ImlpsvA/ua1eKZ0kcanP/qftbTurXycQ
xP7C8sR67CLcydBYnuKFcb86nfBWbPpZ8v9XaLg+wqsSuXUJq+h2X+79v4PnCjAB
J0yqFirrbM5rDm0GlpgteHos6wnWGTUiqOuupXWp4fuWXVsZSdX2VZnj/IsfTADm
gxCO+UXrz7LsAXpIMXfl8mRzqYzXXOIhsipJ+x5vp7CFPQsBEHZBQwY/BFr/YSjq
J41hfoI/Jrhe2Fn8HGYTdDLBtgMsNBvz9eGeE5V6+/RdFcihG1u66OYkV/VPRX62
i26GiuXt2XQlwgP8Paexxs9yBuesqwa7KWRY4sN7ef6t3vQh2dGEM5paZNjCoAtv
s38OZ1MFaswp3CC+KGxTax4JD1qJ0hml5hI6ZzIdi3rEyl46QcnMtZv+f4FeeFyP
hefSODfegWuUMoVZw5NddtEuiV82epeC8ID9dt2nSokb26GaFPh2QZPYXQ5FFLd5
eHDbbTc5EzMJ6vOWe/o6E8FgkkcjUvWRJGLL+vemrDwqnZBZ8O+9/FxUDbxP7R7q
uyaCbeZIDPG6QBUaHrj24olVstW3PKLSFkXTDSJIjI7cYJsbCAGoFSjgs+Wya43W
H3HSsOmr8w3qLk6w9BxkIIAO+41uQasBq+JztxOEBhwoB2Berm2hGZvCVTs0shs/
6IemKVQueuc2b7GW2P5ZXVP9Vq3/FoSJJUMWiN7NAkc+sYCgz52WXrnI2pkYT7OW
rRVi3lQkc3zq0e2pAtp34uH3/1T+2Ws06qAHAJrBXiC/jEojWTeqUrgDgn+rJ7sj
aHKZ/zDsrACG5N9mu6vZPBxcvp2jx7KZjXebD1l2QF9GKqgkKRkENH3kHfQVcUaG
qglKt7xRzhKyaiMvbHEsE+nGP0LdyOuBnzUcHDC0DjEyvhLotfydzDh/kNinKKHg
iJ4/xW750u2ZjICSrWyzbgP+ZzG85KhRoqXADfgSZhU4pgdr7heyMRteuIGw6OXa
RS24pEP/rQJX1UA6cwJHSUr3gTQ6UufXvN4Js9l1Sfo2MqvX2A08kaq9rF7Nv5a5
2EWnawX/DDn72tNbqofOO5d4zfarpoH0SkjifpZHfqfVjzErq+SvlKQghyvREfO2
npQwlXtCjK7TCidNDCobTXeFRuzmVl+ARm2ft974oY+ss0aH5lwIFnuSD09EB/an
fHkqIji9Ng+saBE8GaOCm3jru5mDXnudP+1Fetq3lHfKO7QBDAmxLMgPls3o7onu
Sd9Pp8GrbTZirqRnEqou4IUhfq9GOesSSmZ7LpGW9ZRXGt3En5VbaUu+S0N6BCQR
f6kqNW9bCDFrPTRmGNQU3nl0rUlpgo57sfhLHsq/ZZdfYNTmyFObrAdX1tpUaJo6
5RXbWnrjCmgla4GNCxbXsG66Tip879ZiDE3fckOOuMvzDVgt0sNCH+X8zqnerS2s
ei4qTQgTV+3yCQOhmDMi3I3X7ShHmC6lcmbmqqryPK+Q63Jf11GeivkXSUB3sm2Z
knyKzTNguoF4pmtiQTLms6hj0N6X5sRt6vQerA+ufAv3oJeG1VitclF/Jf7kAucW
IZMgh9/6f6fVZh9/yO6WBfOWSV49fUMHIeFNmGJT2sHM16itthTxP8rAWaShlSbl
C4pAuVWO5BfwJ9YMzyRky0c6yix/TGJePiRcd1bSSYicyAwsrWIHO0boP/pb3Ygn
Sj6n4UroU24sIV8UBXIk90tkjJP5v4xIWiVujy/8772s/By1WYqKwkuWKHnecvSh
WlZ0AqX3v2FeND9JekIM5TQq8HidCfkqynXnh6ztT137vSAxP6yLzQCBSOqmLvGd
+q8Z/ZFzCGY9jjdppzolEuUGvyfGGkFLa3pQpF/ksvXBXmLtHk9534l06quXmYPq
JoUClQFko85hqkXRaRrIeKx9B+I8E1+vb0uT2gdYYXO/G740OeFiOAF0vR/lyR3s
0FYwxLZnbgi2c3+NRg3jw2lSx9I61pUgQbgE/N40+8Ym7oc/IWr03nMqhpDWLcnr
AgbnqYty7FRBwycFV2GiexkkY1+9Sa21yPxY4WlF3Z84A0ls1zd+zw0KD9BHEl0s
7XQop9NXIhwgAJEnBKljf3FGRzHqPb/YlnnTf/B3AzwHtveanH3wPQfn7L159Pm1
I0/g+VhSlelOPp4WWBj0bDsR9O7aGPGE1qPuTiWhlivs4hzUKgBPG1iYu5m/teSY
ExIBJt3mp1YZdM7HZtX5ojr/v7VBEQvOWcSHyU29g6BPmACio/8S5tV1A0s7E4Vm
8kpEAFxDxF5zDrwJxuRFhdFLclD6Zt5Kv0SwdybX4267XajUPg0cg/GKddeg7lA6
Dh2LDlR5JezL3NVVPl8h+PhMRH9/O5FgGLMx+1Av6hLTEElq+eDCvwPRr8Rtybfv
cAJOFJkMIaS3JI/kc/xHvP4Iu/V08DhwN4ZAFTA9HfQ/AjAIvxA8w4DpACmwuQkh
5/uyxZLtCn9Lry4138fpQbQNrNkg6VBDQnoa9G967bvaOIicf53gCEFWVmkbWSzq
oTjrS57XotOjgvJHPwEhh1+vlSPtH9SM4NDmmOl7Igpofk8hm4uGf9XlY5ctcvFc
wkwBY+c6YB1J6xGkwYDKOqtELhphdtdfJH+M0DA2x8hy8iaETAMd6EanpJramAY4
lR+9M3LNEf3LW/P8FcnV965P5hh6J+dCFFK1UdfFrIvoeEPPgR3naMXYh0lTvwur
DSUlh/bD812d5CPqv1EQLC2+x4QhRtKFu57ZmWvYOTmGLyJzLMs5JqcwvI2dxo/m
XR0mLaRUD/JRQaDhwYtrPTijhH862UL3pjDdrjUvB6R9Ur7FTPVsYOt9kKEV6JjB
7o/TwpdPczfwlnQgtx4Kc0wZEKBi6TXP+1yWpKiN/Ofp2Z+ZUDoz4afhTnwMJGMR
cDAX+IRQNvrCENbCaHwBCjcCLYUgKoGGaHmT13e3kXNEj0VJUgIvQ2Uar7SGuqYK
wFHBQyKNQh4C0J0BxVD9LCb2ADlhahH2bIolShAriDD5U/L6Xo0HX6aELCxL0b5i
yKHcfFYgSButTQo28sAI5IYzhmM47Db3QmaDqNn+Ro8ZzVqQP5p3yBH6SGgc3fEd
Fqr9EHzkA5x9d4TpIUy163mnxEZD42Oi9wEt7HZGlkAUqoG+duED3Ctj9PceQ5Py
M2GFumX+ZXWyn++b/ec7sb7dlVTPr2yklzfghG3GphfhUh0/G7fLGDbdI8N14faZ
UUbss1Om20w1YD3bCStyahizyU0Eu31rqKGVq76IcyWM98us6G4jKVjCmisFJpjM
T/XMRx/bixfQqRM5ZnKderBY31+1pDtC9N6ZcRE/xA7El4oH60EzdT/VykhjbssK
ztB0bi4sJ7LRUQAad7arbKn+oSe9BqGB1+ItNjWQOrHyhBz52GI3plhec6SNnZcy
270XpuvQ+pvk1JcJ3FLNp1Iq4meIH1xrSmhP/Qwv46bPpABie/5d0DnuPSSZcw4z
xaIiNwT3NJTHrd3uEGW8FsDjnN5dyg5UTI/2P9Qtt/HBLBmjiFwa17t7OX15jFYv
bAeNrYhBuu+1TQEUimKSdgZ4pMCP1wS8gszsi6Jb/LXtFl99KzsC0UTUwA2XOggx
iCXZFk2IK/wsnuwUjjy87udZPfzNEVmTp8pMtIBqwrvH+BnpwtJRN8L1I1OXTZaM
BfBKXBEagtN+AAVhjIwkYeLyCPT4mHVT1CBnEbtt2bbhMB9vEj9lvg4dhs31zaho
SAySEAkM4LJ/c08atGBk62060ZKZgW285gEeXYVW1+z8ejDO6b9iypj5UoiQxLi3
xUMH/9DAM6npCi/Wndjsy1J4x8ItvGEUb4PymguKCCZZewL1/0tDGdWZkiLmKrn/
G1dpz0zDvWeEtH8N+p2WUDxw2/mI2ex3b25J/74nOQUK31BZPMbKwQu06DXOob4o
mc7ez60S/h59wc2VP6QbK5ZBC38iCStI6mXi3JVlyk+yMJwVgkO2ryNtFZiKCDFA
fgmglFx4Yq0PWpHpGtUfoZ/z3FYgnsd/Y72WtQpwnWORoi0cSdbogsAz9V2Un8Gq
561ZEKd+xf9ifTg4fqR61VUxfnveM/bbnoMgDAFYtkzVGIm63PxRic63Ul5d6CQf
SE0QybMVnnmLoVqWnbuWnYaHzuUavs6UW5MMS+zRX3FFM6xEW/8i19KtZYLO1MoQ
x37i8wQm1QXUv93SmeF0eiD30u+0X0wmhrS+/9JsBfEHguSdZDBtJK2Z+3r+5khv
FHWE+yVdnl+LguUMqvsHygMFMYqjNCgUTxIHI5XTt9abgbNfTwasAo3u8X3AC4aB
tdjQmCSOn4YWZHyhjfw+xUl1/N4eIeiFbWPZqwLE63ch46Yji/M/dZDvpvyn+zWg
Wq5DpQtCHnDKjPxcAfRk7MYNC7uv8UGFNcEzDxJAswH5CY5UDcdcJ0gphXl/JKIA
fDLB9KguQZDBJrFu/oZkK4cWzMg3m/4V3n7Z8o+f6mVpQbDAAoskPxZS0Q4rEHOZ
U+5GYXUoNFmNtetXW19xICoLZfEoQgLyJ0pizzfhrTaFWSzDrhKuySd5hR1XPjA2
w5b/L/IdHCcEbvH4ZuOXeY5Q9Zg9wUW0UfbcKg/yk8c8L51n8oMBygwjmRVBZMPa
DFwd2nvJrSF+4B0zvaleo1oYpE4CBkPRx++zC4+eduQ1JsgFqgNWdL/IJ6MY9x0V
RoYya2CaFn64XTY8XaL0IOqEJLMqOHuzmcPtdpffocyV71xgeTTSNV5wPxJ6wcPn
s4ExgweEcXGJSxmEFM1vuOJDVOhVV/Z6zBEv1mGn8Z+d/KolcrgUGsj69EoY+YDk
c3wd4Kb2Mh8otvx1NiL1myQpYtWjGzs+gbJMaCWZOR3TMNAljmZapne2AF/NozXg
9ALI2F2W/sBlLUqIIHzhKCTcbmPKcJRY/6lCraxKEcj8OmS3Kg1HitJHYX2ECnUQ
polwYcphilAwr6bHk5s0/E/TZwC7c6uBbH7dtj+1BzVZWThMontiQ4RDpzYCTx3q
DYUajFXbjjQ3iyD4HCPwFtOTm6GPwhCoBv9EEvIjynvmxb/DzhoDS9+Nd1u4df8z
A4iYZ/oveZtaULjcrcmlSZOfvXmKPvpP5kz19nYNt06aYcQu5yyQ6Z63P+M206JG
UZfmpyMW9d3U7Ck0vkS3PuxvGX/sZEHCvt9N69fVsuLNf9HyR32+ff7+lM7Ebcsj
sY11pvby/FOnORJFEQv9cMb3KRG4yxkvKVDMPUDTFI+cHorh6rOePPFSDXHPH2By
3m0pcVMd41OsYPjI5ccTUDf4xhXLYBZyz1bUt7iNSXPZLiwQPwdTbOzyaiU7g4g2
+0PbDxFfYe6hYKFsw5uVEgW/Hi/Ni1vOJ9yC+JT74zRAK/0Lq8oCdI0gdKmErIlb
kKPvhhCFR7FVda+LsDGPLyB0q48oP1BvywHwmO5NgH4C4hxl+VDm0XmbY5gjSRaZ
yR54nPe/1KIBTm+o8isk/6OdW2RqyFTIH+UdeEvnKcneR22IiVvIJamgNOa8a120
9vxBDH6P/nKlqq6qaaFRD1FfJpELvHTOlZCHBhXapL9MoIChniAPAy/dy+x0CSeG
s7I3o5eCS3NGjlGnYLWqDLQOAQxko+DvaN8iWCIc0ykkRBiVQShkCZ+F7CW55AkU
Il9FFnPewxL5M0WByPOnJots9nzrP2ZNYs3XQjUJx6ZtFn0nHZLE6kZtEVUd4y0e
oixvtL3hwDyh4E8ZH0JDO1I872uLRKKgz9Kw2YKZU6RI703gWnq+s6/bdqttZNZT
bgp8nK1BbVO+1lNC3+ihpkDxIBC8SSAb/Yu0wHOpfUkWCSy6RkeJPIO7iGdAnlKn
lSLdJ5WqSLBX1aaGyPPtcwDEBLaG4bQ4xXaYgDM1gHZwWQtRh7anXfmoh1zlxF0o
Oa3CMxSddoLPZExeiPaJ4hUzSKxXPJIZ07Hadj77szTIfmJq5VrAxCnJ1Lz4qI+8
3NWMN/S8e619QwAiJGiyW/TeZw9vMlgp2hPfflPkM/1tuGUT/aC4NKRN72i9bIgh
ETg0ToPxIrgBKwym26lFDcP/2y6CwAhg92ghU+CnMdSHquem4MFpjHCe+7mSkHMk
khgShrU+mvjZSt2uuHGGHPTKFRUfGbV0l97q9bvjDZqSU5p02k+f/x6p7v9g3JS+
wkgcYYMxWH27E9p8OZaA3LnRUc/KnC3WdCYSRHAD+7vh12nppV7NWJ6u2IdGlL/n
4WRvcMO4ryG8B8qbR7VgzKQJqilLLGNULt2QGSxbZz48peeFmDOQfbFTAFrLyF/I
1+4DsFzEt2NnkWOlP583nJlwx/WnVdIZPKgJbD+l9NrijMZ1G2+t5kgMAZDBPVLf
sX7hqTgFS25igha/dN3zoHMJ1gAzEarwdjbCvy+jKmr+ZsWT39Y4RMiaFvLzJW/y
vuw5oCkvDkhhcJzKgQf6/woBb5WpISWg4TQ5ftvjdLU+QlTtKSP/A+9rOD+SXUle
stF/4QMt1eJTk/1yvuaAGfgdYnSK90Hx6S4d+QR33OoXUa87IV1UbBIsfPb/aOHb
Yq8+Oao40tXThSyCiiP/hEqz4P/oE2kV8Fx0W4ZFWswimSruhWyxc3+iVtYUXJof
jvCw7socSQmVEZOXrWZSSX1h+b+FcufhPH6mIoLGYfnSkxj+lVKKbkRsFBZSDs41
Q4S3NgV7Z2MgWj41Xc0I1oqfrzvn5QhaMaXcTvjit7r4Wr6v6pEOgst8i5iiu52k
RxyhiYKEnYLecNDcsGF+DtMUCxpY52u7WDqW/Zi+/cvCrLdReAFd1exzYXKIRukR
WIJqgwuaP7zHRnYQFkhLagr48dUy1vTUCHTOpGJ6DJuuUwYeqIHPnmZxAxB7QTds
Hvdu56or2TfFEbKFkITG3YLaJvDQK+n0xZMYBFwj/J166o6fUK0cLsm8katCcPnY
ihb5fe5BzYKy2M8zX8NbAWpd8xYxQMC3OuAG4M/eTEtw1rICexjAc+X8ushsA3B2
xy6zwhkIWpv6D5YbVYbJbSWc94GkzoD43EKZ+KWn0t79TruUBWeq8eGtvPvTQE3z
RuiSl3lXrubuBBKQb/ugcAPd3mg/dVPJz71EnkruQrpHLKBRR2yEAYkGGL97scwU
6qn578ZGe8tgWnWBeZwnBH9NiFH0xUityqOV32V6+rRqRl2aujcEwR9Ii7OLks29
Meyj4j0/aszxM5FzWKpK246y58RJIFowNTEutVlvMZZ0ZD09qQzydJklUEHh8R4l
i7rZlPG2BSVgjl3ZaiZObhanRNAHiyu+WCS0zzTnVaR4YZwZ7EMjZHmyZJHGs+dv
MeK9EMELN9mmQgaSPgkb1u2yNizqwZVXFNFJQ1uNc1ZSm96kuog4XR5xYWNrCPlt
xsl0u3ojyMwlA1ghNfCfEiUr50FoeAAA3hc4a5VxHbp+ZUlocDSkCiPjyOWuc7AV
OA0sKNCWNd5MhCxRGAR+LuHHi9crytv2rGWTW59UUEUGCT/LrIuSzZa2p6De0Cat
hXYu3rmYqiYwuC0I9c0aUZyhtJ2vSUn6FoTqj0ESR32vCUHIj7Cdx49URa1L4LRa
HPqZoMKvOfIM58Ax1FCx0xxPB9/sznV3cPYqXfh6qii2YTschSL2k/6LJDdEf66U
7yYtuH59KQrEzpR5BbQ7VbirENjw1FdOr09JtFHP1nixHn7tmgoO/YW5HNZVWt7p
U4OZTYlCe3ZirZWUnbbIuJ86B4EOgjEPlHNrgF81kknPi0EDW0iKpbbGro5+CDLI
j0wg0zDgBvo23yffbpY5jdqvQ8tZMG/X0EzDX71iWa03lCfRGMItr0KrXwsmhhf6
b5YjNtsgl0E1g++GSRhGKdIUwf9nhdr1AKzeC1IATIFWdraZNNLP1j88lhMHgzlQ
4S+fxA10wZle0yPRgzaP6O6wH9+IO29lc/MT1No0XZkDeYaVjQV9O/Yt9E+VuSfO
YSTCq+NEbm/VruXjAonKDJJVK25+cLkBC2jG7vN5ZfK3mvx2SZ4w+Sa7B80IGadR
JVvx2DMKfxO9er5Ge3ZFArn7cHpPnzSslgQgOiAmZUBHJ1BILWWjlV8qNSxq09cC
16HTVkmUCpdPyddh4B1nkkuz/T2wA9wfK6G1yLV7O7y2eUur8y+t6AEoFFpJ30Lu
Q/3D2AbFBGYpgBS64PbpSMwXlgXZCd3Lnx4kyAFknO72X78kMG/Qh3sHlN5TE9L4
WB1cp+7NI6lYWcJKdNXVx3X6GGpjhSV+VE8H/3oqDS/eJo89AuM19QHbtCdtTBbw
IrnYyciaT0BmJflxQAi62kgHCnyuvwH9vlgNOMWseWqJ17uj398Qqp5+3wf5c+lf
rqgc2ftIJJR9nyY1ZsfAtsVW+8sUHBQ/Nwk8HtzjqVeM2zNZdCEx4NKa5/NPDm3M
c00TaNXo1/HvYd+QAkEK4o5V2bnAWBSvNbCdCvxieGOFVgpTwVcBSotgNEOgkthV
HC5FQpuxRqvybANloGzJi0QsBQafF/RS55c3OwLoX2T2pF43EHF0sEjry5p/Yfzp
I0xwi2EutWadUNGwCbMhacQVyyVjz5yLxVWVu9Sq4Cy+S/dGl4qJ0B5m/P5rQKBU
yD0o1yk3GxMKKqN1csJCSJX+fcBjuwnBvC+FGMSIeujtEhPt2AHsbUT+PiiYm9kf
FjnNtRaEqjK+SVYi0WaF+qleEtEYi+AIGhrMkjXCM48CmwsrMNdtGh7FHo9uhMqd
ea75vCd2nZUVfA8VJV006dgOZqIpA99Kv8rlsoNEjofwuZM7vXXButXQ2zWxNXbB
dNbiYcskbS3iG5jl7VhuHTo2D/0N58MFOLLrr+GYXM8PxRSEItXrwKosA7xAmV9J
FZzpFDKnWXA2qRBiXKfOTkuYTItNJbTc5YmCbxbpGs66yE/xVF43ZYN6QQL0nK1x
5c+5xuEMPpvPijf7giXuVx3EryPgGwmkYMs073bR20xac+ySD4RZbE8NXstH9EbU
BgCHnfvSOf5D5UUV4ueeBo3tsbuvyoYABPvJPA7QtAMaaLe3nkYHLs8wfOLp7Z9c
UnUciPQrX/y1xWP9w8D6dFvgOobKo+sJl5fU9PWMLqyPgu0GVIdvEMzXgSjjXvfa
/+DTND5lnKAMVHovLhPXINzANGYptiWIB00zTcqkL3jRV9N+WzX+FQorw1Wnwh/5
iMiyz75uozMUMcGg4TKAD9xHa1IbJbzu2HwZqv7rsWG1vw+xhNa/VS5BV/Zorsh1
YrV1BKPvUUrCFsu+dudVodonuQkvpPlAR0DdKn8vpd+Erz9kdeHSnS6TE9ZXjqe7
iGkfJiau/labVfx19ogTIJsP0IE93iTl/VJ0AWhuGt4locKsgff0TsT76DNfg7qF
8rcPcepQXU5AoD+Ibns6enEvxwUt0dAbTgxvfgPaAsXjhBceTLYaYYjtpOnOfIgI
L8wkKi+EL5/sLclpxA/0w2I5Km58iFYHcmof8FDhbWVRa7OL0LL18/l6SbXGkVfz
tZF0TBYhFtBc0rQC+TH3gjUnl34WdpXZS9EGJdTf3JB7jfWYdqsbZviDrwq3Bmcx
nR3Bji+ijKfTRfLc9mPOY0TB1YFf4s3sKB/l02NnNKlXwKo5UX3oiMqUMMLv2gfX
e77WRRBWs4LS0oYZGu4eeR1IMYdN5ivUWlF2LbL3Vu75aSyGTo1rv3UzxJnqkwbh
dLmew3Xl20WpjCapHMrVWyls6Zfhx6E9PBbpDp+jm5BBOHVHOGIRkBCPyy30ni2N
1XZJzt6gZoQcAZD1/Ib3sPTN054WMzWeFdcaJeFvINdh0rPGfgmf8o1jAT2u4TRh
VpKpqPdqAu6noBsiMq7jnYXeJIVBDbKxXQ2hKHsXCvJZJnphNN3Lx2rAQ8c5cYyU
rICiolQkShYV1WkP0nzA1tNyOWJruwQ3D4V2wKiivw752A0rN1wzUp2eTpX52KkJ
9edCPrvj6GAA8DzWPq2BM8sHaPz1oJqZkO48E6orthpodVq32e4/2Z3tD4gHt0dv
9m3STqw9AmG7QxozQ19KdlCmjVMn/JYIL9ecgHqRt8AzBMul1VU+f5AooULogDnm
7fmAMhbUQK8fkVhRqoMq6z970/0ObGGNq5BLSSCcsYhRerr7AwI7A+MX8gjSiar6
1gdOVwn78BetnnZglIrz1Ob/91E1BFl5yhwJEXydhm+sW5YvZqvz5VXaiTLJwI9v
T0jsbx5Cvz1KXiLNuxuz4WSuZ554o94O6i4pbcG8zGeeUjoTOU6kFxZt2rGkW/bU
ILKZHPPr3Ka3gApKhU6Zul37OUctGsOGGDFkqtV78bjfbl/vZ0zamAqSjVFLcjjq
wQehEFUyYfcgOqwhVCqku5824mEo0Jt50zd/PRAwu6XE6zpLYIreANADvuqQwGWb
1nPBvFwAogt5ZRwrgqLjOVKsTjaU4oRdd6fzu71UWVgSiPOtaI2JSfsgQHcvgVI8
C1UXwFmPGdbehs98xENgnwwuQDDPt6bEnuP/VCwQvdtyzWcupfdXnySZR1GOk/ml
5n9Ppoutye00z72TlwPy+1gfQRSXt6aq6ctCI1E+0DcO49VRAt99Yr47WkQve5Ud
LPky8UubSb5lF2OnRmudNKG0mxH1CygmKynMf/6T0QrETDWvMjVkIBmRUoL9PYwf
dCfOxVvdzRoUrs/oIMBgodhn2vfiOd7/3JgNVGCGuWauRHPL2K2xpUIPoBUr9Z2d
cP1gusFZ+tLrCdFJhwlfNsJkIrPjcBwRFzcRpdebfTspq8MlDUdWpvjdlbVRbwNe
RYOK05CdRHWsaTJHn9DDluFFND/S+d4xPmZDCouRrIwvMmTs1vsD8yhNyPaD/Q8m
pd0JCGgG+rmjR9zqDxG3LQrl99CYOqFMTP5MLimhPVpX0qDIbJsCeZB8nVPOO9ID
d5RqpW0R4jThNPhntVLCCf2s20EaH2JfBudB1sPzHVEC2LL+jWq+fjCc92Hqr2FN
yzHbdkwSdj0CggnT6smGqaqqEsN95+fT6tnzQ9uHQthSJ91GaFZCeOCdY2jcsgnN
RUuasuIEBf0fIyCyQ3+YmVl/kTjgQ35APKTRZQRjMRLqwoXoJ86CUC1z0u4uzzDp
Lvh0tRJSrkbe7KqyeEYubf/MiDMqt770+3ePF5JUM+r3viYnyEgHSWcq+jgKPaev
E21/6dWj2qx+okxcLBmYZSVhL6tnVMUqgdqs5SxKfTNs8Om7WiJuaJGueAYmiKVD
1bq82pok8BUKf4Mm1zZ+6hCCsvW46dHbaGG6CB+4PEOFUBIW62enIvS/7I6CFy+s
rj+Mscj1y7xu8Hu9aKIVI/dMNO538peg5dNMVuqhFDSCVRTQhR4PoVlMkXOpS8Zc
9wVwPIR1a2AgRNCRbZ1ehaGtulQCAATHucwVplTNzPRHEUoc1Vr0ZBk6WKB1juR9
JIRz+Qp1s+1zNkGub0vvR6gWT3TpWUu6POXGIMQkEuJzYtSWarTSYx1cooUgkFOh
vLRdHRATc8Ix9HYfjFX6nX5wcdgEDwpDF4PYJ+MPaiMWjXHgmusmJcj9BZc9K48s
8PqyluIbc7MBv0qIV6uSS3PQeHk+b1kKp9SaEG07XB46XQk//lbwtgqtsxEJlep/
eQyXopJbR6QP7SzDBfwu2fMWJJgR26nNLODunTI/oM2cYwegBcJT22gFkDvtwwD/
ZjRYOGxCVoXS9EJtNqf9loX+80RS+gRlyqjJuIpFTrmGy4ONVb2Vb1X/o2vu0dAC
wiF4ZCRglV1wTab8ASXOQNDTGUj02fxreOCG6f0jMHVEhGRrhvQkEW86do7yMFbz
PaS5JzaM4J1kuY0VV75piQ9vcaaIBT+eaAyZa1ADk+o6cqG7Y6eANFBUpYNNRjFt
IZ5vREboo7FctzGvSOLVGlPn/vXqV4VeSlp30To+SssP+BQHT6oRCfDK40T0Xop3
2NfVR5uSmQvdh6+dR8+xjkT5eh+x+6xfskHlk2GTzzm4eTk4xiiwGYRuD19c60Yg
kmzboR1sU643ogl+INUKm0+9SWF7Gt3rjxQKF1avT0ukZJ99sAxjFOrnEaENTVOa
x6/+eI9PikCAy6UBKws7K4Kzj5XNjQGY3r0WUNPmcMwW4MsGKYUhMe+k6A4v+Npy
TbBRsAXzDkZYRpJ1cuxbphGX4nuBjP2yl91AJlQM81o5CCIaNAqLUYPrhf/8AIo5
F2nTWmUKpWEXmsciNmb+w+xFDWaZt3cdA7ELBMkg92+qg3FNspMdU8CS/NysWzBe
EltWNXLXkfwFrTEHDnOmbcBzk5lmktR7/74YwCJuatX2ajGam82I8sz3sn3cBmv2
NluhRprDnwNJ+O6pdpt8qtY+5ZjqM0TCk9SHxmEHp+pqMnJMr1k2GQoqdaHtrX00
jTPwhgtQpEST1fCOtktcQ9uDWPIGPRy232a4bvGHaq8Ciay8Y8raDD2pdXP8qC9D
s9HkQ1Z+RH01OeAmnISfbzp0HV/wU/OYnYZfdPcWmWxFVKbzHcILXnjpBZPR5fR/
aoSRQuViBPLhTIxEPhnzg/7muBd8Z/C6WlleS5jd62Ii14T28D4+Y6/AphT2B88a
Yv6JQ1PsXduiePbQUVmyxMCor6/o9kxOhlErIRzm59jGN+5xZTceDOACREjErtdp
1O2LyQp3t4K5gWXKEbfvGbuxx/OELFY2GoKZ35cd2SPJ34fJTcxMvi0ZS+Vzl6VD
dX4TpR8jM0D1n89w5S2A+fYhYsYA5ePCorGH9nOxprmqDnweHXThmHB75XszhUiu
hvM9RHyQwp4ziyco4nw1DdAuTphaF/28W1HQzWeafaBka4b+o7cbJrI9klJO8tyX
lH8ObAEBCTKZP3of2k8OKwWH87tg9Gq57FtzYPLtKOme8xwhz/9yq/87BeTqgXMB
wyzMCkvzCZ7LAmKB2WqBpayhEXFll+I9HKO3tEtd+Rj0wjhVSsqor7GkiymBYl3f
cq0j0xzXadcyvGWt7yfDpePbRrygfMiRsKSMiIp3ZujHMK39kHbAOBzaw+dq5zLn
hR3EyU7YA0BTmdZ1+D9MuvjTFuE34oubTchi0AG6sG3VdqoS7ziNPcI5z+rXTjpt
PbkF7PjlxOOG+qzoyWImoPOmRnFCDqNz83zo0vXKCpKxVJuPXDVCv1cVSSxFEgMl
KbzoAiqHxVaaac4vHoemT+KdDJu5ynFL2W2baoOW7iutmfKPFHFSCCclH2GcBP6a
8Hb0T/6Bc3lSIIeuKSn1sm/LcGhgyaZagnO08xo4sMrRhm1xk8iN8kbr39YLt9D/
BflHq/QQaDYGeD02iQ8huyBpBRomgkyWl+jhEW1Zkn8wFZ3ZMEVSQ/TOQEWfD5bP
ryllJbalouJxZOr4ee9IZA1F+WmnNiGXVrHyjhDUiOr2oZKoBbxC8pKiameTxhM8
5SsanTHdtMJ/kQEAzUPtikMIgMT58tSLNH9IY7JPw/eUVhJQC9tmhYkIcI57WKuo
ywsDL/PEo+XIhGtqKFiW/oOS8bGXaPaFJsRKOoj3odCVMUSaJC24BcdmEIaBM11E
IAEd4Qk4puttXE0ighbckt3YxKNVzP42Ry5qqcSuXuaQ0rI2UUeCfixe4gS8jtjp
jaEpnVa3jJZUjTSL8rCELecw2/96fBlK6wfuxeo0TW/tOEKP+lkusUwCiFdFXhH5
WGYWR5ot9gtKPuWKbcnPQq6u24GdOLDpYt10Mjb7BOnRC4+HeVr3Y3cS7dqNWLWY
PYhoCfOtS5FA/CgsiLwWUqpwbQppgvglFjAJnsqC/3up0oFqEImPUL3+1VHtVNIt
cFPUDst3rYvLPerKcdapf6v4v7HLjCZ3tDfKVr+p/ZF9myZLh1UJiYv1RbDI2jl7
igZu956husN5pWvArMEjcVlwXGskPcES8AaVmoIdGXgajURiieurcszDHhBOdhaq
M+8UUM8kUpUdw6EmWc8vurLqsD/S5cYtrwpovuuos6M5HqJc+J1eEn3P8kAtS4mO
XMLzZzYCxls1rSRWTPkcsdqGADJ5zHFLG/3CgtMyknGHqnYthghOid3YgI8LJxCN
5Lq+6sjBLFDzPXKgN1K1aSVQX+KK7mqHtNDC1VGpVgUvIAOO5KacG23xIiG7W0i7
9c8zMq7hyHceZAZob85cYzqIx0+nERziltasrs/OQVoQe2Kio57JUUyUU/Bape6X
cD3PhoIMCnUTkRoH1PvlBuLLsXRq91TT2+KwAk8MAOp7gb/e7hapxgQJ/w/v7rj+
uAISw7zSiT+zuAOogsi5KMWZ4Lk5215NBYPX/TOYcqLnzxXIUxFFJCGwsUhxyG+Z
skOl1VpLKDmTJgRCCnqhudP3YI/PXDqAsNRfQ+3zV1hYiAuZIJd593VF0GZcop+C
oKz15B0L26ZUKZu+brYzeLP+KPdXpxytnVTaqucC+zl33ueay/O+L5BAt7URYUeq
MZoirPXpP1c6GmZ9ldrqzAJeEXA9KLJWCKXxHOlYDf8l4Kfdi8REZtBAKqHKytwI
m8/JlRUi97w2wduJIZCS6kN8WRwSY4rTvSz/1Zq3Z3kq+JpWypTyUV+/44JQm3+o
KMw35S1dDOx1TgRuCOHEouOh6mrYhWX0iXT1DZegehzQBqwnh8HfQJ/q5uJXvPiM
XOrccAo53JtUgPsCEU8y+X8dhCBGhXtzHw13r8LMmBEbJ14HzNXbIbnyFr9M0BkO
SmtJbxghWaN54ZQoJoS11PC9vpd8JoN2nB73nuF1aK4o4ef2kWq2RXIfFnDzfcqF
zT8Jau1E0m6IX4NnkuqGfcLO8V1Jofzd05I7s0oqPChquMzmHxOFe3UyQkZG8wjd
ttG/slGSbZQ/S16mkNWxIJAZBiBklaM66Ospg9dGwV/R2Z8Mu652urXErtYRQQvT
Zru4hRJsAIQ2OnI+YUMYmOeWTJNakH0V9uwFuWmM5paiXVgsFXZdM35WqiPdnLlD
czBUXZTLEhwgXL+DdCY4izVBDvLFD05wLl5btCQurtDFOx8A3pbDEQ0o+4E0dhI/
uduxx42TsH9jygXuTvkmf4U4ATJPecqCDe8jGEUVp6pr8D5NteeOgcFKQtWf1iez
7vupSaTAt9kfwHXTyc3OU+jAudPdIv6+hE5I7yCjNJq37A8Jo9wlvgrlWpvJ0OSC
gWr5QMQ8bIlfheL3xF4lVEfVp458/GOOBHUMR049ncNW/KYRGd6j9/vqAaFIqT9B
e5jKmdRKEyxqc8zCkJMH9tphqYeGfxegy40Arc/CtRv6506lRPu90uhadPGTkXJK
+SQz6qSI0A30AlS3Jvx5HEW3h08nGp5Gk8fglp6PQZP/Jis9C8CT+m3asJ5GxuBd
4gRgl5cGzubaKWjwiuN0XDHAIYTSLMhi4YEn3Ch9+7W/QsNi+57YNBKldvqlhCH+
SNNEvZSsBpIUCPcClYup5cEKfSHqnH7DcanlBFNOq/GAUzl3VGWUhJIiB/cCP3YI
s6p4H156miNjk9ZVBmr2b4gJtj9vqI6BofvXrgFbjp7f4oDM6JQMKdwx6TYVw0Zy
q5e3t3xiXCcFpcArGE1UvueHfI86n58K1SM9DgRWIfFJXJvvcbxfLyi9lEqxTKg+
pJpAP5TjOjWaXLHpu92XDm/lhYLaT1yTJ0H4H7c87Gq+oQDBqcYH4m4K5oaFfNAH
xeysZYjzYalRvHHZBQ5blbaPoMPvZ/nNH7MB8h7KOm+5q2DaNV4zFBDmGXUhAxc/
MASHEwkMhUiW0iuMWLrG6mG/60RNZ0O2Zn9OZR1c0THKu6cKa32V39LHV9whBivP
1LiAR7mtR/VW8zRISvn1Amsb+XheZIMpzl0Heqct2xOX1cDUpzx8jtElPUI9inb6
dnabHgZh0f/BWBM/3ASpTew4N5sas/PMNawJxe6S780uYOvTotcnPHiKHfFfHXwI
wupCUd9HbUOFJ4CieiknL751mb+tQBGrSo9DJp0HL3uNTXGv49928u+LuAF7iXik
ZDPnkOu06O1lO/Doxrih5L/Rjlh8RF47fl8sIlKn9F4e3EaQdyQv5pbQDpCCyYfX
bD7arCZOvEet51AEcnL5NbVjfV5zMR7wqkDTzTEhA4XPJ6Vf4oKyPVDcBKiXPiWr
ysg77LKYxqRJcOz7gM+djpdlAjCFkOT+7Muk7dAtnSjP5jcR6c6gkntIF6zYSvjn
cGCFT9+yI/RzuIOLpWln/FT45nYMI/dr/pKca4BWsRABkKsUdWHxCeXbyOO1+10Y
Z4HEDJJWhGhH6OsDWYzmR40ggfNfQrq5OxrTNS6w+LroAs4i0wNey5iyKLYv9bc/
oah0Gcvei/m3XDQMMgppxVLvwW59AQ9hWIr9h7l/k5wWCCiFrHYjgAqlt9lqXEft
4nhlDT9aqvSSfkn34TGMrqDlKbWJwnfCMrzcs7JZ7dQwHzoQVJXj9DmP0b8Nia+d
jJyvkDUBhUnPKtCl9Ur45xvv9+rrWjRYNsZl214zkIpuZL8miKVXkr0QMWrl+ZQt
EjhXjWk/wLU0bpSqnFXkwBG5r5n0p0m/uqumGtzdiyQQjm6BwqtA+ZnQH8sa5G1B
2k2blAxOPNeu1mT+S2DkJ7/9Z8UimXW5sz5O50TT4PgyzPVALMZyxGz1I5qFTMTG
CxCAQKAoFGGPuPDyad8ap4uNiwvkh884TE27E1h5M3BnyQGa8Y+p4fSUhs/oXdbm
/UgvJ6DV2SWbasamguuJjP7wZoQcGW2IUzuXYf7NK6O1BzOTZ65DYVFmbHuYen+p
Q2PjzV6Me6gz2e7GriChBqMn7CgaspQChaJwRef5JHHXVxm252tSyjmLDwYE67R/
KII9qB1hOPDcVZiKQrjo6SEHzpqfhQLNqAY+DSvl4ZXYDQ3ZvijjjK8BwNdf4GUM
/4oPPG+3+CBJWRrROqNl//5sTzd3RaSKcOIIh6OBTi0iAsWhhSBdoS8R9PxSF4a3
GuFIWLSvLa5aB+7LnFI6eVb8hECppr73T8bEhXLAEomTmkwt1+9e/PGwczxTkQ+Q
nm1o3cCYV4+0RaELCgXs0OqP7rt2rsOdEMQNPbALbENRvckDjqOW0zNy38R5XLUF
m9i5kSXcH7TvGnY9FDo6P/ffBqJaHiKTSWkOPnU0n/Z8vcbNVRNCpvip4kEbau+a
EhRtbqXzExRRfI44eEjc7R4WZgL3mJKEamYfNKhXQmO/Gqc4v9l54Eqc/9Sn9PoF
dB/3JWsN0ASnvbeqIjbAH6wgoG/sriSDi/ywDKXbSibsBVkdpRV+RlJvMzqDAewq
izvoZz0vpnlkoqzJiDgAHBgJNq2uePG5uBpcZXVApW3oIcztKGoYF7LxneV9yJkW
NSE3gs3Um1/U+ASBBhKX+tsfhGzEoExbyoLkfhsCr8o7D05EjRrAEJWkS8obiBoW
OT0GagfwDraDbPb1WzMTyDhW5VgGQR1TdF3E5rY9Z/9ixGTbPsAianvSx1RqBW9J
t+6kRXwSOmlPqMzWHrE6dlMSOyWdKy9BBRtiTYr9u0028hpil800vT1UoZ0EYhEC
LctYHbJKyTLdSd2mh+7ga16Qdqubcalr/A2oV2/3te20diYtQ7Wm2TOVBEK1Affy
qXjJL+JHElDZy4SiYiTykGMNK7+Dey9mdBqCm6CQUTD1ZPrlCVYCt/04BE5ZZtO0
Yh4R3KKSLKBbP8VmKXTN8AiPATJU2JgIrBjGJMDMeJ0So+ilmhlBn5s2n7cAak9G
HABf7laO/jbewXRzrtX2uyid8gC8443bRyl9pcJvfLWPiy2WLEBrpy+QYFvfABG4
epWmeQ1sSkqAoz64WybVpLZDNYW7t1HJgtAwIfQztY4hyDfgjtrHEhgsWaoyBXy5
FDKLiagJKzLXM0Dyu8iS8KSFxsgVSRgg//kCYM2zK9fdVRa6BHQZcv5TLMvshQyu
MdVGR+B3aguQ5k4dDHJJOrlZ/M1BjlGvNW6muTAIChmCReoEUHAmWIR1cJsqtV9V
Q4RKBca56AQT2+JYZRJIyc7dKe6WNm02tP4ehS679wSLc7pc/Kf409j/sW4E1Ubg
cIgkDVISIv78gZ/c2w3p1CmfrnliptMKKDt3Gee/H0GpIeBRLp6GUqNFdbM+k7m+
vOy9YtL1PFJfUSAL+3fLiLVzB4kz1M5qjHH0HwXKllhVw13RolraAM2wDLziwKzw
0a3Mq8Xh+iTzoVSJo9nrdgYyyjuSWl/Q8KB6oXUKIMnMJn+KHrxZt7dSK7taGcNl
lPPFqV6/H2lEL0iLVBcBGdEHRX/oASiiLmM+Mc6u3OfsQFGjYhiNvTO8z4fzCVEz
4zTxDFWQ4yOU7l8TEuHof/T4t3XbqOa3p+2dpBiTqRgacQlpF4LtUTZCuKBLuMkN
UAaEwqc6QkihJNqjkESVFN/29VtEYH6+L52ZDh90u7H+ErnEWG1/h+KDeeRBEZoY
V1sSWKkHB1up/ru+Q0fq/eXe3om5aQQ0AIYGQe5c2fvdh/IRCZ6hq2LntNEfv9bQ
l6vgV3vhQMuNDLjzSV56yODPMW3eFKyS79o3p/r7JlgVagT8Uxrr0qDJz/ARQ/xY
O+tLRsaiV/K5CAHyPlOt+TR7FsCc8NCUrgtYQ1GKs2H/Fo6DIxdjMK/4YFyxTIlu
dIrzncNT2SHdnRAvgJTYOjeAqTmkoduovl8V5QbtCfJzCsLrm20bw+gF3NzaO01G
sxY2hOvB4yTtLOoxRlBHHhQk3HjfRoJJv+Ylb9rEj87wFl8GFGQdoD1NksYwxwoj
CjS04BBnkFLLRK5RKse3QIslqs553ro0r+FiUg2n4odABfBq4wPlXGyXzp2V6lm8
H1itEBVfe4uJkkKGaHC0Uzt5ZlAVG3S2SW8j/qd6JZQV+wZxccL7okQf8gGgfsJq
GjfZLbhddMdhjVnXb0PdXe3jCosWlNE+dWm2wxxF+Ym7AHIKb67YEHkxCP71FHvl
iG1D4p4G2AmUWtyZX+grFNL2upRZd7QFZghVcy43zkIe+USbsV5h2CfenvEBFkUL
nbqkNADNhUt632bHdxZCah6tMZH4pQTxAZ+SjxkS1+Kj9VAiN3zr7c9I7RULZcKU
6kbciLuz+jIOyvyFKJQ92WX+ZLV8FDQ1TTA0k+XjVKjIU7I5z/XOOF+fia4OgBAN
AVh72x99gRwRK4ObH89QWJ1+iPCzBZIN0nySD8QMCH/WUOvhSFOrxzwebX8B232s
krdyi76/nHxyYmlYKczl8/dZP/DjMFIi6E3lwWDELF3rEnu1fcT3Brub45RHGjmm
jFM74ZzOE12oqKGBVPKv5UDw1T50pMha9QLklWy6nAOiI1IiyKuQ/C6mvLj6FjYE
kuxW9H3lBsfaawJxnMCmR1r4GLtI0JD8VljhdmOH32hvcDf0x79EXLEuct5skkk6
MFf2zZQo/AWqJ4qCVoqA5/cNmQPCKcQrOakh2OlrxhA/rMu1MJrjlPJTJHST3hOs
itrxUmfo7q59hp7QBPutoY+bFtPNuQE5WE1azPyneYyTE+uwbF4BVtMlIgaFzdWl
JXevMUnfWLBXCNvW53N5fsxcaN5Pn2jUkYhrYOTZLkIechEvkMSYaGcEXJKJwMbm
ecdcKEj1p625lMyNQc2GA/9Hz8MIgNNJsBpRCdaGiuslR7ii1OKRA9NQ9LfExxCq
v1VTia/eLO385W3j7hAZjfH47bmtgJ9SiL20dLzw7aHdMGjKZ9Wo2dI7fFoYw/8c
M+JAOIvxTYfGY/JurggTADVuIIPzOP0NUBxfR6Fy8BC5UrOBreg4WAA82a8R5qNc
tV72og7UofAHx6X+4tVmSg08INlxpsmNFBvDcr06cBwUzY2PODViUsZeI/Ei79BX
1rY2+uerkZUmk8lqNJIBwldQd6lNRbq4a2C5j66MIroEzwbUjP3C37xlNI8iJNPe
GYIBQysLR1dFqrC9QNHS2VBQCaMlnOBPpMUw+Wf5HdT/aLPr0kW+zCB+aA8RkJB7
xUO5/KHgWPldxBP5UFDs5W6WsVFr2v0p/EJeYylbyaT3jHPp80161lTi1SWtoGf+
t/fZyAhWpgscJaxEd8h7jsdrjLcExeL9Xxk7eqefe7xGAqbyj2jJaJjo8xccUEA1
2/mn2/6R6ZTMXlBWH1prq2Nzuf8WAnzfqvF8ij2hfUg6llJfX44571HYNLSS/d6x
kC7fTJaHzi4uZjsbx1jHGuO8cjy5lxXhN8VJQXFZgNaF6xfteW/8xw4TtgBNoWRl
Tpf4/x4G867UKr7kzKqUgW4u39Dw55jZfnm1I956qRLIVwndnEFvcHEZlT4+qAi8
r0ChtRUDx1vyCGgIYn4d8mWQIxzTAitQWJC6+gE0JuFW2PUhUR4azDKLTMInjT70
MOqsFUoLPay6TOW54+jobagKZyz+DLI4aS16a5YgUziQi54ESDgDnfBgwYcxeqLK
axBwzYe6aQi+5E9oYO5xseXcCefT3gi4b04rNU98QZjgxACvbn3W2xUB/uWWmpha
birGWTAuz9RvXdl7NSmAXRRiSYVjLdls0xKcm/61mP1maEDEmnBRpgnwMs0Ka+Ew
chqStYFREYah9dLzFO7tPA1H8jdeRR/rb70lvuhnv0Tl22cS7uHPetcEQSxVqkkf
e9btVt4nosL0WVyHwvCynmhA5I6XTQ+EDPqy0cF9xqeVZ374JkbuychEZF7+275U
4i4bVGa7BI8oIDVhO1aO7TgsXrOB/GLBeWuXA92HsOaHlxoETs2Q5wORK4gufbv2
Hf4W71jnOLd6wH5nkUCuUcY2P0ImIEoIYJpFM9qGcZtmdIJICaa79pZ7vc5x5x1s
p5IwW4LmR9O7kDuOKXgUkyX7HB79DUULF5URXHR9gJpdvr31BxVdIQK3+hAI7P9q
oftInez4gTQzrSQjZqR8Q/sgT1R6H4MNzA4A/fhsJsY4n9bVAok1iu4teFikp7YC
na4WhbIkrCr3AAzHJOHTSn6ilTjuz0SmNLKBBhgFFbUgHaRrz0BFBQ7WeQFE+pGV
9BIzlmBikm6ZOG75fOCjUgEjpZSJyPzusvI5K6EnDP5jEg622FGUImJo2qdC+Apj
Vr2AtfTuM2MTQpeo4/brqVt6b9wnIutZU6UWmNDHdOoP74/y2G4qGOs8RDYASRNV
Ys7NPekmtbMzBDoy6hAwBh4vbzSXlhG8wrwuh2RpceFlWk304GOx7z5Hz8nBma4I
JFPbsMJhUpKus5j8mphL9qHpuQhbNFR8DoBN9DaDMlRduzYegyQ5lre6n+mUPlh1
HiVAfZT9eVV+eHGYOhBDf/OsjfxAcT+/uJ33KgFzCC51ztFecRAab32kYcW1CqV8
adWYdYjnrBrMnHSBVmRFqKj6tkMzOBumokgnY+lKxgdZWLnTSQvT/6wXT9nDO1Ca
EUXIjuTXORImQ1Cz+TibYjGOeMJTKPkuZXgR2WkjMzPo3xMM/SGidLB08VtL7Lv4
yH5iO6YaM8Qe+XDLwj4DdyrCuxfMVblbnKo3RbBstzi0UrzzmreADcZLEqrZkwcX
C4EhlM94gX9aDaJK+flDJheS1RUg8MztcBqpl6lLdPWbDtH4jjH6rkprIoYCOi/g
UXoOhTZcrzELVeHOC43QxlJhJd2O6n7L39DDqQ6ml1+/LPd8wP5kyQSlzmOAMiZ1
NlbTN2lqlUi24vFmjZjioFngTk3J5b3vg0xShJu4Csoh8yl96p1PUdEOnEyySRM7
KUiK1NQCkHh5umab/luiksQ63m0EHK4zvuOOQMQSvHXTH97pxnpJmYzz6jJl9O8c
zzntA6v+G0OqwcNCpiRDFv/IpZ5di5lIpcueJXM5S1ajgvUQx+ttntTs2Evdf8Aq
dbeu7X5FwR+PM3TRrzIjCSYoTFhS5wMOJAykPUqYDlzaODzPZC4+zDSlOe2nTtCz
JJc4OdJQHdSeA+vwVUHOT0RnRGprSQ9Updx3vDa9qa8lXAWBNk3JpE7163M0K6Jn
dvpJ1qGGiK4yntuqEvjPSzxIscItH34Kmn+yo4NHwQD6b5mzpkRKdUOI6l1t371i
kpFtTdRQoMfKcRYiI6EVURkasbk5VJvTgOl5d519h1obtokPwMT9ukznY7LknHBx
a3HcPC2nxYUEH9iScxzjQolelvJ3Rqo1Zl+puWFv/jDOOSllNwjAEsdj6rMDlwlG
RMPKthafJghRjQPgCOcC+3IZ5snL/VrbrRv8aEAQJCDkWx/iQdOoMonnPFuMmY1D
ccP3UXEH7f0SsZJoONXRKlOYs1ZNr5t6jFkq29RJVdtROCTIzGsU/Ha7ZY4jZvDj
whCcfa1r9Phuqvie0AyzzRTxtQz7V8rZ9ypr0/dJWM905u9pxiBxqzuG/p2HLUpI
pyM1MlusH28exF2yH7rBBxbkoBkdhFh7HnWD09mK3jHXxnXJur3vssRVasHgbB1O
yesLQlVny1l6uVijpxWj4LOSqUwXQimr++VMHmWYTw1aG6Lk9rag7G4CjT/Fgm8O
gkooJiQ8U4xeWFMZ71/JDeLJIEUT6T/dvrxGbGiWvw2udG+Dyd74Ipmpn7S2tTCl
YAPRPImLs/laSuEu4pBsr+GD+HIA5NX0BBt8Z/K0xi5q3Q+jOb23+bJEkCXE4TPw
G7aeqOSojVJs/ZTgpsXbTV/RSY/WeQca4JgsJa7DKxjgSUfOiLups9iECDtgod0A
9hUyDBI2ZvaRBJH+/05D5g/++8jzCeGYHlRNA3+CSRWf7CfG5q0aNNoxhowDtPDq
KwvoUIgZFFv2JshapW0Dzq3Jf84EVI+fJQHy7rIim83ueJfxSMFQ6D+5XfETy0Ue
H8Twop7xcwj+g3iwe0Lt6lRtkvw9ZQsbeKq/PWbmwgJcnDxglyduhxGhwldw8GVU
5b9XZAIeXXtkWb9Ywa6zqKSNLwYQi7o+OLi8W8ipu684sr27mSc0/sNoC8kSANZU
RCW0sz5mw08jpNITlbH/ENva/FtUGPdeWJOnez4gQOhYNS251DtXKdFGGvjRMUOX
y4DqEKmDuq0ZHaA4LM+6mYS95MAEQCZFbCrrmTKSpu1MJi1pc08jAgBFag21CEZW
o6GrB2W5q3zOIRxFoW/dYsR7N60H83qIl9L9Cc0MAQaJOAH53znKkFOOLQ/qbgT9
SKPAL/mbBOSsru9aFzHcoVKO0Oyvr78rVGzCDHmV2lwa4iR6/XLAEZF3feF6HrIF
9mWay4EPuntAaOiZHXe22PtQwN/0YL8O098aII0KcZ3xFsaZ0oE/FZTi2x9bdgdx
kpKEhLFGBYWDQRPrjjhZyI6SlY7sN96slus5DJM1AMFzG1TkDIwnN+Ajvu9EpGBp
AbWOrIY2ojB3uOVkmCwU9MX1A4psZYMSfYb0lN4QF6fiiNJNo46CpprqP8RYgX5H
fB2hPgVsx+3A4yH0K/jtovyzuH3jXZMUGDTIunTJUq1Lim5dZurhP+mt9QfXKnfW
I7XErnhuBMsTBoyqUd8sYdZWjt8BafOhSGGTf5TySp1yQtAaOU/+sAObjpxnFzpx
Qu+0YBDRjUITViIgT7hSCaEKAR0tLsipQTO3eC4PQf6Sa5k0dalRtk1qZ49SnCLN
JTjElRuso72QEDEVTBvvvDZ2Kkd+S3ybV6j+KQx0rRRNz9Y90Xrj02DE0uBzgfi5
t2jB28UWjP4IPXTTxgSqQZK7GME/EeUAbkwRAPb2Vf+BXTwMi5e5P32olh2aGBEM
7AlvFHsfqk4RtXCJbXeh4dDBnV/bzu7rYQCsViU5KFS5dr7h++PYxUcaTye8poon
EOMP/bZKx2bUrY+CeODJzopoxCKUekU8IRIOnXovKK6f3RD5lA9bBDB1qcZhVBqA
+VS1kab9SuqwyF95NR6aI29FygiKYX3iWdZhl2DG58PyhSppW4ZA8ytmHMS4+iSu
cF6prlJKDbE8qz9RKyuK2fmQflPc99h7wYfLTre/Co6Mfx8saz3qUoqcmxAoYnzM
HQsUVe4qF6a7uos4bq2DQcHX5y6YktviDuZVtWUoQSaTMbqmbfezELQgD8vTBark
i48MiaW4OP2G9WPg+9f3jruzgSlEy6FZs7JZtFK40emfPlpkGNo8rSnuFDjqIPTX
KmrY4vegMhK+oDkhBB140z7UQQmxujLUH18MWuSnxuJZAbNPAy/NIee4vRYd+MQm
2eAI8UhFBrgOQYzkYrNtOpGZEzd9DfDyxwkf1DlvGAUlC7M/nXiHkDDHDWIdQTFX
4M62VjcA7cY7xKiBTIH89d0EjBFz90a2tqaZjHmlCON/OgwKUALBGilrn/mZ7fMN
gEjUq4hHOy8oYEEDrSfSxWxD4RpftCVIPrMg9DAnCNyAg/1hIgRsAFmJqKMN1621
1roYmLcFmEDD53iVbMbkinEQn14FeOjrUK7vueSD8TMcMPfo4cAeYR4KOAEnvRGI
chLN4E8E9VUfEDwebBKsB8FikEssXGDfixxdxjkGSJtM+jUR9cL8tGmBHnI88jYE
6nKeQ5nmfeFORW36Z5zrdDx/LVHHPOldD7v8frnvn73KoFmayaZGigjBvIGgXZMl
lZjdDhHKzPao+oYzfkG8I2AgoZyrZ0rgyUmcy90bQtNX18Wg9+nGBGFx59dpIBCJ
hj/3S2v4DEz2hhd5o/WZWPyN1wd8H3XgzfLYqxPQzBHGHwvruR1/GdEhDnm/L3iu
JMICsRrWkdch6Hdbiabfut0czbvchGTqSI0Jxtyc/5zTFRKsVVeJEdsyMig06hKF
o+/dFsJXDG0bZFOxcgZNTlM3WZOsXaP5bC3StQ8el4ebv1Ggfojut0aXezRNGK6Q
WlvVtiqEEBNnJnNw2Ztw+LVp00n3D7lAE4bsuc6w81fmJtmOiKA69M9vG+XV7blC
X7ABsb+4rBOnnKDGKMo5+kS+3dQ5eG5HG6POIZKzxvJXtE7fJhuzTvPjUOW2oQQo
3/5YRDmA+vhMjc0Y0pxtwPp7EMw04HRCUaMC0cjTLAel5ZdU1Y/NwoCAbK0hJVHP
9w7/LGVrvPDd78c2Nexkn+9Mm4UFHT0lSOqyXoyOkgw8MflSLuTR0d9AKT6y9tBU
Gxv+kyYBtBTrqIrKeD3xm/yE85xXh4Z3ZgyPPv3DqCzD1dzwe/O34R7DfFF7kWnW
934fJLx6SY9DFMEpdUTXrUvm857/HhMf0tOMgKga3Cz+p0d+Rd/2h55yUQNCtMtZ
zlY3oLL0Y81kQDBXFIK/C5MGWer70YpEO6ESa05jrFcQ3ijty5tMt3GreigoBw+U
bcah73moYVVTtN0g9e4Vacv97BZjomzneClJVRKCoWLdTXLqHEnNbUo6BE1nCfQA
yz9Wsk6Ioj82xklfCrDiznRbZCx5x4CH2c9LoX9FyDltg0weKRZytGo4mEbco2p6
nZdbebM/75NgdCFX9GoViot8WOJIrvE5GRHFFnEpLSbXW5fyuySQxtf7K0Idzegt
MofSQJAwz+MqFDyoub7rn+pyesdc8jfJlCyuKzR640XnmtSrzbpXeEcsuBHsqSqe
L2xVFzDmZUJm8lTHZUC1N20Hpz+hiuaqHFbeQM4XBzmyzlJ+gApZcndzjw8174Tu
Xy0tz+tyIM1+9q7g8Q3vpZlHxOyuNf9n/zu/jho54k6N+gRj/KNKgem0pPlXiOje
pt5B4YtGnFBUZXwwvuVMMevUlnZDLTubG78lcDKIAUt7QUzZzrzp0pE4P7EB7nM2
FXF+YODoHgg/0J33wQGXE4ryes8yAmHOeQg88B4mhfwASLjkflBciiZEpJOuDwLZ
0OeRO0joH7Ndzqf5bbzxR/r4/fuiAkJcnw59K/P/8xt//asyu6Ibx8jl6UDpSlDW
ZSBIisFY24IKUO+dk68ntjnc6W5xsvB5/ajyI3xnijzZd7D7AbU46i2gAXJEWOt5
h1zZdROg4VKYCKKwp6cFH7QfKnsQJAt/bgUyqaUeDBxTuCyr2Rw1lBTBMrnxWyOR
hrORmWP+F0vwnWRWa92JSpGce9tlbDtdaQhtUNgYeuxN95vwHhH2ZhIbsXHzcH8u
+aNlDINjZwHPN3coMWnMP/NGKg6knJU+TvkAt/FWN9PLkSTvM1TlqW7uymV5TYnD
9KaKeJjAgtGILCXLixhkBDReKryKNI1cOaMUzQDoLS00W4dciGwzHamtH00w0EJv
kbW+J44yyvFRQV+5Rfwliy1jq5/LGcFXkCxcZbDwwyCr9zg8/TbZEQpjAjOnQmBH
xatREJ3276VR9SCbDaEn4kPNdmi6L28PXoCdxAsDnm4JMVgy365YFqXencWWPW4y
RDhFVQr7VDIfshIUMTnr3ASvRxnsea/OseIZnYvKxy4z8vSLpng56L56o7SRwYA3
NDrqOmnnMUN7tAtETHkux1A9+t92pIbAQied2dQCeOUjA4Yi7UOdgajxIJv4SQUG
jKxO3JBy9qKm8ah45Ybe4a2lIIZdLVKjpSSgWocoGaw70TlknksYda4w0hNLD/5g
EZUhGo4LEnlwfuxfWP/ZQyPm5H5YwtNmyAJT2rO/dRoVdoAZh1bLJS8l3+B63YTY
2FM+55dwWIUP3E51ZkpTMY20JMwpT4Ewc5A7yGsT7JYUyuZGwOsTDZ9UoVy1QelY
wRk3RqyDl6bLq+vaeqjzxEgtXblhexi2ccsYDz0U7YA60aYmGPdEpm4OgB2Yb4ud
77kb93nxgadk0jck7HLk/6LpsSYmtm4Poh757GDUZo4VzDJDaJpbCNSxd4faubK7
ncSuyDOeIurOy1L/0cdS67Tv8et+z2gtV9xpzlY4udaoNdGtzpGjcexawYbTQm3/
xTCtZvXRQAleKVpFu0vCZFNuuYku40EF5ivTKPVvvcUzkwzUf9YduM4a10fazf2O
3//AAG63I+a7myeyiuWBxeS5K4iGieCBK8xCITyBd+S9HBWicbyTRjHiFPSQWBbC
Rhy2GH7yZaiDfrrwpAVX4dy7gFlRMMIzE7jAkWFhE0yPSs+H63JLEFcJ/w2vwvqP
og/8zt02WYETwOrCX4vaXtoGRaA3r7kbpZSvEZRPO44d+ruJdg/ndFjfE3Cz7S3V
hOWDwm6XqwhYx/9EzDYO6mYGgQkVr1w9P6qkgLf1FT7lGY1aCh/8SD7ZHwy1yJmL
Sk5HwHulrd5cI6ygG7Lm274rkjriXcAcR2IShwOGh6DT05AEf/CvkJlsS7hawqYQ
Ok0YDrOXRzPCsIOhypi+W3vTWzGdn+tqg/4dFN2/TB8fc2UK7fsoPvxbPInGEvPD
Px7m7JtNVdBWcaGk0SQsSYcTeVFz+V2Q/8Tm+6mEPDmNrLjjMYuQJY6Rg+UdjZNq
Oaj2CQ7gh1aSiUI5k6P63Q9XLvjF0+w3Y0jtjfMxjL4FREcU2GLeWEtYnbLAdkNU
gW4xS18BaN0+jREjGX3ujCYYxsC4b8DKHxU11W/SgC2nmIPhj6TTG/CnPEwRea9r
hiZKGntN4ZjItPfCUqsX+o2FD1HFqxU2zouk6p9WjMUFey364K2r2Ltv4TuDMNGk
q/OnuIQ+7UD08c4BbQe9wqdHaGPRtu19fcBKWZf3FxGX4OPICvIQSZUqCan/r3Zh
/VN9bIwVB5GqLgOjBrg8ke/vIXGHCjfHqI1VD5cVr28xrogB1nrii4z7D8FuOAT9
Id+Pa5WPXkhTWE25WLx45On0q4xeLp6aFFNunTZMQPKr5gCMymjBMbcIt4jhaAM1
QRYlm5BNtDJfzy6/G/EC0mupWQ3MkVu5GeEo5G50ARmOfMIg3GqGtcwiDkZ1Wy1G
V+L8pqxE9qjjWpnNoVpgFQHVy0zcZWhAw0CxpS25oGqLTXUruucz+gDtLOhuovRj
pU1FRUr3uC65wBwVf9MG4YhwDdaYCc9PhhEg0gtVtTW2HMH2pvbe5OXzY6VYrtq8
RwISR09E3ixqHAqdg+FKfe4uxfYuT1eHlLQRtxLNSoLlbfuT7v5L21LInR5x5ZQp
5lXY9SP0Y+MJMQA5PrVz+R2vUj/uT3H99cmcSRxuDVRLCpKQq9vdXKCirbwuHDRb
KVvJTb8oCxY30gw9ey6mIKe0YbLI/ACcJpp8v8BkgHOB76RRdDoHrmCKoxvg2H1y
lqtUCGoG1LKEIDESvI+u0d/uethxztFI50BJ7m+OvDzcrhDVzqvdZlwwbp4GiDAD
jCZ/ngwlhLQeupHWADr3qYJFHbhTPuPThbDyVvbyIES/n0RY0OAgiGeId+pklaJz
PamB1nVrlXGudXSda52+kJxe+ZTmsNIzcRS3aEaO5z4XnpWz+nxfcWiOuayHkU/I
fMDj+rkPEXXQrj5+DDfZlJR3Dd8+p3f0Y1gumSP/AWR/PCX+iIfOov/WvnEO1Ud1
+O2VbQx8yrPp4wFt+Jfnl0jueW5kZW+h0D0LgmhNoAtTD3szYWR8iTVlIo6uVNEd
cBHmbCJLQDvG1aWwkKzN0A5nG8xirvYc1WkN0JrNOeWiNXMA3n/n2SNtIJHco5k+
l7hgSHKhiLLdp+lDbQGrIg3qNXVaxFH9Chp+dwGysTBRTDVcRv7HqfSk+UJNaVEB
7e97mR6pBg23seRDcL6gfnHKcQcApOLYzD1DGpdRcyB7RvkJSC+C/JBHIGhLAjf8
Tm/RX8u6lOZNp5Zreg21oYf0hW2sEjb34cQaer/8x2Pfr91IaTb6Td19Kmwf8V4X
Bpy6HaqPuJ+fcnfK3wHm2q10YYAHwr61tMFel3QAkJJXMMYBocRYKYwFQ+DxsNgW
2fRSrfw0iAcpD63h7tir2+fACFyOensIenaxxfz6AJ9/bpDGzKIXvnXnwDLdeWN2
LWP2M5T5s0dJbzsQRKY4QwA7G5TsL1QGTk/gnNFhIfFFA43NkkabFWSF2Q+5xoGN
xV618xkTsfOlobGuP9yGtR3lymwbStJD1wPvKa/BFVAEefZtBVIg2K/W+xABZAHK
YnR7jyFxb8e1Z4ZAwt8NcXcaVGJ028pYEyo9kmwkwLKsuZXJjZLoIfdeG3clcV3K
wqL/3U3LcXAOSU87A8vVwu6Z04TDmjbbGLuVfyXKhnY4B2dIFafin8+rqmgU377/
CEq2Zc193XjXdyGc7C7HpiAz7j0AVhPhFTPTlDTFZOEziE7QGRzjIOq4aNyCMgIN
fnEifzdFyyA2A5JorGOTlqUzhu2vhEyP6YCyWn5pVoG4e1ViXJKHJfsPh3PGaPiv
HWvtXUXOZB7FZKJ3zv45f7OyzsW2Qq/RpuYGjT49xiPrf1q+xbjzNPc6c8FOSqyq
j1Y2OC8vkVCL6CJRDltw4aERvmR0UTx8At/c5ET3+QYGPjxAa781nC+YGHi7wOz/
ht+hAhuJtYGv4+D7WrzHGVQANHMX3rpN5jnvNefLXbwNAnfkoje9165GR6uYc6xO
z69vGrna9rIjKZWNspevctyA++5L8VTU79Hw9QcFMraoCd0iYiudxRcwQz2bbVIj
4S7fvF7P9GCcX7MbG+M529xaqNay0p3GkqOHEZnP+rcFWffNVnml3Ef8T0w4LnbM
3/G6x2IjwMb+kIKnyFLy5OncbW4Y5SzwW1CqSZw/DG4T2FhC1LFb4637rLJ7rQiF
cVyrPnEcW+yX1pLqQ41eMa+hUtCkqSuB1f2iThgc1qwWHVBy6gpofkgIffv5rMS4
3u2lZOi5VnvNhRKmL7YT/E19zC3D5umt7s4E+VN7CpjXmgCawXDE92xiwthnK4gM
6oSrgn7HLZ+b0SvjiRCZdrpKuOGKOxWzjDbjJhsC/veV9WoiEd8LEDOVOPPvbYUQ
6HHWeJpzjD+Kon7L5U/dm8fcTfu6g9uWPIrDyXC5UIQXRE/f0u2rCWcZXsnRwu28
1RXJeJFNefcs0ZCnh8Ngl5urmJm9HDLFz2cfTknOhXnkKEUyXLjP7qsnlt427/He
jZ9Q6zfEzjNJXFfqlja5Kngo4a44nIJga+YS8Ti0Cn6yG6iYk0wj89Q8QF51Fuic
vB+pLyYPG/Ge5CWwTBguo71MFt+/UZQXqk93acHe14ZKowOHI87t62Osw7G4wyWo
g/4NWIVDIXRZFlUzCe4vYjWMExCH+N0XVbMyttd0X5Gr5WvlY27jOtYVeemPZ+l7
qkYPsSuYxPCo6O5oTqrdATvQ9zqz+3F8vcUM2jS+9Nf3H4Vi8+tu6HnhmnPo4TSi
pBqSxP0IfcE7dN8K0akFQfARDxMMHLMI0NVyvIoofkgkD+I82C01El0gmXIths38
1C0mp3QS9NYaQlATQsQ2+aAp4HF3oq2+f9R9uxPJzfU8aDABHwDH+YLBHOXS1z3C
4A8Ym1mapO++L26+/AT7hgRCYj5RdJyZbEZKqEzuufRcQdTmSrFjIRQKn9iW1dU1
gUUKMJCPQB0YSav9DZbBTINOPDKdbNobSZBbzbqWscggQ0D3ecmXTbBO5iff6dbp
RndyEIRr4ydXkN6sd8kiYbidF45Wg9/le9I1KMPlFBZlDOuivNmcwiFUybOE9OOW
baQntl0MMGeaTrWwbduqTzGjqRITdRoFKFOCYaNm2m/1jnzrCAy7S2NfRuN1H63E
xPRnNqvV0MQgGPg/8dtYKEVPPvWzXWPHSynfY5Nxod9S7oeVOZcaUwPHbkLkxqei
YpCoaHLx60+VTGrQkvDUUk1fs3HdK04oY/NoB9xB9+pDxLy9Phnf7uITHbhu4O+l
6NjOkHlMlqKiHUf3O4GxwyHrYIiD4K7PJi8Y7ZM5x7Md1OcLw8AmXzB+YcTExDIg
RbiwPt6l61I5Bbvsh5PXCVa8gLQRmEtBSrbS4IG6GjjCo9hB5j0RCoWlLZdKcbDU
0R+Al4wTHIet1TfYvMxAP2XcMa87+l6wMW+L1i+sHQWIb59btPZQGrIktuswRTxJ
27CtMMOpTHuYFeRjVLa/Bfocr+az9MR2OUKLGahSpQDuiCZ7d3MxLkTLUyogIvoy
31SErcaiOUmSTMG3c01m30v20cceoDyXbDyDzZ8BShCyMICQvg6CBAOuYeI3RHAM
1yu1OvuSNH/Lgu4ik+qrnbJFx/XVlm4sUfEUOaKX1TRMMrUxSbbfp6mn1+rkUTVq
E3LrdhC5/0L/yKFSSo3M+XHD9sEe607kSrlW4fiw6VAmk1Whl+okmfoqdYDsz7ux
qhKUpmz9Lu+Ou/djxc0HIN0PEmhyeT+OsEjLQqwO4IoEIifIIpDnuZU2OFE2swxx
dAgCRCzX9lhXE3UYJHgOi5TQQaSsgKwU8iRE1+sNGMbySu1/9YHMrSrweQnb8gEh
jq8LZuZe9x8pP/rNUpkipmO5uDSJ3EiNJ0TWyF9YhW+jQ+h5UFeqqahSJhYgoZ5D
o+o8O3AZTboQUbCx3RmsnbI0g0+T+OB75Dw2k9ZdFH7/6Bv3HUVLh9BBUEnLNxPV
wulOzKa5XEge0XM4ulPc7bkJAR5g/uc8NVNgIw/SAM0gzuDr2Bf0VtvLFQb7cKhk
GuEdQZnP/G3Ut7wlZTt5PeyYYiuhEgUYSB7TVY/umRtKbOldnBSgZ3qjHrN98RFV
yDi5u4/PdkXgEmgJpNKo2dQZNxqTn6uR7UJgiM2/WkmDGtwI7WFa+kSIJmwG+VbV
YBYhArrqdpgxDzmHparKJr8CCJj1/hwmE7WtKtc8wGUGv0xmBuXbmAcujw2S+MC4
zwcsIx0gHoEPAfzRtLuRwbSbsS3gJL9a+cPa7cNlttqyQvfNndmkhJWI6EWSqKb2
t7q0ESjRdevNwFc7PMYAxt77wYvybNBFiMJViSqyynKE/+iGAyp2QcPZ4ykj8IOw
jFeZn3xIMXX+tMBFjyE7FmFLJpO8m/Q8bVip77JEqyeBzX46RSD6GeA0demG4mOu
qysY1nu2y8q0291GK0zpsXoz4PnwmiThWNZcICn1+aPRYtOqW090tcgy8s9Tmvpq
E4ysl8LXruBc049RpX2Ku100RRHTxgh+iWoLj9gFgBOaH/oPAV6Bs5ogqNZe8A4c
JvMaPbGUcWr7s8DHDC7Fy+xYNMdxp0L4PE0H5j813YHPdcQvjN8ygnYuXkO11o9j
/QzqTUrPVhY4WxQ6msCtqvIuNcXLuh2nQnje4bEfAkg4fxatqLsmONBtY5bbbQ4+
T256aEGZfxiTQgJ2i61jUB3UlrXQKytqZ0hllWn5cCDsEwaJaxm42T2ESL17fPie
/JrmbXT2SfG5kCSBp0CLASBY2yqAwT1UMbEIm39YIOGYaRF3TOAFPHUWaAeuI6Zz
9WD+VQBOlIlcv4PgYjsV/j6npQx18miWJtaG8gvEXOmh5l1nka0PVuKM1oGP+7Ha
CvbZlDF9p9hcn9ZZieUH4lK1EnPj9EQ8L8x6mAbsvKtPx4p5CQNav4Ze+AeLnGx8
8JMvWo6CujF/9iFwHmeDJ/LrYWYnM+REEJiI4s5JMgo5RluPlLqUe0ixhkVDvd0Z
GCt2Jm48pct7CvvcqZqBZl3LDEy5d6/+XHzkkfuFArhFpt9jfljvMv80aaZmglB4
GbZiR9z6M0BYDJTeZvBsA6uRmQJWU2RtKgWhH9sud4ugiNukznp04MhUnA3ApbM5
mTDZshC8b8CxuM0k6P36MSDUTW5FxzXUysTkX036iFHePd6ohJyNjM/LZJc3/U9J
o2DUF9yMlBTbu9Mz0RIp2WkrxzhW66T7v/cQ5h9tju+u0B9tXPsiqK9UcWh+iak+
N32qm42lbKF7tgbb4yzYvpLO5DZSvkjSiJc2a6VExh1MxyabNL7HDvkkHq8p0NOE
hxfBjKC4jPvo3HFN2NcJNKgyMJOcPxXvcJAO/sGYddZK7LfcV4BzZRTXsHjzZhck
QMnjzX1JOjMaWh8Npbm/k550WnkSPhUPq3yItHF1MZbhchX6YXpFpuJ67ESQ9fMz
BWeDhJszMqQDUhRuv6pGCa4wo+nwcq+AfdAKnHsi2dMPKDt+daHOCfKHmxMlv9VS
FmjbEra420SYa58gzHh2Lu+uTHSSXpC/MGXr8jdz4MVQ41VXiswUBWAFH2uZT4pG
cJaUdTRCfNZZPBHIXYL0uivEIoK+5lZrDQFW9s+dGkc+zBG6uq78JmBnyi9p9dt1
3LXFF28QKMZZGpZKgUkNYulWUkIilSEBU8po+8ds2xdWkSiP3sXd2Vz/9LLPmK54
pK2R6/c0Dqmu5pscrg9900E5efIyTlGEgmMB2TMMQfZnexbY6QK6MsoWyOkj6IRx
Rdz8zLfr2RNeLc0RJP7ojgjvHkX//f1iQuo4fxjA6FruBGtdOIJDUpUVlSjLQcxh
YOxFldsqZegFUOg4kdmKV+EPRtink0ouIdMMAWj9T4cRsaXpivx1yr0n+mps/PQk
wqHvJMO7g+8WCJVUy5/UjK1lDoRW7X0wcq3GQIFJvTi5z85HidG9WILPe6bW28Ln
L4kD2ZkyyyqSBvnssENqzPhnWMgX99JGoe2bVgKEOttj7IlAs21axzen0OROKDUF
oKgpa5W4k3vi6DluuAUIH44HzGkwRAgsw7vj5zuHApEMrWRF8RCT43uaZgEHd8Qf
nj5yno3YDCmRU6Phic/zD07w3RBgOcjSGXcgBbq/HSI3HGoXulOqLL/MDT/I1ezx
DDH4ma+t+ufe8poV/YJOGSX7Qo/cMsfdP+qjYCF+v5cTz27BQjiGkDApsPOSqaMn
iGG+uG3sAAlbZtpMzglQSrsYQW8vCzsuEmCuxpAu0FWCqFz0ykDhOYRQHDdiVRvg
7ucCCEB+aT6jV984LYhcNPES4ShVe2/YZN5RN6C7vbpt/HGA4Rs/ZLN4Wa9+N71H
EgFCalLc6dxS0i9/+iQBYxy3dZ30fROdiSlNOo1IAwmLoFkcuH7aAtbILS261wiK
4GGaHpjQb/RJ5GQ7HzUL/iAbw7Fs9iNhTRSF7oKjufCY/n8njOTwCKnXpSk6puJL
sfRNZnQPAzX+hl/F7GhWCpc1BWmiiD2VxCVDfAopB/McmnTQ6GmLYa34ahDH+9OY
m1pOTDbJ+KO7Ag0gN16lP40bgrf6jZ9ZG9SkH7jtywNlfze4S8hTZKO41vmTObIo
4UPSoy9WMYY+92Uonn27Kb9Q9wTrVpKEpSiREnT/XgoEv708rvJwORq6S4LQs+GE
UnIb419gnw5yKLlfweGcACVNEj8m+KvUKU/Ug5XRdkUSn8neUNNdfPRkbeZdLEgJ
SPM7hHmzMGVEQQUJUTGV6E6MX2rNxUoKhGH8eXvaGUUnTx6N4qSK617/BXLaKIwt
3DM0Y+jt1riHAZMF8NNx2K+eawxh7CfsRZSC823zONNLXf4eq6yV4hkeX3QcvSaU
Cgbl69zJkbQlxuZFECr/GAazv3No6yK1vzEjCYqQCAtUUUVWzzt9PRZOsnuZvlfT
X7IV7uFf4wBb0kAn00L1Z7xW6WHoLZZ2oHtrMWsmUr/aP831GZ1+X6qidT9EzgpH
xfaBP6A1f4bQ9VNWMRuG11zn5mL/cq0ZGWNHJe8ChxrapXFgtKA4UWLpkXgQQWv7
ZGZTwAi0T2bLVImoqh6KG0M01rXTsE3DiWmTiIyuhVjcXNm3urQvSxCtDLlABOhq
MCSvlNdaK1VJkUQ24XT+VMIIOg4rtN8+bQU//D+KbqX2Q4OK/NCJQG1EX+kObDJp
aioXqBtEBYSyIsU1+EWS/hnlOVHKYSUT+9AbiVO5G9Y9ohzYZ1GWb0WnOEx+cHtE
jWCbWERH7RG+XY1/y0eCt4ubR/6p5vJgQH0Hm5Ih8r3fT/Tl5oPK8JIdaC2ld5YL
55/CqyAj7P5PNER1qePoL6VMFvu8lwFMPoixhgdh3j55bco/6i69AD9Yaq4SfjwW
CocGFlBK6L8AQDmeggDbCqvCGaufN7Oo7GjEmwiwe775nnWaZ70IeIT2L8rDrIT9
HcEE7Fxp7+zTa3gQKfdTAWTVbiTqR5o8MrqmnVPaDvlnNp5yrW7Znh9Bx4APBx8o
KgMIJ+cUbzmHhiOFGYYt6GMw7TLZ6C3tM0i5T3kFG7wgwK4QIHrfAUoNjk4BB5lL
ObUUjuSTiO+IBl2jCX88GUFqI+o0Z7Pm8VcEW+rb411NUyeQvoyhfzwsak81iH6J
WxEIZi5dUITLNu/WHT0JCrltntrnWFvyBm4TjQ6F3yuJguT9ERaJGUx3kT0qHVyi
RlU5mfaskBCyR+GXYHBuyEu+yd34DARVkhic4fc6yNYhclu15hleccYcJY0wbFDG
6/MoWpSDM+sXjw+Ja/KWkPQjIBQ2UzuHHBcpmeSyJ2LjDSXkH9MsJc3ERYDi7T7E
gPXsFuV8N0j8nFYMYGdKA72Uuez1XJys2UmmIIuS42uWYmaqRyUgRossAHWSdvAt
t071v3jCi1depDjhSC4mCtonSqyktg033W3seEOALCbNPPdz05n9c804gl+ABr8f
ruMoV0cJPY+DWhZwnbdtzUlY0D8VLrlk0ZDZIk4DvhjabXkkI1EWdSVUvVCZOEnt
1M8/CZ/uOe0WXN1pw156loKeUVKL4wVEl6htIGsbC252KovVktbN6bCLNQEXefMs
nnmhVMahmQ8Z3yUV8Uq5GBzVWAKuj/9bY67S1MWRx8pNrBlfogFKDh3uzbHvqyYq
QnCRT4RfOweTeges1nTq389Tj2ORftnzCmscXX0EP+O0ikPU8aUe8bg2mr/JCzIA
N0ItC/Yqgw85wLvad978nLrokSwmGTTjdMXxxbOIC8dCp3cZROwqNIYvWjee2nA+
0GYXut0nDSioBJSADrE5YfHK7U1EwAsj+CThfkAtv13DmCmWHoJx0sm7eqiiL0Vz
VO9/+I7dJQ9613QWxjx8kR0TQt5sXD7pCMp1HxXxOmCp0ka4FfO/FTOn6+j4Nmb0
vPm/5E0yRdf6YpzHxtanoN9pfFDt0u7Z7ZobWT3UUZ7SJ6u+KTfAmJn8nJoUqXmy
kh46ZGpYv4eqBGUcMh0fQlz7DmPTwytSi+sSF4PMV4cOuzUNHhlB5M14G0K0FEHb
Te1SzBk0gZJhL8ghSBR5cOUMNvTpOW9UmJAXxeW3j37u0KjHuaGKIKhj7UxLv/LE
/8rMKbY2BDj6OCWOUSicc1Gks6osLVHEo5K+j+GBzh4Z+SumzYI98NIJ0o7miAar
cOm8HMK7Y2eorxrsn7DubU2a3p8ReQ7327sY8JdcJ0IQUG0pXLpK+dhBeQtQBDrV
XkBnPvQrH3MiHC+wIa1AfsoyOSoAEeu//q+B8A8XtFxzsLPk0yjDyTj5A2i57foN
1GHMhU3W3JRm7znsbhdmtTa79d9cUu/Oi3rAovSGz1eMXkW9HfhPUxxtqe8+WT5B
Q2giKrx8b7kskL7IQFcrmoyDQwIRpj/k7vdWqXR3x28GVCZKZ2RbcDK7dZoc9MOR
edjnLP64ei7GlEM0l5jq7kjw3qGN0XdqFyDsDxx8a/JDbqFUHvRixaaXViFDx8xw
rcWDJKob8kNSSEsvILbxYBDE+mNRgT7a7PgVf9bhPeEzRYYC0SDTbZJzMUpzH0/+
K1M9pDACBhC7EeXNY0EhxOYSu3v6bPjI85zDzcCP0xpnky04wl/4BpwgUgwXXgYv
63dNliznzn2ltzxPJKO14S4sq+pgvcR2pOUFHKDRumqzlKveCMYV8W0+Ov+0fTa6
Cq3HYwf8qdF6qg3ifpI6Ik8xD9o5xYoyXRySdAWOoXNVtzLBHODP6THDvH7bzwU0
/wFRdXyJtoPkUh87A1oVvNH0+rjGF+6g+nlNlRxNqW6BxiQV8jJ1mtn3KSLgGKG1
9pJiNFuqZiGurF7Oz2ysNRRJGGNNJbpKf8mu44+qYF/7SVqIMPBO23vsdCUPHs3e
ITOv5x3Dl9TfdNHdMNz0XZoMHzkmOAHs7zB/pfHjpGEQCYRb1TSE7k8n1NAp3boM
c786DK53bT1sd7Rch8GbZjqtG1Ryyyh9OXIELDLpBJ4clv+3L3Uiqm3b5Gc9a0xb
qfugu1gocE59liLnvmSo9dWoN46rucZR0FVM2DeIyBPWuPy6dYlN8yOL75vRMfT7
Q+uc1sdWuurERtHR6Nhad2Ym3+t1DEPuACkZYUhy1D5cLLJHofsgQiihZwPEeDhN
XHSIcsWLZ2MWzUU3e9R2D+vyjHMvzxDdximN86AK56saZ8c3Se45PlqGOSxZgG31
9zwTpYcTcsj4LrD8m8TQpKKNflxBo6etCaMgbvxAhP4LQzjIctSyKikcfDlKdQ9Y
YgCwQDMJIBwbyXg1elO19Fm3gPOJLal61+O5qcWar7PoDGPwnZ8476LFcrEpny5k
WN4s2+miGZ/wmxyHnIp53tZsf46lF2w/S4eCKewudauD8pF3t70f57QRFWsZd7UD
K/RNwh+yRmabZ0/jpjY3Hs4BbwMYWKKbUhxRkXXYP2oGXFwRbktJ4uBW1s35OxdH
vqfUWQjF9U+sx9Id+gxl9+c07zPwI5mLAOsp1n2eZm7ztgtnPigRkEk9+z0OLyBb
uLHSi3V8JTLxrD6VloV//g9wPfOYxQYp4SsdMYYwUaJ98AUp15hiQHvp5EsOfmBh
VBfOLzHz6NXQgxOrb65eZkVHTPoAdTYe9oxfWqaJ7Y+p/oM7s+fD7P6Q07LDfGcd
mPa9JWGRRf5pzQkFg4kGeg6XryowtnjlI3cYP/vxz5zziEEIMSumi239BJSswP7U
x5AcH6m1YP3bIAipLuWI3Aze0k9MnVh26Cn8qPx67Fk7A/7abUGkpIGFoHdf4JGV
hQUadBYPMDFDSDrfpvWp7hFlbFavKRdjAA1d1iDQEZErcEIaJdliGTdByFTp4wzA
50WNoVlKyktuzWApol9p3ricUm5pMBH593rCdTo9RECCAWQN/CfK15/NS1+kKmbw
czbxhRcuiGceKwjAegJOZhI873x4ZLgQm2DwNN+iut0VwGlM6YAg/q29oBNN/IhV
1fwhox4g3bPdYXP60rZE1gLVC1DytHBIzYx8Uml3nDnUSTN9QIPGDGVdaT63w+lM
9C5b4sCPpiiavsZcwyEmykQ/aCEFYAj7OsiEJNUp49aFbzXpg8tlm2UQ7YlvmxG0
+T0dGs8+U8DSdBDgqxMKQfyUjF/7QmZgtN9dEhSQQIjmPgIcgyD05Vm9+QKh1TkY
ZA9Xa7hClohLHRLZDzzv8jnU5ZCy8QLHF+yMLLDT2DRp9QxtTULyvZMxdkEz6g4D
0N18YxDoJma0wPslavYNgaODBF1rpvwO0Lk4cLFgXh4cJuptTOAGMK2tX7um58UL
gdj6KUQoqnz4WX3GpSM6GV7KaYHpME+3ME+iIxcVfOG79Y76S0xHEiwXChXXUQY2
5aDcvqZVLig2d36fVztnodI8dVsnOwlzJBaLMPdRkxjDtQUx60S0vJ+17Mvb1LGJ
W7eLMA7Dh7FSNOvhVtKe3iQHYQYDa5eYTYlPtVmfjm4Y3TmTLf8LVKnmhh19DGgt
RGODyWVoF+OQsmE9+Izpo4TrvZVr2GNHujDUo98iySSSB6DFqz14b3rSXv3/bTDA
oP/nUv9V0DUmJPt+eSFBOWEq6e2+8PpMsdIXA/uhtfxW/XipDQdZpR2VyHXR3FRB
MU2s5mwIFNxjsNzFB2y6vwGPnSf56x3WGfWzCn/x/3AeYwnehq05LIfUZDGRBqmL
PIynq6lKxZt19ARAH+b29Wyj6K5xdLf+pXiiRnK2m5XwLDhANhN0eGtR8WjZCOJa
IB0GQvrfP3ELDq/eU5aLHaPED7Y93g7C6eArg724d1BUll8LuC6w4ZIwSDTarI+4
eOiUa9YgahCYVvLWESElBFSaY9riBxQQ+uQK5rjYiD51owaU3PWhPTnD7PRRfhuM
Dg+cV2lorq5XbxM+npi8FEBr/e3Ea5VlwEeOpFF8dBgwYO4OsbHaL5VY9lz6JnSW
R4YIhj1lIok/WltZ8/C7E0pFdv2v7U91dd944Z1rPF8/e+hquv6LAB1kNohXjpOx
/DfuDbsZGYI+pbg+gs0br6iejxDQTnA4weyiP5hGTie1H5FIpJ4fNxFrDdi/awO3
l0PRL6tyXKBH1NsxkwIsWQ63CfvNfDeAjXcy5v5AkhrwRAmtd2FL3+eigs2IQpZ+
FVS8xvYUq4AHsC99th8Nvmz0begJmluCn3QoZhmpL+bJHJlyy/wSK8P8rYVUmhUv
2etNC+awUD3g/VZrNkYA/OUMzFwJ/nO9vSOTIbaGtRJgBg3JTPL1UGqrfLAQIKyq
VmCgVCWMB+l+vu+D3NuVyCjn+gHndpoSZR+oOuq+KqdJFkhqYfm/I707dfiLHTKO
EDNfQCiIXfsVCE/uQ3cO0zP+Tl/Z1WVdSLw47NI4RKeTtulAEdZyeZExgTMyB56x
f5P0w3TEawWFMlxa0vY48Bbk4PyARHasByIU+hpNLdbQhpsNCwNUr/qWn9p6yI43
aZC0UUQcBDKBhB7HLIorcfimKudUxg3kGLqey6d4e0k/1jsHdXDdUciINXi6TH9Z
0nt6ZbmFWJBzrWSnXTiZ56L8v0qlVwtIkflXcJoXSK03GTiz+gnW40wHpsYYwEXH
7IPmh2iXncOgIlww23GAM9XNLaLsQlHyMUzyMIqTyKuLZcVWRI7oQNK83C7j9cx8
W4Pdxek+8tJ7R0NTavtBPDU1pgUDTRUBkVw1OLq+l7cDMiAe4hW/xrL2hxqG5/6P
ipcman/VL1KMg41pMtNUYuoYG0lVj9s1QV/0C8A0cgrusJjLX1iHPqdC5CAkpKva
wi8r5UOQMyXgHJKDpwxSKRq1rJDmYnpTMJNLrhGs1jjSZvfdLU2fBkr2rPAuls3C
3KkoUgTQoRC+YeuX0ZU3iREq2f8BmcrZ6RYeMPqwqbX2rur+OhKYEbyhfL28rg5m
Ic01Db9nWkNvUikDNBnI3MGolIkHb/wQbXUMOv0XzGibLv+Yc4/1oi+P+9DpkiCy
FvT7hE3Y7zthgCta1GlBpGGNeLU0ObXKMPgKF5UldYR/r3VFDvGgEg1WdUflmDjo
IINDENu6T4iaP2PT6Z3yxfwUrxC0VbXc6/9lO2+UEYfEUVyj4evpiW92rP41RFGr
MtW0noNseMDXWllgLfJmdUFKWfUj1xcvuDy2wo/L4o2FFF4WedMPe4wZmslFqEvI
KkIGyDKGXD+vG2yklxodcg60BlQoYINvgN93m19H/hkAxp6tF0zuVj2E6Rl84AZh
wPF23OxOjDKtOvU6EaVNQOYGUEc2jzW/t1PN2379qxnmfmVW9PhYMLNwG7OXKAh5
C+eg8dWwAAgmJ9fRLEz1CZrSemJbUInv2uNBteDUFLSVtWwJWRMhm0Xex9Cb95AP
zMhNl8B4xWVVh0JUweKXtrjoqlhTuqfPGdOGmsJMQLgTHyoRWNPcjFAsXdM2IU+j
BUbmHGY4SGtbnnxo5o+zoaCJspsrs3EB+psl4WuWinxQk4JnnytaL8LeA3Cmb5Aa
ovoUkeO8WfJ9LoMGKR82VzAE6NQgnT0xiqck74EJ5sy5TDUDHVXd/nihDN6jBwOY
UOM2W+HW+9hQrH02CQBGfG1r476Wp227bZqbEGQx0PR1i9OHhjS82apjdkCOu4SK
27c9tVq8SsXTvLof1Rrz4Ze0TOxeNiGGHv01BWMaX+hTUceIXY1rbc2Ta7behqw3
ChYM5SDWPf33WVpaxWEr/1IsSBVainMfM/SCcZEZQlXQ6mpoFdUgwOvD/WY+R3BL
ZcIe7GJ5/sF82/kMdmIiPaVGNFgBlNwWRZ+83VNhVzPxtI0yx9j/HOYdaAwhKdMW
4ljZSpE2LLo5PrLEYHBqUk6NaULcE1b770dBWb0mJjr+K9mwp+EOQlsUI9z//q0s
QPSJ6ofEQbMbVeoAkNF+HpwApBkeQLjoqLSsWrcEW0v5VhvtZIugqAzJQQ9NfNbX
xr5j7N0tnUD4jYcr0RNk7GKkVGSW8zRLQLirAJM4eRn8b783l/oLsco8R9uqbIAX
k4kMY+1mO/xkFEyjVmPYohNzK4NAAxS44uC9d1zkWHLe5Fw5UIOlVtRzeVplkAZl
pJlROTYCQXTrO+dCTNYUGztNz5zjiIUpFEYWwnN1Hv7iTaAgYlItPrLe+gUiu6Zh
wctXHo77dOT6PHmYVyhV1SyWSZ394OFO/AFpXdHOc7JG8i3xrxk9iTpShgEvvnQx
soeKV2Mpm1HoOVxQzU8PDshn+8AkmGpPD83Lt4V7XT4FsJMa8p67oLYG3pZDDKpO
l0HqL7laKpMfPOF37Di644+9IRYURwlg/zHIa8ijPNzLOj5ZAcvDKI1RZFwqzN2C
oPG0z6s4Q88Obf8PsUvN/vwzJZ238CpYjmzcQ9kR4MgtneF9ykvOjT9E0HdtcegV
TSMBP2P2QN9U7XMlep3mA+7btFqqvx4Wq3dd0Bx8G+bgVuiM2Ku40BmBhL7Q0IRx
m1tYyYeZD2voAUDdB05iIvKsNv1j7wqvxuo+yTDlOqLI+2CpaObcUukJuHfQXNiW
7i6PJgBxxVyPy8xvK2VRc9VS420+TCa8WWvt2ljTmBiMP346IZv8HIfESK/IqDHP
lzLxtMcwHTkZWUVzx7o0oDnBK1FyQ80mZLVwwy8VbySJ1w5J0VyfHZFAhBgyRzOp
LvBYYj0Ephemiqmf+tOqeTw7CCHHsl2CPPhtw8SZt1WMxhBkb9S5Rnb6u+QYwH6T
JaTfxTZ5OeiimF/vKApGBP3fmhbKs+jhlXhdsOphgaffDt+qScWkcpa9L9iJlC4p
IC87rSXDroHGFM3tn800OiumF8WqPJCmWgL0U0U6mA9APwfHPsH9cXynPw16BigH
1IeBGMTO1YwiKU8jv01XwYyyWwZZJenKNPMeDBG9ul28BX5U/ZuSluy/rGPCOSLn
tDzvqRG9N+ROrKnMhDZ1fZ/e3+TC4/tl1q1mxFRHqXP2TQkula77H9xdnWbAysgg
MbNY0/ckNAimAUlzw5BkVELgFCLGyXGX2pq/gdGvymOaP46ZZ6/C34FYuouulpwx
LN3On+xuhlZJplKYPb2rrAlfOB0erMu1RVaZf6pKHxg1t8sB4e9NUNz+LHE+EnpU
vzdTy25M5GHEqYLmdFDjWut52FVZrbHhBAQRbzxbHybyk2WXtHOMkEPoi1lq++Xn
66qlS4H6kpAJ+lOsSRzYyZ6TzYhxVztB24FwhHGsf5Bbq1x9VkwL7WBvazMenLSY
hE5LW4JxBW4v00XyLEVc3Xm1nvpET0YJXW0kfZjm1Tgiqcc/7OfceUPJlXM9Lyfy
t+KCGqtNDKQ8uSX5pBdnCSJgym+pjgGtcaZpCaCYZsL6Sxv4E10xkhBNGvumikgF
pU1nNajpOF0vGLpXsdgy+mVPsiMbTUSBJjuMyFYOfF+CGFOXgwZfyT0vLLwfOGml
Ckcct6SjEfQhbOCaqOM4ckHBHoxWznwbK4w6/pU45IBR3e+cV6+8F18kRxlNU0Gx
dwImvsylRqhea+Ed3RYDloL2O32G6E+8keo4WnBSYl6dKNoG5ovTbjkJ2ryPVFfe
+aD5ebFfOCfawXYbFJ/Wee2/Szil5L0vdRbEsi1Aq1ST6YGm/fgo3TrdsT6rJ4F8
fBHvaCNdKNqed0Q/RE+6Iy54VCMiY8B9+40CrYU6mqHpU5ds3iKF5FQD2topi8lL
YmgT8DqDLa+EoFfT004grwKgYcPBxDqJEy3hbL2XB+Sqfb0NEOIv3864j3rg02vp
prfF1BCkyupEAUxRXcgb+huoUj1Y1cG/U5jyB5KNd+VXEhq3FitpCRXufR3NZxVT
m6bJEKq1aEVjpG4Ed+Y/j0yy+L/iJw3rwIrMWHsTZLWJteabk7JKugp2Hl2H47Dl
X6FrXllAhXobwK3YNmI0JDcfmfiHUhXZhnX3DpTWa7amOd5Tl33/qT6ZZQ62HolN
h94WMT4CQ14iXz+x/JYtTzs7496rypv/BPcyVoMe1LABsD3IcwHlxRlUc28X2PHv
VscZ1wSnk/6cSCbcb0Y2FheRCFm3Lza0YbIJH+MizrKvrPeweGeaFfGJzbKYXgGw
dp6xRmD5ARwiAOQGrTw/ENz+8YhP2Dgg8i+sZVxDyx3RDmERdAxRfaGIZ0GfzZc/
gSB6olaJRaQ0jrskmOthTEFjG/7RC5ZkL1oFQSd35mpb5z1bF0nc8uXy91ScNaq0
ZijHUScjWHuvJnSKW3+YiKX87GWkYunNeShhEgwFNIr+Ud9p2idRQE2snjIWw5T8
lcbwAnRd9bWJLKqSYHmiYMaV6RR82e+n8U6AqbJv8SFphrxwAr5q/vJ4xi3sTPnc
jEAo+3yo6wtilQ2+iIfoC9qfAYfQbtvXw4nBGEz6VmjYIlNoasGu/Fn8il3+xGse
nW0DYb22XSAPZaymZBKubwG/JMvoWrFsv3nAL4/NgW5OyRZeqUgf1B1AGniVmFy6
LVHFw36RvS77fNuXK9NfGeVw1EJAfr4bztUZf37kBVcfetexYl3UVbqCZLkIQpS2
kENyXpF6PJvXJjLhP/8ocEZnO+VTqYTI9Skbhe91H9D9b/n7uQECAgltDdP82wFX
IYcRpcVJLctrsdcGeBaRyaxDO8vfvPuNoxNz/V4kimJK5NI5Ni5xImbM1+6L1gDM
Eowv6j3Sfi/SdVyB67WpPDigP7UxbYzpQjY6vUdfac5lE6XNhcGrKE13XRZL6bLn
xDd1Cpu3IqrglWON6aRQFVf6HcgA1ORUo/XHncejVzUR3u4gmjrA/HXHQ+arja3t
Yy5fp1hpTJfug+tl1r9jR+T1fdtnySeN9gBlYBlAmrBHTYcxwcXulJ5ph4jkbwKf
Mj0cpyadYL9yb5QlgeclBda8an34cEPpiErFqYQroWdob6b/ods/zrRxLzc3y4sr
Ir5zXCW3EeD5DJDFuYjMONHrq/NaWVGHb3conZbZU5WcGDTR5V39FGal4I2GCyz1
MS8pxlHv3+OYtxSvh/enH+OQb/FjMKnjg/NV+SOwoDuauQFdVs0YfiQqqNJ+2r+h
MWWSuo5L8JYBPBSb+lRog2ESWrp9/3S+OiODyFnEHDiWq0wRrawm7Vc1YXxdzOMS
d51+Tc27tcU6rbtN4Dn4HjNl53LVWaPPXbZwMAi6XkZc/O6AJnVbGiPiFLKKUuGB
NTFnk1SyqhgEOdmtYlh1KqQtLrSD6M3H+SeNNS3gWDWB3fPmprng/x7oTKjRC3o2
P+6Xwnpkfre0emckeBaMr6B8GSJv1ce+GrUs84Gu10wjmfz9WdMlCjwK1+N+rdIH
3aahumGHEoBmat0z8usgyCDwmYXn8oVFnwpSb8X470LEujrOeOKrhUtz9worC3qC
TXRj3qr6kC1we+UjvNHbNySw55qQqNUMjF378zPGxwjWZHNllBycgAgRPtPoJ2Pk
TBSSdXFmv/ZMW0/JszJv5Mu8mAZ/EdgCg/KwquTE8ehqPYm5TWd/18sm3EcZXjiQ
RlfyXTfvght3b9MBKF4rZw38LSqYndKZ9se2/8XNhTGekuz8MBdXPN1N0EvgyBdL
OAHVSs3cN0bZ4iuhO7iRsUZr34Si985o2OUaM4sp2TAPf7pibjR5akxGIIQ9I0NR
J0QPMhG1lwNT+v/PEZRH4y0ZciesEgWjPm1ZOvGxVAqu/9Dmg1zjxo3rccJGXW2H
NdYmB1T6B2N1e3URiC1OvpCFhCO8wizJAqmISkVjICweBW9oIvlEM2lU5POu5Kmg
eSrQeN22KxTeAYln30nbRRUT/HUyraxso52ZilFZbdBGSLtlz+U2zD3lg8XAGSUx
fPVPVdjNPgzmKaxXSHY1SVlK7Z6U7KRLjywCETxvCnBRd8tSKyGWQVXmOL7zQb9R
5SK1OwtTCx6HxGhalF1eaxIjrQK27crTiWK7Wojs+9EYlHssNHp4LggnYHvAJiPd
23gZXWufDX2UkJgPUkRnuSuMmkHlIIqtRlKcj/UO24UuG0n/wIwxEx0p/pHeqDbS
ANXBhFomRojo1RCQIYbCp7t/oRXglQjb9vYtFZqqd9cmJHHu/c84x9FO9n8w1W42
ITo16bOwqfk2hZyl00wp6wSHJkWdPr+BQ+ImQCvjTkL3+BSY2Q39XIzuRuxawnn8
2w9OsVkLaXQIcBkelmHQ3N+8zyjRudjemvoypEAMn1VzXJyTwDDR6M8jxtWUuDj9
dMjOk8VVQRcUC13N70VjPdW0/JLzKXAlcHmDBt8UH1f76SFo8OKl8xZazFaTJZpz
MqEzQp0XUvTtpSvZmEpEpAc7IMijkfVQ959mnFRLxGWA6c7m79uQ+WrnCZb3TtFe
11+VbmSVINMPzpYbrY0T60HebviHGQbAibzptke+EO7qndmnJI/JLu6MKngjbeRk
9gTliDERmCvG5FGy1R+CRjieKf6UJ3/RoGK49fvs/m8JzLXRynGmWHHFfc3wwt9G
um4CN9nxyKjjeVdXUFUP6K+gWqwmeosYmld4MpAm7ND+LC1mkA6dNzkgDf5gBjc8
zeIX7IW6I4rXb/voQESNIxTIOuUprSqha49cHQT73I8hOrw7PyHA9TeSnlqKYMf/
/ivEHnqU4BMyOjo0n9bB5be0JZ2UAx/ytifHGqD21MKsNuMCYxCFXNF0O2gGRTjN
lrPv3yKU37R+qwquVxYa6wDTleFyWe0vt+Dw9WA+/0ltRRS76LjWdDe2Lo8lHViG
hCwOcF6nw/J/aDFeojbHFdjLiDRiDPD+AUAFH+W9Vk0Y3C5IB3Nc9g3LrCe8gRYy
bPDqToWXhnP2D++8uOFC72Z14mPm3xh7b/bDZNL8wr3DyPrGszR5xf8iBE/SUoe6
s4gG503qYXBbl9lT/rQjRB9i6r+8LIM0vIAwWJmMeqCpSTWMAEqC8ZrV8HLBQ+2p
0Xo703uowmo3ci3OTUsd1JzfJLuG5nKVHLgw0FYNgzElHKXC1zKZnm6IY+RI21SU
BFWVfChbbmjBC7W9VVL/N4Mw0Xh5YoTpJjTMueZaAH4ArJCjTtCeHjvDvioUCy+G
Yqs9cENAwx7Nqey9dKErbLhgQa+OszlwYMVWjUXrT0KpmRsUEMaZXHHDySbGu75w
mSCdTeeRnKQfOAZx2vtylzFc9CmaNyzurHXFel30COsAv7kKFQ0GLRFR1wxlgyUL
Rh142M+rUBG4n9QpmsspcZsY8mle3v0HPQNIg1ntcIheRMhafj1b5Qr1F1StkmM7
Q5hWx0R/CMRY6rYciGmVkjX2aas8/IA9E+gXGtCDEiJ5ca1ZWxfFUX49iHw95C4y
/JFVQUHdnlI40cI0O2Kv5D9XHC7MzXt85DR8171H4Hae/URBTWFfE88Ul+olSrtW
+8a4nhOorIA58LedSfvSa3XYGuORdkPh29tfSAg7bawf325Lei84r9JRjrwVCItV
br4LQ/k8n1NRah3RAOsRcNDH87S+zcyWX14EUjQ9KU7ks+qxhr4HRkoW8o+d9qj6
cTWD2e8sT/IZWHrr1D8NVXTr0kTRG9s+0z2ZKJN0l5x/eRZ7MM56/e8SYgnXR3Tx
yAwRhTFRdoZDc7pEwnkSN3LFvhNaVg6jJ+wuf2KdE+sG/KOPzxARgO0gSW30M7lB
dIl14lTw5kLhnJgU8TPhR8k6EDXpkbNjDt5WMpuqoddBJY6xf0/gebH8EDoThxN9
U995FEovBoP+r0stMfs/Lk2H+QB9O3L1qAYY3C65IapGqDa2p5LW9zrhIiBPu+d/
Mk1DRP8OWWCO8qViCN8sZvDa5oa1dxnLwinpFR/o6lZAn5zqXbuvg9HmvywRsTqQ
Onp8Z9g1IM0MlGa7LgGndWWbou2KAPEfQDwNMPj780M/Kb5pdxSxn5UTnu6YutAt
eCy95zAgDqB/L6dL1ewTr84dS3FWWk+NS/vdGuEUMWALDtLjsgmeAD3fBoOY2Ghp
smKijYu1ZyNmSNd+uBy7r7TUvJehSsOqEqyguOT9aYPoV0WaF1V3q4NcKD5XZN9p
irTPrpZSbyFubasIFOJZP4E89Hdpj85VajmoRgsEX1elU3xwAD873honSa5gA5fY
nwMHjI+6AMZcfZbRkgrbkqpWqFbc6CORdLfpOoI8P/TkDSvCjmHodGIUwwv4qYP/
ESrPXxH+/uCECh1u0fP8oL/1QtK2xv366bD7o+c+9yuGI8/tA2v0+DKxTMd+B9kb
KPwKBHekwS0rXoIYcmrgzsZ23EfLFJ5q0K25Z280kKWPAh7QnVF66w7MqjCndw8D
JVqkV5+sUqNOpXB3yuppd2ygU1RTugQKRNB4C2L+Pd25PXhh4965niX1FaJ74m+N
bSKD+gRPjQEW4i1Yx1X0yp+N246wLXtGFMX52s0StI6SVp96uV9XAJJE7oGLuyy/
4PuwJyomRZlK4CrkqdXRtLQUzlNqc2foEJC1kvwKcSe7Ibt/9qliMkk2hBDcdMMu
M5Z//tZyoGEBXnKXQcRlZNOXRWAtEimxdGcMrXcSo2i9dq8fMsizxfcKF6HckCpM
i3Tp5UuoGTqIZW8YdzkjcZN0kJqWkS+Cedma2avK4iRQk5ZUvGCmJynsieIb3EiO
Fp1bsNLDRasygyVy5BGNU2+FPernc+IeZUnW8dpfuB6fIhI/9Ly9+a0jK+HxFLAk
YTSTc1Ep8k8v5U0qqGWes5vCUzG3NBb81V7rhQwe9168PPdSCDj2QNESpBoFIwOo
s/nNq8UeYD2gQGojTP96yDGmhLxOh2EiQAYk8ucvOF8mptXERsGUSzgoKtEOXdq/
zL1hapOgdapKeV3RQsRdbJT5OWmN3vL8ynu0l4hCJG0sYoFvIcKmii+woITOVFzt
xwBJ/C5iaUaGhevfQx3qWUbaofVoY5Y+S6kV2c5+QfCqeNUy1PE6IDLbC5MBY8qm
DDZ9Afn81D14Ekh2adBWdtcrlulzCgPMumhDYNRLbvdvINB29qblgKaHq+5TeDiC
RoctYrbB1bJqaMMt/lh/kONQrxgAGt+jPBaXDlsR1DnQ6rBq5G4NKgampI2oC03n
KFNg7ZqzCiiYHmXRDi/el7ZiojtThC/Tvr1QVFgYKkzbkBudJCyT2zwshL4XWqVI
eADp2OSYe4/4BTNHQAX8f0qmo4kk76voxibtzy+2ljj0+fWNpo2marAykiveQsDU
ylyb1Qe1MrJD3lir95Micpuo2AYEvriWo8Uj0p+hgySorkNFk8B4t6qS5ZyG6J6k
XBqjzJjTOP+n2DY6fh871nZA2ihoLZNPFv6/8ClV/bUwIkPYLoF69/gnJGZuaUGf
MN3BBNTOUzMcbAy0hRah9LaXtbZrAdwXQQgiBLeWnC1egfPZcgOY26uzr/ug3bHZ
rPI80SZYA1t8IUABo46pGw3iX0tLyyKjsVxUlnhbVCPvsZeorzEIrsJn3Z82nQut
1xcGFP8uCzU6yYyLcZC9z69/Mxa1dKw+zVt7xzSTO/0+TGmzWN01OVXlH0s1uXhv
WOoRAGTbffxOM5YOAhjY7rEWPglN37bvjibcEfHAUtpoLMTVDbQXIIT427oJVIEL
GxcPZTDQDOeE5u+VZ5yNa4CMbCmrHBjGvXwpR79JmwcKLllTdy3O2jYxD4BXiTi1
q+ypFk0+Fe89+tsCOtmeuAPrPAgwT2VUkVKPKJr6ac26sv1v/CKsRv4ZF4mKaVsU
dD7Xipxt3tI3xm1bSyddFD00cZ+5FoMwcpAIvRun2gWaQCqWBYGRlJ7t943WobbL
Zt7hHDlqnEt7i482nCJKtUs0CQHTOkDRbkg6WR5LWifZpV9iM+dDmBFWhmSty6EQ
rG8Fq/xHNFMbx4hLJvvUPqkRfGg0n8ufYen5n6318qYniz26BgNjQeDyIipo+IPg
wkhFUgglNmNqqr4cdgsaDEeppr6GBbur0t5zWjdXTr29tXsUGWMzskIf6JqCbRu/
HHjCUzHZ+b33V5LDwzJFPs9PT4MuI13QZCPiMMpoUASssBaTso7IAOTG8TCP4fKA
Yp6CDDVyyQa9YXe/6YJHVCEWTkgVpXpzzj9PQHvmpImnSIFDyzlqImEOOzWXA9XH
clVwpqfWrcWDnxTqBLQLIYzO6w+A+r9pWqrt3bYsz4KjBoO+TMCpv4Ks4G9JVMho
f+sLnC4iG/yWRe6ZiuKEIrFQxWA9hI8P9AdySRIyyVMVQG4p29r5lZ86wsw3JJbU
scGcz4AQRaFDgAVnDDa8iJ2aBDxQv0U+8us9eUpY7jcSRk0MRtzwPgCT2+XLg+pc
Pqh+ITDu+2yCh10Oftij07JnNYtXVQLN/3f6Z5efUrWlCawrxSuMSRbaEV+ASHAZ
qD4FpkVLvul1kQoaW29y4SE9243GYbLWhEinLfg9BupaVGfH+74+5deXRPZjnMMR
aJfLFBVsfxx4iI62r6bbbTc+9n+6OFxgwJEZFPghFhG1Blr6y7YNlwh6bWJ4f8Wm
i7q8/K1YKhr83lhcfwuF54V766VpvuU7CDrXnp25GYcICo9a6P3OlKs8izMGNRMD
s+pEqZG49Ng/14PjTM2zj7ZX6rNCq6oVHdwLFRZNk2nRnPIN83WLSPCx7BKdLbd4
1af9YbgXG9WF2Cy8UZgFwtl9o14Jeil7H7MqL8hIbOl1xXd6h2OD2/1Lo9vUydK5
Gj7NImUvumatznWT0t/igY0FfpQNihrHcMotRV9DJLq3rCeMoM5svYxXJFWL32h+
rXt3xXLispMPYyBBElhqaTX8/rNFS2q7U+Qp6DWCYivhIahkX2pNScHQEdUQcL59
UYP/Q1f9Ofm7P5kpUmImYCY4pRSaoXr3eyJU5afHvWGk4gfJCXN1U5o8RZOzeN1w
k3xE4McrpEc1m1LtJQ9w0rP9qt6t5I90Z3pciR55+NO7wr1d4/0iZv1X34N4CQpE
SmUuhl7BP+3UQpY0FH7PMNPXzddsFTTywT2PfKQmrOgWQcRzij//0sXHHpEjVolI
7j68xixGA5+ESj2uW2IeWrUdA5Cd4sj7KsPHwi+onac29P7dxxQdaBW6qRHee2NR
8rTl++TaHTjymb1ULeccoAA+gpSYleys+nAsk/8rGCjfpnpMQ7Hd+Pb13whRSRXj
xiTq+/ZPsjAttk7CNp9PaT6WuNfeMrf4pbILuvhNo5Nr2s6hUHWE3/UFEP3s8IQE
OPZ0Ye71gqDzyWAecqoisQNKEKHxpqfMlK/0mMnO1XHrEiWW889uPot9FID89sLA
JzhxBY+rPBg15Ft8ka8/zouJKbOf1Z3Z3Q1/aO2q2kjTDYI2rS3VfvkmFMOvAI2v
ZNNZwS1AKIsFJan5ZwH8lGuc4RvZ5zmUP9DomSI+FPkXr5/tsKXFNot6Hi4rW04Q
4DxY6HSu6Op1HHzsUUTCM5mSIen8mkcccPq11+jqkZ/+H6QjbT/PMd01sNMVXXQJ
0GgrjzcTSeXMcawGL1GerebIFqErt/RnRoEQZj2XKAN0RLx/XB+0OVjPhFzvz1qr
Ng0/8pY7wCt4OHYygm+3fkVnekRks5LbxmKnntcKFFg/H3yuhKsZjSYY0btdhKa5
N4ByxB1UoKMMdvsQTJFgtC70MWCuSqEVvWwq9YnhSRKY+uMc5I5b0B+xJp/iQ786
fO16XphCl4hmEyRNqTkGHeAgM+Cr/bVg0vP5eIaA0fbtDj2aUxu7YPaWRG/0GFa+
k9ZLwTYt4f57Ho0BfiGwTgJIDnQvrqP1+GOmwKT7wkBAFK9HH/FmL9l16wxt8prE
jGtTGstBitipjYFZ6fuxHUzBOnQpKm/fb7R+B44Gyo76gKRfpqswhDiE/9X4recs
SJTY60hyL/5sozY7IrZSmspU/+6cNP5+9cqD+gwrdddZM9sRkz4zDg1iFcdal0U+
aiD2YKd7GzpqiZF1t+NXri15QXGUvSGEc8XqbnK/inDsVQk+U+TUQSEKkkF8qt8w
mif1AdsPsD3sL5wXIbB9G/R45h4mffoLvK7HndYNE6t8AdMAdyc6Dh0Jw4gbLsRJ
4/Xq8Z+ULYYDNmK03pq0Y5nLsnouuCXsawXX8SxDKp0zwa3Bq1lvZtGnSxDTIWmc
h4+tiUIXyajVuUH0e+/AVbTnPEBkHLEFdkhxkj/UAxUxpeX9hRjicVJKxuHHvdSv
DvtvBXoyK9wMf0ST04+2e4Kbitc3YsMFAQaXnfYmUqmIiaA2tmUCYjUOIVip97j2
KAqUF82Y7Ges2EYo2Irql8vtb0Fz1Lnes3pwCP4AziNdseOXfvqg25czDoJMSbry
cCCmzR3mMymMV0rVFa56vfo8oftMHQff+RqUMLwYxFBTLwBAat5PEgr796HqGeMO
eQEdw2P54wyO6CL0BYDgLlgw77ieuMiFcOUEzywXq9emEDwrdtVHp7awUvfzVM1k
uSwlD8JN2Pziy/un/0kKGJdufFVVeizqB3BjmtFZMq74Ieoou5WHMhfpp8QpLinu
ZNWOM6zd4FJUrWvIHIp3Iqta/b65gxDNvuNAL/ivAsAWnhqJo486qkTmJPCENZH2
DkNWKQMvYgK5gXJyIy+bJMq0e7t4m0lAlnV5RxWCmG6fVWcYtnxj2JJlO8yYTmPn
s7gq8eBnT3HC0L/poTGe55nMkM9w8KOBMaCju6U6zGOafaXyXNC106E5uxvvhoZj
jo4Yvm4C8xtnLxOPzaI38mx+xa/fR3igzWy2lb/StzCx6mwLH65TRUWGcVyFJwD0
3h3OJ9ck9Y0FMwtIbFhTwsT+gn4JZh58nDf2a9MzzrfimZkKFcuw6OclSdtgc0Na
MxMzUPZenoq6r1beV3HhKDIMMjMolKiKVrYcNlUDuo5fFnhZkV+UEMMGA0a4EAfA
ZR07DD2UCWZMc/p7wA5NbVy8VJtz/g48WK/l4GZ+tIGuYgicn87H5F0dyXj0Wnc2
Eg/eQ1VHV16/yHxHYIO0ERvYK9fRC/Hsf1megLGPsqmn3ztvvbQExuAB/RTCEXO+
1yl4cy/DCOfPV6FS+2QuB/jv2jNePJE0QsuycWZF/B5iG1zlGQ5mm66KNeApP9Wh
zkLu42Z1tTqC56CVZl76Ya7FPDdAkeyCp6o4by6VQ800Ip8CqoL6MmcVHhbMCpkK
7Q0XDG4wW0UI1UDuNAJhnBcxdNu8l4DOTlSI4piQAZq2dMSjzenDmP24zV/wGWO4
3GNVcRdxqSM8pkDLxe3e6PwOIMTz1l1QEz3C/N9iNvn3PIPvJyl+4rfWusahakEE
oZeJ6FVbK3pxy2qGisIl8oNsn1NHqeSgQJZCoMD4vuudO4k8ZwhvuOe7rAzn3JIH
v3nCBDZdSfQwRDQrK2r5UxFuEYStKLIk4tO2cHyMh7750UahMQB7nDuwP0YP26SN
IKVidzZXviSSOIaMjmjyGY1viVzvD96FkpO98KHUB4IM+dfiwI/ZrqfnuQZmzA9K
HlpgS0jBxDVG862l/ap+AcARmbELhVf9kJeAA7GX55zgE1hhXLB7t7cSLSzqZZ5+
rLBM/9vkntqZ5BZR6LNNKIoZMrLpg7OphNZEmwhYozU4qCi95Avg1XUw6zWZT72I
qQHdqSXfiW99GjDY+rH9oZ+9uLvUWjDV+7ss5Tu21YcCJ5OfV7fCjhIA5+hL0FkT
JN+22tqvRexQC1wF+WrH0eJTVf9ZaUpBoO0d/swZh26EZ72EbLMMYT+eiyfbmDWm
/0bqMm+AG+pSbxFexWXQDWt80czjO+7NdDnRTZH1tcdFZCfDdsRPyZgrGCGw/l1q
9c8rCzE02so4zBcmvXZ6c/urebCIc7dji0nArh/WCCa1dZTGUq+xqyblP0Vmyk0n
Uda9Mxxhx8VwA0A04lNXFxyRX8gBf4xrZb2CEwBlWvPu9RDhSFfbXsDZMYtmAapw
5xqMXyhlG3hvnPc3PK9tNMgNXNpvpmDehB8dd11pYESv51mMcnLm4hwOejgerLFF
PjIi6/Ke15q1elVI9LjXFrevfop7ic4MqQZDPK4/Rt3gASQB0CJ7WRkCWYVwcNSU
Ym1mwvCD5kmEQsmww7Vf8Ezjlb9tMrUuPuvVD0K1hfGi22gGL9b3bImKacLuj582
aLd0cUnd7Rht6lhQalNXL4D4tL2UTwMI7jl94kxIlv90+0fyC4W67dxxtRS7RXW8
2MmPBieptZW62p1QAFkMFCCySa0rBi+1Vh4v4GLXD+u7aqwdQFarllmVktnyLwNl
dAzP9lKiktVD0FWP59HFpmMNttZhmlRYP6NfWvfyRI+puRPnty1QtMcMoxfS8/e9
IkX5UsFQxnTx14KkH243vXWFmbRiJgpFRTbkXkHFkD957n0he7GzgQCv1auAYnQ9
EXRfsFa3uquLgG1cVtcM2gGK1/gxYe9ReD7I10zOeptp1kY/m0nt0/WflMVxhgrN
mI5vCUqXCMxw6VkMiACam+p0HjaZRlyXWlZ8SsAj1At+R5shPRpIg8BBFbGo/5Jk
hrpJdFNL0PBSOmo+IROugF+uOdmXcsarXYxB6KgtU1nW1ne67S7fqGDtoIMspTgT
i/n+8z9++DKz7N+BTJIQOUMhsBFHvCkOg6z4EXuHKPzuI1gBeVhvqAovKVjTd0vJ
FzMplsM9RRYuiUs1fZzCzXAUDZk8uEO9Nkg90zeKqf7ICsZoyR/FHX8+RLyelxoC
lrEXHtJPUvxRgDZVxxTFACgzWdo7p6+GJGxznP69KkpSFiI/Qj+k5WBrXuvjgBCP
1NTtLc3ijiTB/Pgy9cOALbtDy++EIf0dZ97IuZmEIFkBmbvf4v60sbuPiH9F0hPx
mwVPWaNcfEUl9Bjp4VUkL2AGnwokVZ4wJ7Y7YUI0rzHbhoUIxJE1aRzBi9F5AFC8
FSfxoRy2hROzEWr+pFQevG4nS2rbwTnS76dNsXxmZC5+Q2zFmaUYcOq07AIwY2fa
AEjRt40QEYb4wfxskQ21vZ0j2clByXp+lOxWcFIXItJRv9DHiPCUUCmOA05wOmMc
zeAwi6KPwVhaAwJ5I25SLQ1hKDJc3p03a7KP+AsRhr89BNiE3OTj6pOCZmZad7HJ
fP+JzeKP/Ai7ezwRqFNHjG0YmSdlaa4zXF7VSvAU7ekTDIJBL3Rwp8n4DJeP6V+W
cfld8pwmEDLnpeiXI7jMweyKW3V2XenFi/aprAFE6Hahsd9j1thKoSwQxBdz1iWJ
+qdXDaR8NslrMttRCXkaMvnp504V89R9K4K7/ytrWJqp7J3Uj9bCUNqfYDc4wGyH
ctblCngnc7JNMGywHcu+removgaTIfLXyLVH/EKx6wVoUyZ5zkGFPTlc++Vegf4g
mG+pIKzJY5RvoL+RBMK7vAKd8U1ARM7l0jc1wBal4s3S4wurYEPafPwgsmqCyzT/
xakw5ar8L2R5i65qGol85gSr87dM0z+0hBAtz6G6y0wCTPB8EMhXBjyjhCiaGp5q
Tli6C4/DWsDEtP2DY02h0YQ0enbGvfq8Xhxk2EAhBYv2eDjdGTPPMYW7VgdyiTHi
tOjMqd4Pd2YH7UJkmotS0Q9s6oRXoVQ7iQqP7m0bHp+ZGDgSY6LrWI/ghj7tGC6J
Ib0EcncTN9Z3nzwqCprfu/frHZqo/MRpfDyk6oYTXiM0P/s0EBylrgLgxW3KHgV4
PUgcMZ2MS+E+4nRgPo72A3xwZjddNy/hXgJOA91i4ylIsVkca74ZU0Nwq1K9exP2
v8ae1+kAlNAngfP3C1Dz25eo1181TbL1M7BY9iByArYWSHWEOBP1YHj+LUmZmHGZ
ljvWAr2GEGWT+EKCyHV7W49zSD9/tYMefQn3lc0dD2fkuChxTbS1bie/cK4bAdBq
I7REWIPDUV07S21teKsKUCsAEHyR4BCwuE20S7l9XHWUfOkL47/gtLX/n7r+azEQ
rQy8xUeG5ngntAMpMZSw5q5T5gqYyqjFdsiKMwDOgy8HUG410dqUelFQhAm8p2HP
uTw9MmwVO5iny+octtuX8VvexPkw0Xztl32YupXmQ2gb6/IQltREI5IJoSLVy6Xi
IK7KsfkbKMgO4l7EGMsp7DLP8hEr3Y78fZRNhmdXcsSeANZRxelghDzMfEU/CCk7
I4dNWbK6n/5iNY+uMaID2ohjlY1Npuqy3h9l+RTIxDueKA9x/ogt9Qi45h75Xzy3
numyVPHZKdlIe2+G9iQw3xY4um8PaIARbvrvAxmxtudiqjeq23s48eiXzzd7gaEY
RVARb9OsjyYxswiUXxrrPPMJeniWZY5WnRrO/5eBVtCDdhHgiLLhyDCGl8l4Dk9R
3wYXEE83vEv1n7ya3GEPunECBgJiSekBd2eQ4QnjLIxW6XPG+KcFW/bT9d18Cmvu
LUXwTbAvNYV5xo/dksEGXxRZMeZdOR/S44Z/c6LgcXyaJ1ogndXxvl+gC7j8rCtK
rcKclPErbFy3W05LpkNObEGaD+5jo6+DsYE6H9Y8oL8Q3PTs9DamDv25RPYZgcvw
URsBFXktzQ7VK9kQ4SaKKcnH/VKjlaPQSC6YlXePH6ZCzVgg4PYSC23M1x51FSt3
biBxdJ47jty9WEdW4kx2vZIU7WJCIaKzpjAAOeD8VWhYD6PJYdYtH/J/HifxOu9R
9xle9DzRkctm/EBq377l+uSIcearrmQgjhFLZYua4TtIy/MsKSJ9qk9kWzLAIZUd
gZg5i0oVhNnxkYY0DSbdZN1WYg1TsNVOIeA/WU/Fc2+QdKzzPhF1g/cq8Iiw8Bsg
4WPgV8S+Qy2cA1s/zRkz6V1mmxoAYeZRPxE5jsaWMBe5BeLKHThbt/AQa2dGHjAl
sOxvLSPQn5qgYOg21uPavBt2LPtv3G1H8jt33bNWP4ek5hZLM6XJX2HwYHCGHs0M
VOaUsVAk1MYsZsI1Uf7vd8xjPm2vjPcP0bIzsMfKYbIVn0h5U2aZ0HELVN0k+EhT
asUOHx/eJIGDLuBplXqj1+NE+yzt8DArORLPXt8vvKc8wxd4yN6UKOqQvPK9/Am+
0JVVFnu/LfKZ0GriTJK7lbM6U/vGloCmCJ5aT2LnnYahB4l0I4ZeiGQwPHb6jPOH
dGIfwM35WA6H0FMMM3bC540DeoeUBRHJNxc9xLjJk2gRxiPptK1IXC5Pc1FLZunQ
7WH0tmlniMZe0nWgS+rvWDGMN5HODcd+aa1eaqjsHTQW2Hswy96O6Aagljso9I25
DEyBFvu/Hl09qO2DTse7pKCAVTbiAQi5zOCeqRRDiFYdhlJhp/Q9Ail5SM9Vadj7
WqglSzF0LfCBMdM2DCySXLK2OgAv0h3/Mbme+tTUGkHMvOd1zK5euA6up5EIkFC3
v/ApQoJcthKgN4I/3+vYukGLsIji8TMxylvRfmCypYmbcr1kMhLPEfJwkES+weFe
oQZFyNObJHQ7Zme97Fg9vHAVhrxFbSP7pO3wGRp8bw1abQyn/3Q+b/hYWmerH8LR
op6Sjp7Qkmkmd1Dx3VR7nVW1/5SWoDl7CKoaJXUtRY/NZBkxISw/5fNOvTQyqIRf
QCy0ieyQTmNZ6Lj14dynMY8I8/lNi/zxqVk66Fk1EGkujrvEKgw9oDUqDMVZbDej
y1gKonsDZqNAeWVkuF2+6BfufGIJ0j/d1fBupoqwOemkNMlQb34oMGn+0iVkWFCF
yPgxo1W/iCUCZpIvWf9lBqv34ycMoYJ+TWSaGJA9dKxr/xazEV+xKtORr454DdPx
GII7MQin6zITsZfr1ww2U28NZQYzZKHUNe63eev3aIhbCMR844g6By4ukhud89q+
phmurCsvz0Yu0bLvvCQpeCcVHQ9j9JtlzuOtsuJNJY1g5Rcg0Z6FSZ5f5Y7GKrFN
8fbvw/PVwIW7ydusOuOU2dYlb4IjJVAHOt2/CJDFD43DoSRdCyrc0o5gfA+TzU61
Vut0WzBe4zUgSBJEqRRBx+9ke+Xs6PxsXA27rwwF8fylgHZlVnZDXj6kzoyBwO2C
dBZXtT2ssDlkwysapqLUbJfYRHgEZpmpSmka/nEoWG/Vuw9rqByQLR5cWVpgE2eL
bCOUsPBtSHEzDtvz0rXHKlsgOGy2zntQAH89ly3w4d/Fbs0H8cbldUdXoLzB7SYE
PI47n+yE/DYF/rJnbq/2OdNV+afRZ4PDRVpB45jH++sbnPP6zr+VMDVDMHt2jgBL
e55gUeKmyz/gbOSdOpcoL83sT2FYBfGytIapBg97ovfCFG8AEgvYy/r3Q0oIEHHq
WCJKgZsRFovhP4Uuok7HKcZ/Z/FCotvwxDLpviKE8JWgM+rE/tfXt8qS8BMEROug
C4E4JMBWjnW0woxVFxoileK+RRx9NoDScyNXK3VQ6jkCM0wWxJfUNTwcL48nBIMs
zUdwSCToWHawvJwYkaM+ZcBcpHbToa2KBX1/XSf83yl2iwYAPCiBQ/XDdKWqexjf
7+tVkQ+7QyfdaM0rKqqG80jEofVvGKw8r8vqc3HHNXS7KjVL1pg1pZJ1S9C4PvN3
OBU87lyM1aS3x+wXGOiWnUN+XMHcXQ/bGqOprZwZYdmfscYwuiJ2nQaMy2BfeyOC
VJCjnsN2LJF2nxZ4L1d5Vi37LWMCq3T7v2RWyOEXIbYelOshUJqAOsNlLizt1BYV
oSfLRVRIZPD3Cm+U2eTY1c2tQKXoNi35x9M0J2SxXMHOll5Ss0yMChn9VPUVPs/K
1y/hMz0QKad2EniFPB1dbDe11to134Zg5i1fAHOh2YrxyjTFQNE1Ler4B5Vu4THn
Hj1VKjF0Sy52LO7AB+VwRKcQ/JQ2IuK1ZhAeKgWiIA9abUiproOjUzS5Hdccllsh
khfvmiVx9nI50UgXYssDY0yGRciFpcAu7Uxhq60d99wxuZY0MoBvc60gX3WMf0x4
I//5Zb9cfYP/uAD8wJv52+7qGrFEQkrKtQcHkEKTHaL9hBZVEVAD88jyvQkDUO0U
XKAObIZO6G7t8Ak7pWJKGw3gCO3n+rtsIApIb+gpPQm63sKvZpWDD2sYq6FAWFjz
nCMrAPXGpgOAyoLPikEo8uxNKhSz0RQqNmFmMIiJ4uZMyP3+BcBOhO7nEGVyhlQp
NRAonNgScJWKchmsY3/9XQQTjKLSxhDZllD2Ykr7fdNLX5cWRyjxdEz0GYmVtEOh
0hSKW9ZsmT/vZtwJJz3imsAtFdwoYjYIV9biwbdc4ZTuUQVqrWqiBN6IahsVVwG0
rFNBzmcs29CosX4xAQwCKFd8al5wpBzzDqIOO6sWG+tvtz74fyzofBw7rgg0AHwV
yhQog3iqUBq94hzEsTfIW5B4MRcJS41POkHSDfcZapIX/FlWFh/szFMAp05n62Wf
qsY2JQXAY0Pafy2TEW/Hn93o/BORu6OiNVjPT8G4/BcqQLn2OnUCwS4ZvqBS5nu8
f+pJSGi1fRe1YcTcquUpFfILI1kpLJEpJB/9b1+j11Nl59vI1x38jo3jssxM0NVz
arq83rNSe4rAMqsAZ1ZzRFPrfUwpcrzJaJ+VJ/jE2bUS9ByMvNUawMW6EbItoK/l
WzZYiReRpCt2o2/vWVCInEMfIR1j0QZKdGQb+1KJM6OpVl7tPPNoS1wlIHyl+HGl
sZa3fDW71Eif/BNduSzTY6CgfcHXHw0b0v1qol/UF/pVrIHJ4c3yzKuiM2UDqYKJ
8Cnnv7agQoQPhncD6+N0fHg6j86JMLoaxgl6jZNyStNRAEcVWAMf6ZL+Gv83YlGT
Q6Pphu2To2y6+5INyVxc4G13BGh1lhxk/6Rf2ZXIY1ICDdjtBi+Z6KVJb0Ik5/m6
EDSaCZWdTdZU6AuoGffKMVq95PAZmu5sVQzGHHDG1iRfnFciJbEbG8RQLCS8X+CZ
J1iTLQ0ix4Lu2lisdDp+OFL9/8NIyefw4o0/Lu43zp0Z+VIwhr86qU04AqgR8qIW
SeCdgZw4fX3YuynMLI8L1qPV7EBHX6ZYvhVTE0Cqn/3uTomXP0hua0LOxpNjmlYu
WNuIWo3nymV1wSzVNpIO98ADx31keAxL0mhWwVAfMhKdBIFLGvQzVhJ8A5YtZEx9
MQlU0L0OechlIntl4fItBRDc98xCPltrfGVgXWVg+8xAx8EbDLRKGPq/wIEM7ldU
rKayMuk0ogKv8LRzaHgCe7ANN08s3nXcrGhE3WZdIX/K1YNSe9c03r0y71kg5EUi
joTW/SEsFVKrxnsRPIi2V7TRGjTCCUbTMD5Cv9Igx4Kv3XY+sYwganYm/yyoblPg
Duk0QcAuMiS/WNwGLYHXV7mN9/QdOOlZ+1a705sMIWV21oxss0xF8a0zhhGRlcYJ
2BvS9rc3eWvL868f6fCo618GCHR00zEz0ytCB/8MfUAPdm1TKg9gNmqZFt04FjNo
0hv1jOUycfp7+eeoruTCbzYXNPIjmep5rmKG6mPTZz8OuSrHckTZNp+DHd1EX77s
W1eOTPmkFxWuQGoYYvK/OCd7dPz3yUVYQV+HSn81Ss25DfVUOWWYpASKV3aqxsnJ
LoJ/1ZLGnpSHKApXR8TQ8dcQTnPC+acoobNx6NqKIcTHoFulE7NlkGSka5v6fzSX
D4NmI8RTbVdPKXKAxu2aN1+cpK3hszdHR5pxWLsQZJb5K6CAHdHnAbR4rHhlGIjI
ZpL1bk9I6V0HnBTNwdl2JdLlBlTNDAjNTJt5dUwiV74yVDFD/fNKy4j41TAtsURy
5GowwDepFFguKvlfCsBHC16N3eChy1G7nnwst8+zmPBKOUBDErBdozRsJnT21AsW
9GrvmUKwHqMgpSRkFrp2bt4oN4slAw5u/ebZkZ9/43PvVdYysHKCR3u7ZkOXXNeh
ipHRU3iB/eICKjR2tnYdAq/DNziDMSWYUD7IQUjjFw1SOyQxfkJmoQjUzM+hQ1R9
8xSwk77SwGSR3a3GO0drw2pzso9MMqDbVBgxgFGjomh+zvlw4kEAK6jB9H1oFHAT
DNQiqDyWK9X7odrXXmOriNSdpcS5BlSQlbdjsoZfw9rw0Xgr9kNbqS2N5Np3BlQY
JAhKN64mB3d4XP56KVvbs5tNUQXrNqkI1g6m2fQcOa6dNxmP5ccfSv7UpAmbctxa
cUALrhAo1Nl+uo51O+cg4nsZ6jnpm5jEOaJt9AHjOLZX6K30OddBLxI2/sppRTUc
9SiDDYOmO0Tjef0JUCDR/sGMQEJvzaZ9c4yS4uZluhpelmuoxqnwqrpsZ+nB6sEq
KVpbvHMEiNJSQsfkW1M1PAKSHSryRFiQePXG4Mc3aCdpWN/Q3NRO1VKckwMDIbPN
ExRtFzPp3Ue3jPWBnU3E4+s0gqLbzKzL0MX8P33iOV2//3CFwt1iNHlQ2R/TqyHp
gp1ZcT/MruA1CEcO85w2yJFKHVB0letDyXAkBh4Ges5kG6ELCZfXTynpAW4VQPSB
NLUv/7sjgidTu5ryGUmK2qsi/80jcWHicoGIa3Y1jtEwl1R7qQwvJ49wvsoV5Mie
Q/ia6Mvw8AQZ6TtnLwiEdJKplOFYgjXRA+A0lfRnUls8SXby7miyGVtnbtvjYzFK
DeTF1BF0/0kvDKflvD0PO5C75ySM0gs/ZjCugYOCBa5oV5gVGzIj41jFKuAvtY01
PQOd8Dh+ajXQGrYNJ2rUIubm8oxbcW40fdHk7u561f8qdjeMHgLtLxci3MpoXMn9
oLKZvZjyxjjSmtZT8nId3fBqgcYtvkc0uVgejb3yJAEdvu/J4sDsL9ulUDN7M0/x
UL9DQZE+ki6nx6QPVWzjU9erC9xQEq5WchQQmJ5/ZbnAY83U2vYX42N0vxnLLxSI
lCTxpHFeB6g7bYyttJJS04dsMfdtPK4EeTWIlqzm1fe62TK0NYuy5xQMEVImFvFZ
hST6r4RmNrUcXqw2QA3qFAe2F69Hg2wOcXh3XkRk3hT7XY6XzN7+Thi/uAwmvkF/
szZv3ig6rk1uI77b8vMad1nW8V1eRDqHzKIM3a8u90e4bC1DY6x0jKlpi6k0rhKX
boNIjmC7+zgV0JmELJOGc7as6PL5SRZfP35WHhq9Oe9kPqW/apbz+U5yOPnDI/Un
esOKHTzLq3680dLnv1YjG9GMPYZvdKbCHh4ZVRrw6w0uQ3Rp2mY6QvobF0RKUvPf
UE0x3c751eaD711RaJHjry2my3LDdUSUCUelEmwhOvgzJPJ3Z5cg1paV8ZCEA6sx
Ryn47drni5878TgjaIld0T3k9SlmYyTC7C/VoIl++MTf/GVc/Bvw5Wh50KAueCL4
yV1T44ali7RM4iEm/hIxgWbvOX1s3ZTFo2sfg8/f/tDZan9NT1WMAqYydQG8QQMe
f14K8Bs0gIx/lfNpQm2RKAVx83wlF3LJpdyn8RWChqehOiFzQbjvRfOwNYE2kA1V
NMIIKdEmR5XI+rqv1qzyJYuSn8mdgwcqO12Oodth/F+oklYXfdqFnBdKUWmGYbg7
1KnGQYYGqd8ed27YPgRom0i2aDRnSewBrB5sH0KqS9Sp6e3lYqRZA2+xemNBB6Hz
C5qd5GjSk6wDkdh6HwX3gilQluyd8nOM0NzdWMhiK83DL/1hFkezF21TxW+UQLDh
85LVCmUK9bEZiXsBkgkMOM+FIgPUo6xaeU5Qqz/yEnyqHf7SMDFhY2vEliiRNkLu
GdyopQ+lrcjqkIeKza9L/n+isBdlsgc8TIHPH41gNy8oCgSuX3TfjXYAYtBEXTXj
LFokARj8VMgJ8h9gEa/Ag49uq7kmIAQ8BQKE6P5422kEPuHTf6mOkpHmfdOA5Hrn
xdkYMuGwGdtLE7QzPdPBn2u+Uhy1S29WEKqTidfMC1VAWFkHNghQyw52e9TwTvB/
DQZOAi74EPUNNfLORBtMqEv0YsIKlyMAZO/6KCbEt4sCOyVEel2eI6PXHEwhuZj4
piBWWWlEW7BgAmp1RHh/KjxuZgWBCNXykJ2vhxLR0UjGnDQ7ItVNpvU09w0fclnF
XcsTwDcKOwi8nlSilquC67p1G6TsDl0V6IisjQRfniy18XkdPBMB5zaSh0aquQ45
ZwQaDv7S/pXehjLV8o4D8/YC3H/okhDIs80uHR/iX/HKm9B/RperADxhd6eeMzT0
kc7+EU0SVElTJd1btm39d8QJ4IE+5W/4zT1HK5xT4LksF0Z136AfB0iGVHvVXXEE
JWOLIDyeU9kczEkXpGTk+9Tztzaji88G08jkwQtpJdjjYEJPsFkGgUlecMlb/b/1
aUVOWUeV0gnl6ZB3oqm8EVdrjQ5eSacC2OTryyjNDdc049GA+8FGyEjPiyOgVIhJ
+Vg2UaEu0vtND7e+lpWvP8X7lhHWokuFochIYuVo5so0g/jfQZ7iVpcAUi/tgBPc
GvSHXUQ0FGyw9bODlm9Gn2qpJGHHIB1vmxITBHX+UPdzlnpQZAVvDcMdLopfr5gl
LIGKbRUVHeVKg1OuBOJeHe0Krrm6u5cHt1e61mBtGJs0ptMQTicCpoF9LNDef8PM
nxWW+Brcfb2FXEazXzdwtnMI6/G6dRMKcIOmx3raDxpaW3+GW6abN8TvHhIWBVP1
C749HYZMDjffXEiywgFkiqOhIXMFT12lcuTvtMN/AVVJI9t+W5d+Cacevc3GmF3j
xTz2CCsPAq6F+kjS4SIW9O9RvDMCpkSEnItvX/2F9Jinl6FjT8O76Ka8oufBKz1q
+vAUWmDuYAMHB2baioZfN426Fz8SNeuQz8y86Wpp+JkrjO63ybdE9U2k+uAQNd/s
7xZ3WyEmgbumMRvISLP8yy0Rg7w3MDmStARpf2uhJ62OV77AWJkW2qIPV2pGsP1D
Ik3p3/V3a69/nHkWL9lmD/tZ5aJMmH1JyGdGhgHL/airZ8PXlaLLzeLV6VBc1I/V
IigQzpvn5+GLnjMxrDvnDzUGX7Vxmbj6LUg2hYLz9vpUlHDEESiB973Yrbv7tpz9
WyeyHXojzu/luxqyu6G4A0z0jFjm8C2arRW+kvXEEOwgILvFN/J8sIWMr5McbIx3
XX/LoKNuh/9ZKbum0wsmvPys6JoxJbx3EG9/Xy/zXn/HY0KQ8vflrbpltSZZza9S
g2eXrNB0hbFD5a5BP0dXi/6zDuPqHzvek2nmj2f/beW9YC7xRBGvR3+He/InwDkj
QQO8MKLVbAwofXWbI4+gkbqjPs9Op5RKdiagzRW5NGVv3AjUx7t7ho1T2Trn/AOJ
s1r07BiL5gARv2Wlj6RaGsgcIGMqFRasQJcFMq2YvBhA6sXtGPBKWZBdaLwUMRvD
OanILdlY3O5RpSxvcyltR+neqZeDH0ok7AX72TPNb6jgpe70k5NsD3sU7bbJ4EaB
Uz0P+OyRcAzJhzFe7nj5vpwdLnOiX+BWPLrs/KLaoBN9EQzxNfXRycNKBQDR3cnu
5hA2qc8hPb942raQVrPyDXRm6Jj1eCs74nStiCfpxmnNLrikmHVroo++sqvmj2L3
New12CpHF9haHS/R/h1o0PerC8BN7X308aitN7vFTJ/wTUEkeyl9XIyL9QY5nrhq
U6iXXmQlexXvQD8KtqR5wcD63RT1pUbxaB0GJwVb9uKsnNUlez3JegikPxvNVuUW
MNtq/sp2LiYmGsIRx0xT5CkezjCCjYxYiFLu7TtfURBkTXMSeGwhSQaiJ/ityEW9
piJwQiUYjWJ352JB/TN4ftTdw87YDomeGn6gs5war//qnI410hiCT7Cr14xGHp67
fN6XgPmRpawFKzhBNFyUrwCQ7oV6GTNOtDb93CFJxiUt43a5RJJ2AizFHGpZl6cj
tlpXIJRmRmfUy/e2pnezIY6u9T+LrhMLjxHoB9vu2DxA+LpLcMq1ze/6GEnZ5Q3h
m5js+Qz5X5Cm88fslctkrtaOePDV4Oyugxf5UgMR5ZtI3yJkA5o9VnyPQPQN1hBs
J8JjmobcYz8cwJqP6DdvOVg+SD/eLRtr5GwEuzCgzFfsWkLXPJ0c2VBcvyRxg8R4
xBqCSjUHDceyiFMCapGfjdt0oDXErcaoE/iStt9AX8yRWt6dq2SNDwAIpL4/C0bW
e4oraVT8+beNDvQBEzE5ZgB0K63lbXLNhYKuma8n1Ff4wsog9nCO3P8OMI6d162e
cgfebdsZ11ZuPJfeSz2kZSnbsSYeBfmMQnVa5ZkbFnkfKXp6JZF7JTOgilGIL/T4
TnrxVt+RmDliRbDFdezb4F1HO72/o8QyRr6aOuMq2yeKexCkNoNUhPENA2FVHtd4
sVcuvZiTmGjvmrXhnJpGz01mCSBFt607dAyR+rfEW9bDKdqsj6LWdLtvEtSnN12O
8+PuOr73Og2F5znasQEVpxZ+46uMUZZNRwtcWjHxb1vOtDG2UPwDSqN/e8xmgoxZ
bWQt3AdRUGeNk1lhd5y0M47vU53/Mf1LaVcCWM5569vX4kiXFu6DYOG7ryoGy8FD
9Z0Mh3RTvvW1KtZ0vQ/0IvvWRFbhFGOVyhWRZccCUrHH1YE7v5wScc1KhaAl7BgP
TFy8Um/ByN5y+RGNH0HRfFi1V3V9BQDGvd8nE2/didFcm8wY2013JuhoYcVEsNfi
Z3+y96S0okz/qhbcld5VFD2g3OYKEWsfPbpTKEGr0pQJbi+RHVs5diciwfDqVXY6
jbRYPjuonGxo2lMqnyBA1RJy6NRq/VRIvEd5qoi70j+qQgYnTILxHT5gZA5ibj5w
Qc4Ai6WbGXxZh5IWEy3BVJeT0WoHa5M1ODrwwYl0f/6fKHrpm2bgPpBdVvkYKY42
gjIj2jsO5XAtlWRxyNuspk5NWWwuHjT3Un4Wka+8M62n5KRJ9C2lmaJfC/I6Dd3E
4OSqw6mnTc1CLE8PPnsKy8f2s7trxb62YjIWEyPrXoQdHEXpkt6dpBhWmplx/k75
WUmyTdXRfNxZIRcxLMO7msE1Au08iG1GYBCStOF4jejyRU89oa820NF7VOTFBAce
278qX8qSs2gCXNOrgwqEL+q1Me9XWKDCF9fUMZxcOMo8gZ5MTbSHctVR8mhnqVyR
kjMTqy0IN29jL3WXR7k3dAs8q4OO9KQXSu4nGU/iJhglAN+GDh6UeXqjsFf8IMm2
bLlZSCE9zYTC9OGR75RlTb7gKBoRcLPnRSryrDmsvYKnGB4CJhrXcNMpR1FsjIWD
nSNv9TwpARH86v+pW1kEWA8d/VGqr7A2zQYoQdoyNyyqRjAyYO9FI2omCqFP4xYa
S1JkRxKTrnpcqIu+ByzaAa7xeNkPZdtbl8iVxul/l6QBueHzCAsfIMop7qqjjAlm
SPhqLrfU6ZPOdAX6ZSfrlh/mG+Bg+gkWSYkZZMTnGPo8LbMzRudsioUsRhqA/Nec
8rScbQkg/7xqJmJtwrCNvjM8pbDx70Nyu3kq1Wd1lV3d7qaxx7ezMYnGLdamh3If
TiKjSirRPG32ilO+AwVPXTwhufYAktMPQ/Bubzvus6Y1NAoQAPdNKNmeoEhoJCQz
P4+//3XWf+pgRn/ZASU7h6ghj9Hslmrc91UrG2WiuNpui4a0uK2bZIUyqe4pqBBn
WgZR8meJWTbEtxIDUn/7Eb/5IXpaoCyaeO0i7s3OzkLS5x0o4jP03rrpgNu+1oqQ
qPfuEqRpmdKabPoIAstlau5nQbFn6KTYgWjHc+vJBmB8xCaokru3eMH/3Q1wxBRu
hPu1To7B6Qiuq09AiCpGvc+Uist1ntyyc9ftHxOj93DIc3ONwtMEUPJlmSZSQmA/
MyshElGKJaY/bL53bUNL9F1EkJ6076XSZQatPFw6C2Isg/lgX5HQClM0jZ56dtEc
egHID+7okwlIRfTUX5PtHcUQnOOmGI08Hocky4UoRdEiOapvYzj9Jnb2/pMH9SFg
Dw4cgBDjnLdQtK3atpfP9MD3k3I8m+K7a4SKDtoopvavw61EtHkwF0aOvyC0ajsI
k4Tk8UBVPMGht9VrBmRjKFoovEYS3ZjlFFTDEpSuyIGEY/7UzM03J8/5E1a0uqSa
+9wgMToAa+ySgmZXFod8+kf6/XEJYfamyWRz7vC+mepEuaj3eNtJ98dMBdPW8J6V
dZU0MrR5KlTIDIRbnhoJlY9ts8xEWdSDdxXPee8SJ+fYo4ZWvr79nb/piF9+/tY9
MsWZyV0GJzCJ2GEauRlVCRiNVmvye8IM0/7e28rxwegPLXzriRV026WR333KwTXb
bV0HAHtU/eOs/zDMV2kbZTWvbxljp1ZYqCtVHhXzS2eGu3pZQeu84+v1gFj4vOwW
PNW6I8zMt2WcnVaNKSeFVKHbYyNvFs12BP1xLt9fQ9mRvkbBcS9HZ2NLDSXmseJ6
h6xVOcYL/KsfCycPyVY03hMinwV5f6uEih486GLIRn7xpqdNXIqpq6+9ykxkrqNo
kkmzOHqWM8CGu/UvMyN/Ff0RrsHi731igrExr93xxGOSVRZft5kAIS/xNtFonbza
rNhmJADeNIJa5PqVN9IARckVfZRkchDZTQcC6ysm49aNNdVxv1EclcFM3fszpvQz
k+ed4X4pc/+cuTxMW1Nkh16a2woRwksa6cScTyZuw/zrsmdrDiyjQAZ88JAp6Qlo
8EvLdfSdFHOleY4rBBHVZ1jPqC7ifpF9c1AhBEiV6S2sYABfODu0zfrdel+/g3AP
MyzUUkIrDH108KSbJd8vTLXtbGNxCVSMc0dhtahl7CUSmXgJzFw69npTC6/iC+Eq
aOFipgR8WYXp1CjZ4gDXpN5RqAIzEmSgh22CLG8FXP/Jz4k7bLM4ZqH84PYgpY3x
mgOiddUssSrLY8D1FOK32884Xgl0NWfDjEmGO5QDAAKRyhj3ZGJoNAEG68GqK6HN
WA+DhPC114msObMJSSpKz0MyyVuL7tbes9lmgs8d+nhJhi9Us493pRRmjahIzTKw
pv35dyrSenNkzOZ1r0Ve9XP9JvTnXa81ztt7+f+yo13scugg/7/QonDVolIE1kls
D1RWbJ4FKVKiwFx06tE6O/WMbgGf2HrYo7uaZYAtQiUrfgMeeIHYl9otNfU6YzsJ
eFRb/HdaUFzZjhb1l3Sq+qC8KkHOrK7coC8oNtiKgLmd8bdbVYRDmBbPJ7n0/nns
nle6zs6zkSrW1IUKksVLr4CaCpN16gNxvdEOS1ZfcYHzL/C7lLzkA+0Rq0trmESD
hA4Bu0shdOADotfHRsEIU/1Nn3KucpAXleqoV37cjrooLK8CjuOjKeZQJBdXwSA3
4NHbxH+90xRjhr95pxCNJ0sxmdiucplITghVWkFsZBA7Ov3mavLKXBfbv4jlElHZ
WVxeEFzK6S58wuUl0J5Yqo9xXclo1T2B2TO+Ru4uUKeiq/EV75+QDzAf9HcwafNx
Q67LHW5NggAQl1sGN08QliQ2WLPF34j973/+ALvK15wMBVURqeM0RBqaxk0SF227
xCRB7FTVqBOaoxPuJpTRsiPmsPo3wVbOFblTgWhgnVTJypAtk1U8TtwSQuICWvMg
fTPXg5wwyEQzI5aMkE8uulo3qJ86AvLQi+L7JQ6aS/KIrmAjKFEULnvAoDCNS9SI
uLcwTn2rsT9xfHv0IiVBcHYXzRXM75rvP/28PDLPTMXN9AoYPVZpSDQ5/NE8uH+j
7Gu1UYFlTl7x7M2qjpirfcgrWcVZ6c2EFtNZHApTzjWAiot3b7hKfxHI4VyZ0Dwr
n4teVJrfRmZsQuPnQM/NBEPNE3DR2g2rJjxZWnw0uW95yMKH4+kEn0ehAEF3+8PB
psa+tR9u74TuisWCFQfUYTVNkg1syrIXmGsLbgYoAHhuFs3L42sSGTRGTmf4mHgl
Ffqmua02hyvVf0IJcz3EPbAwXpA2vDdFAJ2CAINWPFS7HTzY3MVnGfnmrA0GjqqT
uekgPT5pHuORnPVVbGOx7qBJbmQBWKxA/HAoPHTB039MyZjztS3HaWxifH9JwSkW
IAGqAGrvohPaImUd8JPsz8+dIpCLeLTd58yM+LAcJh/cRGGtMAIcqXuADZ0wMQxY
Rda4P4z7K2f4DNgFbK7A42oF1iGSY8n9JoFEmTp8E63IbzEG09QOADkfhm0x4UgJ
0qnE2FXX3RkBjqqc1FuPVW3LleVT/xJoWslsKMbV/C13kkke7tmD6/Scnn4csyui
EbJ7Ke4UFcJK/yV9qeuEaNi2imxRv2geuey963PAxWEb1Va4f5WdB4pNRU+I/76E
nI82RJW0Eerdocb0gAS82Bp3z7PiQ+JU5nh45pfvjoBEzCJMGSE3JJVZMJYrScT3
Fv/+/S7M/NAfC2QMqkemXPsusZ4lZ1vTbYma+85iS89/uWzXw0TMDxbwhWqgiODJ
Ix7XNuImztHX6HTLzDDZVS6EvNxmNZmpyJIks9eyHr2T8LjflqqeyyRjcPW3ZfAQ
gxZjYZGIhOV0qqRG/wYyuSgG/glvxJfzUKg4oj2RECy7b2aCgXihZrTohWkNkxVf
pJrHLKfCDBoEqqUKNnzSVj+pujLSihDE+7P3ttl5Cx3XrMy02ZPz0g8PYPf5TNR4
+Jd6uYjSY9z4bHutspGFED1O0KY/mR5+12o/E749kkxZ2E4+KFFgNfsk6P+i4ZyN
zazfZSKXIqaTDqU0Fj6dVRrr+GkxWJV7E+PwyUetoVAGtncxKesrBwTJ6d74bXB9
JJZZbUe91NoPAtmGd7pgChjRYpuUUHVnkArIFsFxgaZ/A43Vx0mGoRV1bneqsoDu
7PObo5sWAMUd347NwjuX6b7nmjx6q4lEzmbJpuDtP20ySgvki/NqL7U3wDroshZM
8twKt7pIUHephG8aaeXmkSNm++d9R4D1oF5sEnKHfqn/qfGYm2KbCJ62kdGco77T
0RbA71wlPqrDVjhpPEG1rqaMNVLNgG15WhJQ4WPMf2+diaDyHBG0KoW4dL3x76j6
Xi9uZSBuuqwl+syK/RaZ+8TWdHT1VR7tevYmjAKfzreWQu5IE5q0gDKIjnwuvu37
DRSRLs48WIENBJJpfRCaH2dQaIaV6KY85QzZD8SyrsHHTRf4Tfds6Pyu6TSmuCbU
+k26XGV111e9+2vcf0kQ6r3PanakcGsGIuKPAxw38lv71ioUGJxJapZDOReoikNw
sifY2+TMeCF7QFHAL5RJPGr9bEVwhL0DfoXT090XNNLo59psb90+nNib8akQgFcH
mUcfv9I3jcV+ZyR/czFdOO/3HHwFTTiooo/cBBLKf5T+CpAbrLl2tqyLUh+UbrjZ
kD5+OqMXpyZyOsCRLhLQoOB2/VddUGvxYxbRJ6UaO0PfnNrUntO8DFtg3aPz6jpH
gGL9VbtapQ/VOshfeSZ5IkhT6Y1EdirUVYQbM3dLoZU0ptT5x0wGkuGjXnINvhSC
qMsSfQhuOdctIHbyytjBfFTUvF7wnyX0sc479cdin7+9Nv7PU6bbNdOGiby1Iw46
AEEW7ULQo3vjLDgOCM6AQCSxpMpbzWGCcBDdJqiu/8YOFpuwnjiMcldT24Y/6boP
fyLWsDBBEpZuAhF5vizaTx8Y4tt5pkyOfbwdUuhVk4TrI1e8VtLq3d9x6gWBsbiT
7O91qpPbXO3Y72WbgzgzsPuUOsdDo0IULuZqtUnbkfvGgKjmR7yWF20A8TqP/8N0
yvNqZbHypwXkn9MlPuHJDY0gAsGxR4xlCR5un7lyoNlyjsLy9E/VpZhQTLzFPzOE
bioSQP3/W3Sh3qxobZgebXSwLHhIOqGs0T08KM9UhRVcsGpZAmswj3AIp8ktytyM
QfvvZHDBfzay97PNgu2H3zy5o40yYHFFfic01eTS1QizO9w2AMFuQBrDXmwCA4fn
2SAW4BVQ3JV+b9/UXj3cQyZY5AxYwUWdgCWNLOqxS02KL/HFxo4OTAAtm1M2e/bn
Io0esluKaQa3lm7nPh/BUx4HNjazqgE9vGP+nPbr98jg0HaXHvrwEpF7x5cA/6en
N6dY57Dw0jnk3FMAsMFgbhzbMliCkbgyul2KwrHD53mAUqt/KFecHch7fs+XipA0
Wy04Mpa70zipo6vrX6y78lXU54+YHc/Pv2YeXtsYqTyIWGf+s8FS2qZ/3rUXLEm5
Jz3xzf6Ua7oXWRsf92H1Tm/vbvyA/ait3Yps8c01HNKiQlGG7MNQ01U0X1Tu6C0O
5CgDWsfpsr1EUZ549aXvk/UV6nQFvhMe5cbk4nBDBcF+iY6OMypKYWGSrGVgzPMi
2ltj0aGWRBSeRgZwOJqGwl0bw4nQgo9xRcWYG3xScaXAacRPaEczxaptKV5eJ4UH
ONs0kngWDuHaXu3g3ah+cFwGcIaiqthuj6S7dlbjHN1zs+bwu3JTrTaP+hS+GgKj
STR2Hkpc4xXfCcNS1RswhkfDJJTDLvHFX0HYrrAAyJkPGsnUYLwG0J/Bx9iwCGsI
0erviWoFNjBpxWkorUWNxVjwyGoEdOBFPKPkuykC+hGow1kke8nY3/MWc0bnUXub
UJqxEKKbORdqg28RQmGHAdl/Kiv02gj+b3LiMfL4lY3LjjOPJS/WJcDDhGqMK23T
M+64f3d3DKfymRrFODd5kCKdr0bhxmVzdm9mTHwiT2BHIHroq3cmIMRZg/J5ZBuY
68ojdJpB716tEagHlhINrnMLYVgXlPq/FA48wVy8UNp7KGUl4slZHJ6Aenyilm8H
aoN16Hf4h/NAU/bRXx50Qql4f3eXlZaxfhMOGYeE78XcLP0tMmpOJ6Eff88qF8nS
nGxBAIU3j1Mx1mdBdRFjkX4Anz+86nlOnwDW4VtpXtcdiIGpM8QxTrFRLobo3BHD
wpM6+kttCLE/CDO2W51Kh2+Z+Tysij3dvZOB4iguh/Feube3LCZUx69IEcYg527n
kpfNQ8PjxkpmjaRPy5OmRj4mhkqlFRUnn+1nlBGVsVO3HflOgoPjZ9E+chc5Ri7/
TtRcDcCHVE0V05kA6VNQR36qMPWFI59unrYHR12bAt6TXrNpY4PaSGZBFeXSALUC
/Cwri2H9fHxY6HRMhJwJptVPVvE89mENVDMUuwqIAtSSdZMdBcPykKrInKVeWPfa
zWxQvBlwR8XGPhg4V5BRSaZgXxKYKZmg37E+8aOVI1HoXnLZm0+2OyOxw9DRBftH
LPBWgf797JyPu2owtgv/fhBnh/90DR1U4KwlzNRqdP99JaCCUoV8uQxjU/2+CsqC
u4WkYh21uhHTM3jn6sA1XDcxAC7P5lMnXpY8e1SfN07o6rSshKZpBMdCPNlFHkPU
k127cuMvsZPhZ3qHrnmF6bR7KheiwEZaeFIO0LyX2HQJcM+3Szv7uPu/lclPKg6Z
PZAxiYYOP6tbWyUma3ZmTkK95vGyyrcz32LF054BKfun735hVn7Uc6254HLk0vQ0
IM2tCbY3tMmIf4yj++zqNpIcka3Ewuqtuu5YnrQAp2+1W8xoI5ETYyedX9weIrhm
NyU7Dt92tuUsOVE2XhdfELHKkZ4uMCmtK9VS7rRAp+Hld+ILUrmLX6CPBOV7fJyb
DUE5VYhYD0S8rhnWDJKcpGvuIlhTO2dBXaTGD2MJEwyCipvJwxdn4NDneQKrJnA7
xLu6dCS9o1V/Xt2qcH2Mo+kGVPo3B/slasn/G1eIPh3i5I4eNw/AmmfWNRmvqyW7
8ToR5IV3gfLrYtEOJe/2SKxEIrMhLocPblWMZaxLn+etEnHJfIrfHTZvSkRDFzID
q0FZuXgE9acNKyJlK4p+vtSkdcQU2EiGctp0zSkWXNwgQZx3D4dpEbHcmQ0Y8rR7
98niT5i4JPSm9KdQ+BlPcweqTTL1VemfkUHau5WNYazhfrxCO6cftsdl0Jm3aguM
eCTGHQDIN5nzghfZqWdmorOoAQhCU/kpcS2AL6qgywXNPmpxMHf8IMF8tNhhlxrU
R44Og/YNRQV/DlbWKWgcOizocn+77SygABkS5ZWHj0Iy1rzxPhCpAMDV/g/z7geU
D23rNfJNd8L6449Jp9vJIEldxuTDhzcwxFJ2zIUyKRdjkFbaml/AHjRCfqHQMUUU
UYMHxJy1SqXaLTAmS+NazxRJm+TC3nWnCcGgaNIgoVJWmBT0cyu3245dtq7eNOQC
WsY/a0NSQpBQMrSTeLHL26rJsIlkE9Zfcws1ulR5SoevNcPGJNHHEyz97nxiXPJ0
JjxlJvFEkScfLehAW1W0kyGFGRCqaBYxCkaWvrJOvLl0J3DX9X5rJM3UraxxW8r4
bDfVQ1Dx9e4O5ZIEaBJGEzhQoKT3RX1vGTK1YChmp14gxEpsWRl9lB6iLtFCItoa
EJxaOaqi2CF9CZrKZBGe2xHR39muUURiEkZWJdww4ShIgLaiaUnio48eNOfEurhj
si8m067A/jcpM3aGu/F0mC8dN4vuwps9xazRCe5Jr5PZmLo06Zk60hQRlP8ul4JL
XbzsbcwkIXYTIUEU5ip4CrTF5zvle1gas0hoCeehjwCtNumYuUDM0JMR6nQ4eKLo
rGAgxnKU3KCEo6cRrAQhY/Bq9BfwEkCGRQPzybR23FaoC4kHtT4Hl/M6vEghrbA4
dC9WU1qMUtdvLV63teDi2cJmBJLH6CrQCP77B2Ub6AFzosMY6WU7K8/o4wL2ZzP0
YoSprGLi8s+tbn+rMAyOtAkAAYp9Tt9cuHs+0x9iD6er/qt6SvdDS6RnbyfyxOWS
dJXo5x2wb+q89rp5IW0G8/zRUVr/mHGRdemWBbqiQZaf/ymtBA3UXGGEXHIqiInS
kYQatCdJR9kk34COwx61dq1vKtRytY8oBLvQxoaR9DVkzEoXZmVHmJV6oB5dzO8H
i0mq+pTmwNki+AvvB168XJeIZ1EJl9ufL5G0IzhsrpSfqeuL+y6QAwtir/Thc7SP
Q9daOlRtowcr8tR98FAn499nNb8JHg1t1xGcuzOF6gkcCGGeKJBFjGt2O/b0hSsP
pov8md/wIzU7pzWE12TiCEmDQQDVFKflVJUsKmEo2jQ9tdaTFcftGTY5KEg7MVZA
CV/boOjLrQkBpM9jXU3NhI7Fe21nNpNoiVsLyoYTsnPWeaG561mANv/KcMmQD1Ni
8PIfcWUE6NVGYBu4hFBtot6S6pWokOGrABvTTI74dJTXL2Za/VUio2DtrGS4f7im
1cELr2xdOBpFUo4HY9eQO1vV9uYDVjaR4RrYc2y6nN9qs6PioYjYJJxpW4QsKiv5
6yZGYFG6m70mdmMWiMURY+joXgFXwSpAeB8tyNDZ/wHbRmc/6UqfmK+ybT3AOdMv
qWKFgPMxR2UVJ3JO3bHPYFgnEyROU5+gAR0TICJOkM+COql+/8Z2x3pJNpEYyh6o
eXWFsnllr8AtGQQUe8xVzGGYzpsCi0KOYs1YoWd6ooG23z2ubDXXF8TgAlPPWNiu
npt7Wg6FCyefCkq1Mf8kbNnO9psasX8SXoXpRRj1WL62QNLwQNlL8Y3/Vnm7Z9ui
GkJ8saWx3A90OjZGm4OwrKWU25vyFQIu61b2DWnA1Ojbsherj6eVcQ440ZNEXe0c
DLXpO0QJYa6koi9y56XdRoLXJv/YzF0miIyUzH94MYI9q1A8aBfAny9j33+IgHPA
vQPhKEUoUrQADjFQ3jMTMErLWPDlEYk5CVi6IGn8Cy8UdIPCv78bWC1IBiZppn3u
JJOnXgB/Opr2EdN8P1yIhxEf5akuElIuY3x7c9yyCCI4DcY7ZduyLl1LqikT+uDW
VnJlKvfrZ+e5dHEvs41I3R6m+d/W+nRKrGejClighrVk55RQUd9eKBJA51J3WhYP
Uf4C4YyGZl75QcG4lSLotFPOKTjrVSoZ3JSmUYcJ3nR5q0ReJJA+TyyyL2k/2ySH
i5ZXeW4pczFzXk0Nq3hBHPCdiUTj79oeZtrIB5g1sLgEjyuZoucj570kWrSW8Slu
9NWrAFlsrdySb/ZcU5qBNaKJyct64fV3pnzXbZz/2FwrL3S8QA9Nk6Jzgx3A172h
8M8b2pOCvBTE3bSTNsoSfwb9u6E7kgCSL0fWYIlRLBc98oiFo7l0mvE2x30DEZP5
T+v5WseZSoBt2Q7/4zdSXp4rjPqdZNXHkPQ3f3WHoLU/v8+LoCqITN9RYgoDtY6Y
KoE/KSPXSrN9cYt05JvaD1x/Q9Ta6s1KMwtj29X1nsuGfvDgd6gg40PTmyT3fTYI
+BLAj3tla3szlyUxcbYY+NcaOdIKlBBpyc2bWiRpVfvPNEw/m90ZUkbQMCVyOBfK
TpfuBwHiJVxS9gzYVwXa1RX4q4UO7WUPexr3vk83EWCplFtd4d3WmtJKgHkNAhPF
WrS//Jbwv8v4Y/M54bhuMwmqthdkIUscmV42DTl0Xjnf89r11I7U6iN8NYKZpvkz
TD1R8mvSd/zqqDGcpaCYFrcsLBbdS6/Q5buI0lqYhLpQKnraLWxEy/6519ep5nEL
n8RJd9FzLOaJmyeWMgR7uI2GLS4ncd7ZiqaKou/fWHZyPfgiETFPsCj/xOa33NQv
QHEcgK90B/K/3H9njJCgLAJjT0D8Upbu5tYJ0pPTgTaL2HUoeyKQVB8MVBubmLiW
RUtmMy15H51zzLWQFDLWVKPSa5W8WpCDQr+aHgWbrRFVHPSDaB4VErwJhlXCNLDi
qk3V2Kpt7e7NmEa8VulkMwklg+Ly8DAyxuaNPEJdx+2FDbGYNvHJ94w4H8Vc+3n5
42fW+lArx0vPJ634S0DDjX71yHRC3wNdTjBhVJZu8Jqfm8dFTPSExss15srWRyZj
fbxSnByPoW2tbl+rlLNpXsp/T3M17xjrtu6i1oiJo7I+Jaa6JD9F2YwfMsL/Ybyx
J1QnJApJpye4zTbcEgwdzPqU36s9QSPrxyHqa+wIBBGFpTObfyYe5H704OPCMmSO
TMf8XAVaS205J720LTwI4jkpyUNl+YSOh/cUMCHdV+C4yjZTEyUGx9i/v1xPDYM6
CrpQ+//CQQ3TivpjA+aZ8SGQ06hRu6v/v8c/5rS6WbojzrCUL34AeO/1z97YT5BK
Zpg4XclizeqMu64IDytupo5jQZ6P3b1Tzk0OzqbclRvglSEtqIDMmuGbEp4LRyoE
fXj/cGkE5KhcFuevJFGVWFcMhsbemOuhx+nuiCnB1jRV3Ah8ZPQwlb2Kf2an2WpL
NZS1l0D8AWfilJgu4XgPLHrQ7GwLVK6b3RVOD0TvZiF9axpOELGwS5eLLCD1LnQX
4cKIBQNlaJLbxx7ynWY9nzu3IQygxQucxlQe/p2vGiQvWkhO6WB+1JWvfVGf4zQT
5mo/uyD/c5S7nauSFQE3Oeu3VzFGvJoGuGkk4ekvsjgFvbhvImsH4f1qOdTJwpLi
jG8XHFWIAHzBiZB1z7EWK6b0Zw5VTyx31bfwC1dgdx6qu0WfaWYczkhfaC62upUC
yVyx5ADPDlgqHv4ReGKjbc0RogYRt4sBSLbrG06DwqpNicnydbTQ1dDC+yL3kWs0
fgVLKjx+KCBDbVxLf9sSGyi+umxM0e5fqjq1F4G2TpEFjYFieumNgrxh1eSavUPT
X1fL9p2uCe/zfT3kDv7K+szngnYjtUWRe4QPf7YfKxIIubYCJUV0xRxvpNFKuXUL
dq+kkpqcJw0u/2OenuZoPJdw3FzhsS8OPy3/PAQJnhrYKhPpM5dSUrEpzuF/L/X1
Yt+1DlgiQkb8Yf31j69sblykIw4Ol9pigEhR+xzwWWVCC0odMIO2+A2uO9KO9xvf
3J22ki+aFuZ1PM2t/OkMUepfiZA1/tqCeYFcOAN/4MhRU1m7UyL0L+uwwX5Jh/H1
J2l0EE61nw/hhRy6bh8FO5ugbeiTOihSOLpCa11lzv+6KDIX2A0UTD2gQBsO5Gj5
Vsrw5XVxuoux7PXr6eDrPLC0gEcGAvQy8XLe1jIBDy576Q8tPzGmOb+DcmntlGy7
k3LeVVK0KfUiOm31FiFMyjb/I2qym7XYipzkhTQbvw3qbw9QF+FXDdCxtbWG0yFA
Bq41p5/vhfkfc5tsIHX93qZOv+NOFbTcaOOv37hS6GuT9DxcdP8QrrVKEuuf6DDP
XbPUxOoEUhTvS+LteAeF5Ey5Suw7BvMY75/fUrm+kvH0p9tgn069ZXEYSxZit50Y
0PjdHS7vSJ4Tj7c28l2d88i3kc6/NG/dlDycgw7aETO049lS8TOeyvW9s1FxvVrm
WQNYVUqh0+e8UEATM4o28l6anJ8nr8rYmAQUwAIedaVVrfj1onDAwf7dDpU8yrIx
CiVD8V1ByqWe0HURPAYx+qrLz+Ej6Z8gCmy7O8Ga/3o4Swl6KBtuXDlvzEiMOhSo
PsXbybWTweXiOBvS+yEeJVO6pt5wuKbvvpJuTUP6sg6oMxxcofajkvZXF/jtrMRe
s8/BVnj9f065f6Mtdx/ntr0X8yubMuAeeJwx8SZyk5irk5dSS4YaorpHi03wzTn0
q8Z0SEL1pHAQ3wsTWx+eQGZZqa67YvMopFTkIRAukEQqI0ijwsmgrR9DIqX6vfvO
nQk0RwD1F6ZHenoP2vrOy+PxqjFXBLy24LII1uzbUugTqOp7yatdPjE2avC+wsnR
iE1U3gED4/cB86IHMFPtoq6oHOTsyAwVSTrI1nELlIyMxKotXS+cTiBuFdWlcf62
3jaEV+IjM6H/0DBkS0zOBHXKSoeLaUAnzi5IBG7HlLHDHI5vlqb7pCB0tJq9bAp4
x9PhNR5UR1iTMnaT3gUdjSzinQruuZzy4J1LGOan0I4kD96PMadsz9gbhUNug/hC
z8+0PD2un1crDTLfaHqQ+RnbJtZIJ5UUE/IpaqfsehEi5yq1vXdUYWtDVlLNC7u0
w0H8NM6xjVcyzsJugBSPPtpmmO6JuJr0ZBhLHn/0fQIPZYMeUf+AjNI5W8RCX8a4
5SHHT5z14Fiw/IKLZE8/dpGUTzBT1nuML7aLNM6RYGTZGLW/rphPKd1rmT9fZLgv
8LGX3fwvtQ0EIx81rpVVazlMvOCQzJvABKSSOHOyGoij5dLN5j8sTfOGhlAaOHaX
dOlPwinNVW4M67HiPbA1ErVuJRUka9khr5D2MNsey+2xt5PZ+KwIH/cyXNzrv/tP
x6RY/PQgIXqHFrZjD62qAdnB3lu15e3GzZIP10M1LiJ3DTcfvq+XN5VQne7qn0hi
zF4o/iVEQ+RF4hRsbJe4G+BJhHP3i3VMPQs47XHluwa9q3UwBNJjVK48LkDjR8xU
tFC/f8ED5k9wqv81EaDwlW/025lDhwEVYxNjokbWG0VIEUNBQmXqxK3/ImrqFbUo
NTiC07zRqowyD7p4oYxfuC9wZa0xvVCeUa5ynTWTMNn/gpgYscRKaKUvrZTSmxPF
ncVj5/wgCmcqwfrKl/vGKykojl8FD8YlkRPMKW0O/eYOJ/OxPpD3mHgnbMAAmol7
DcWPL5Vlw5Al1vm0xuTAkto43UD4zSbDyFyPV67mmtcf1HDDU0eES8hkUFyRcm92
FW6Tkoz3ZmxaYiiYMQuOntbGDjs8e8wxO7jPwZnOq6oXfLYRsFn2Om150e4YDVY6
mTzfUFJm3PLREMhGsZW4mKs5aC/rJV0eeB+k+3S6Z5M1olnL2OPG46nz9h032E+P
9AvMQEvvq8gRIgnVISGOs+1WIFT6tE75Zf/joW+ZQEcFJDltd5z5JX7xnYVKMSP8
NmnUHO9uNfepGWF58EHT+Ln7ltVQ8+o7Mo28IopE+yhX4VMUi2nan9LwIzpbAeC0
OGu3HAviZWDc/9Y/j5pb0t6Epqm4RUP7bceI8j/KZm8nbNXCZfDwqnItzGtTIU1o
1bUF01QErICY3fkZ3a1HbAZJuJ6uFQRHHnYs31hcudX5TYKVnM80U2QmHz7MaVto
OtWHI7ZuFWoS4gnMpNCMXEycDDOYDY8SnT4pnrsKGp1OYvUYy6OWh1L1lsjA3MK9
bFIfmWSVIRNV4jD8waN/gKGG8xZ6G8OKvBqo0ZfkiZBe5T0IxwWRQhnTTSWALvbG
DvRVu8mtWSJTwYovvfMxMKkipkBJdMojg4v06qvDy2Q62Y+yfITX9h7E2qtkZvhm
UbUodn5dsxSk97+0nPbH+wJeDYKFA54S80X/RLKftvAUOiS+SSyvxp7YyYoxx5uw
Kay5wAih05dpGC//31bpA7gN6+CwupT2W6te3hVW30MC5ef8w1jusOmVAEzjDfLd
obqLrr7SqJ5SxH5erZicwHYvmcDbo2QcNoA/oRrI1IAxTAvTunHbDKYrXFGhMfv8
zBM+kDqT7YyWjLKXrNndPPMD81Xdepny8E86cP6ivNZ32UzppeOn3rGnUW7boMQ7
ptwoC5sBAxjlQgPdpBpjgGLsiOFO/1XMt7mpU53y4vyrvSkEugGsCMjxyF1Yi57Q
n4Ka7UcHU7diG+Moro8rO/7ZbzpDpmzXjFsUZxJ2Qm4vD3wudqxUCYFSZxEnjuqM
e5F67d/xugQl3Ac20CHhyppfEGR/QUPna0whverrjSvEbV2LniDJwLwICnWyjl9R
/k+/mY7cLNS8/Vq81V1k4Rf9NwJBNmzbktRHiQJtO5dHQbGkjzklHvlNyZb9eSV1
fsJrV1u4LY4Qm5JbEV9d9bGYb/ms2P+kv3aqa2br50DXF+za4GAQvdwvabuYpyaZ
hdYSxJqSAFf7w3/WWuhW6ERRO6gLEqilZ/CoMYlHWZ94m22MTzQ5tbHHTi7Ts1zN
y+LFWPfrlqLm4LsCcHUe3KT4Zmtiu7fYPpQ0I4cvbyJs/VghGi1Y5KEYPu8Amava
csdvS0MKt3JQgBjuiDFY+UF1BzteAcw9gHTDyeshHmW4rTaUZ5FE/mOfEgaMN/V1
G6WDWNZybVP/83jUKR32vDBklISYD1vtUTiaYey+5PYhVa8hKiXfCP3hJGAA7QRd
gCeRvizBTPwx4SI4Ec2y7VKQ0zAthqaFAC5Fb38S+VeoO9of6VNLPgbJen+zBegm
ehDfy9fU94qY0z56HkP8XorgnEFkSBo0rfk2aXsvr3E0TXa+RfHmRVod64IkVkj+
fuwosBq1h05Ol05tPj9s2bhSJe7TagdZ1SYve1ScFVxzA65DamQojGtne1AsNG3+
npL8MVgIir7pnqqhHI6zchvCVduLNYtrCNJonoRXmUFovh0ETS7ChSmzLIebzqrx
FfLhD3WPo0m0lxUzX3Ws4mfLQAwjgkNAvtvSFCigvtIpq/fxHjnKEGg6I5eJhTWg
SEytggm2sULweuYOGfXOU8kl3TDQr7z4Bwj38pL5H40ilEe0oi7yH9C6arUIP+OC
+cGZQmEQ6/3kvzDVCIwXa2f9n+4FVvQjPX8oPEmuQRKAnqrESUWINhgCxZq8T/ug
ReTwATJOa9mrdRVaeZ4TQUz7vE89xUpV76Tr4z/IKyNVTUIRR7CVwGm75Suq4Tk8
d7wOTKk+g92mXpAaP6Jirl7WVnRNuiwcHLcfSY4Bt8EKut8L/vUsND95pfQ+lkm1
cAj6MUwGVuE/JcrVA8jiiGRWs+PQkVQeDDl6y/i/UTkfgc/bB3stKxvpN0rwxUDG
p7W5xBraUcN0EQ6FvrsWi+DZaU1oOHicrhOH/Ei1Btt+iPlKG282uqCNgmAhfDgb
QdPltej8IKhPKC7CvjmvXPilzYfCD684A6V/Rypd0E0ET/pkWHf2PRlUUVvNWBw0
hTrjmnbzuqWKnSQ3t7cENmsYSHeYvBHODhC57KE/tDk7MQtj047HdoWV8AEutCVR
cs+UO1zI60YIOY4aRdvNFwUj3GOTf7gordKgn5LxV0hZU7NMjdjqRAqsUyp6m1eF
oKPr1J+mv4MSYwYxiYiSaoibmR3FeOhNFeuR3CKXoOxqiskZv8Z8HZwsi/ZPFa6Z
gke/42HqylPoBWS9gWR0Yyh9dnvFC83IcYyRuCTABwBM+qNSpTwUeAHG9wQIMM+z
8tFl1xFj0Ak3fRvfoILVYH+qXUiN9i3iJLvNBelsY6NiUBGgKr+bV3zZ5QER9FIN
A7dnydFuzieBJZfIU70E2fOp8OGJs/fojVlhMfxYzSS6wXwDK2OK4R0Y/PQsDlEb
2G5TCDsO7t2MOvmGnhldt0NhI/QXtCZ+3oO5W62SyW5ylzfhIyP9XphRtEYgvvZ7
B0Igvbao9mA9mwO/NGlRHzbXQQyEZrP6MHv19kXOF7A2fDlEWx6ZJJk0XhkC5PTv
fRSXKD2mzMOK6S0+TsJjlbG+tmrOMCGnncNn25s86NcU95/btMLDhgEw5WPZb8cm
8BFyo4mUnOpQBNg9ThEOAPetvKopJ1ncyZF6jQs/5MFzzO/Nn8DIWr31LNre5UK0
Xk4XOuc0PcIJZybkjjlODj7ttia5dl7Gzoj1K3NtVJGVZ9VBmGzpJ63TBxa71rSe
n2O5hrdrmYXk3i1XeY0ewmgMNY2wTnWpQfHZKpOfgl4p7V1sEiiN+pw9IsYwxQBk
0cY41ZJrnD5fKb0At8WaHW+EGLgfgs0y+TfpHDQj/kwGSXsThlOJo8pgXT9Hnmai
ELFauagJFoNFgJhkydYMYsIcFYzWeoYh7Iw6bmPKi3ShcoI60HpFKv3wusYqTckY
WL23vqDqnufnkRTx/TmVQbztt4sTXlJKTukofsbCPeo491PRegG50mB6a4S5uAhW
39P7exzwA97RgLPhUlONUzuFabrjuYsy4Dk4qYThhYoVsUTla367G3InY652xCVi
sQwecWyH/HYNGoh5nGGEJL6TQdrAtoVh6uu+fCCa7fBfIR1GSwasyX+hJtgCSVRZ
1dDSgTjCacUPF0cOZWIR0zhIL4JsRdqydaXHPLFLZ0iZAWEroLhZEtIn67nc16H1
PDnTenwk8P+B/avMQHDhJuR77+dnOrfxj0TyFaSS7iQ1Vo3NBa2L6bRblQxsRr5U
+mS2i1PhQDH/FfRAQmjTzqARq3e1N62eymRo4p+2qRUlExg+UpIvI33HF1WV72ZS
3LjJT1R64Z1g08shgWPuoNLweD3b2WPd9C1kKmz9LRSfqQmix5KqaMp5kMkRs54r
cNhHbpMgp4Lc8IVBAA02Op0xGw3eaAl8odkiXK1lIGHYiddNCgjHlNOKrxnakScf
5U9RfyqYFYBMsb0Ek+Zxt/uY5d0oSYlUb5rERTuQ8FNZN9VvndJOWZAF8wX33PHQ
ngZorjlolJUPNaXWYHVzedkwDXGqgkd7/w5sYnTEah53aYJc50hnnj8aKJ4EZ6Xc
AQlOTF0qwkPVn7K23Phz5S2PnyxUa6kPJ9dcBzwqeeMc0CaE8WX3YHrVlZWZGdww
7ejMPCbtSZiQKrjx9Ou0Vf3M18cbvzSw6JxnPAsX61A4FW4ziZnClGRNMvxYetIN
Vzzkax5czZU8MHAfhlGEe86S1zWv3VPpDnziEwfNbccAiWgurVFBNFSlSu4BZH4N
ZDclmKJI/3p0cnMrMmhiDHbz8FaDlHv/H971RzeZcuEcnfwR7wYobYsJwqegr6UJ
MVK741ZxYcdJenYmZDsoio/21sCRhHhwYhZm0SQ1HlMQLwLWhu07Xf5ysfxtg6cO
cH47mMLGlO9zRjM3Ob9z8jQj9anc1oqUibCCYtRtPz4Df3NXXrW0ESh5ZfqHo13X
JaBcmvSAAFLrrYQwryRCsmbAdBnTtGrcAP6hlYs+pUh2pNhmkU4hJRkjGKQoROiF
dOyW/DDpLFo53d7SzwUAOl3lu1MmbIAzA/k9EomnkFYBqjutboP9Lq+1kGPb6/vH
Zd+LIjI+F8zPfSNlL3acmVzqtYV31omuIk1UAmxCAIyRMUkdukeNxLzW3FrX9Pc3
8p9ElOCuTF5s61zAptk5M/80C+c4GAtGnrD+54rkYU4xBVPqW2tBbe9+F0Xfj+VH
DsqdwcnYtOnWF+O2vGf2rJSV4C+U0rO3R2E0k94I+zUwKnfYlHmOOk7nNqgJ38yg
MDznRBVfsjK9Zzv/lDAYNKjLAiC3nV31oAAuHCllhD6SCB+ow8EDl+g2rn5Mfp8c
9LuL7EYZVS/76yUBGeL2OG/eNLUpv2kRQqntW6/audwiXurELEm+xOHqjBY8RLzF
lQ2p4PiuJIO5TkdGhjOYIaBk+h22nBuZeZ58OevgyXDanw0ljwPkw4+7XwnIC/Bo
4LkrE8gmHQ/2x+xPZVucgZ/4wT/w5r1mcvt6XHE1TtN7fy7SNq7B17y1QTjYsd+m
0BbREJayrs0of65PiS76o6gtDXvuDsbUO29dpsYoiLHuzAkbOyhjwfB5pKMI/fTr
AXWerMopoAsLRPCVppfMvWvWR6pFeSMzN3eiZbLYfvtkTW1hwWDt2PsnItIrShsD
NI/bMfKAWz3S53WID/st0MPMQ+arpsaFI51lMt5GXQh58C/uuIsLC/2gwjIzEx2W
CSKLZqPf2S25TF8/0VlC+rW8ignL2Yqt7ud+aiFn+yZNrZqMJNnMAepzfnWHLAjU
UquaYcqp5S+yfybmZyyvUHOFIssjMOq7DjHxqkOgsuI2qSLvdyhK2y3QndTS8N0f
nMZqMR3vhfXLr7YDqPdNNaA/5JXjPpQYfh9E/VJcex9x593MBHyGrP2IQUuFCvpQ
1keWrev0JsAQ6GjBtPfwA1MIQQ1IwI2NIaEJmkEadnoY7DI5PJvzHeu0QVGFOxKk
+rUFq8TS1wlvqXWxSSKgyJR96m9j5zJjf5f7mZaXMMp4459fIM6Jo0kRA+Dr83a2
uM+K4TE8YIz1pBLIhXEs7yWWIz4vamTw8roHNuHVGpYA9Ut0zARgyu3X1bW/0EY1
XJstjyO/pz3TP5m4HKr/JonYASM7UAW1x6ZRS/E4L8zgV5Yh14Cp4mLz94BSPf7M
jZ2DbeS5rjtp18cI7loeW62t0l9JY/OrkJTICPEirGZgBbHMGnJx6/1PyTJ+I8VL
LAywgJ4hvFbjm4KlSWcTujJc8jdQcZmBxOiSpeCUSO7KI6oobLaFXCx0A7sMFrRs
XwW1d3HWUI1abMlQljb0QKwh36AYPEbWJ85SOqM7hJi87UGxQvCXapOPa+/0yTRd
ibOtjMWOzjYIW/qhJW/JKFctW87pKkMc1oXrIle4igDgSsG9I9OOIZULd5UPAI8+
Qv/BFsGWMso1B6GSn4SqKlaKq35TOuOhPsVADmyJltAtk0eTIps+BUsBduMlDCef
Jy7AkxeVuDc7Wy9KU2zhBEMsaPZDBPFLwlsGvPZkTsSnSwi29dhp6NyntiQSkb4J
fgxKfh5RvTS6mOEsgadKcd8mbeo3eIsALNVf5IAFQvIV/RsNPaRfD2kFJI4L//xY
eEOxjhx1stem9Fkw/wtpyqY8SlxoFwRM5DH4CpD4pkrtfgYa1dJT3816ZzmBxZZR
SrEFT9PdOy3P99aw+DeKQHUcieJpLbv5HEMNmqg2mfHFGd4+fLGl/RF+iF4omoaD
RJRmZUp1wFmvW2ju1MtcPjsxGrb9YLsTvpvNK40Vip+IAT3wQgbTT6Cxe8MlWh1W
uQF18ogM6Xl24MqK+yaUtAgZmgOthnNcWBsmpKSb8q+LGmCIxRu8XvgknuYC1QZI
HvitxahH8ZUSBTsf7V4Uwn7B5OibntTv67fHaHpAQoM+aFZYYaZCXfhRlzAv2kKW
7YhNzGPgvq/fs3zWficsU5VVlj0LB7QQr8lYw6Dp3qY4U/rWrTLFYM8VDyP141RW
HDsTlohnT01LflxxFjix/TkzGwkOBg1D/HMsqv9gxnh+d+OMG9vhWO0DD1ZwSNjy
3Ow+e8kJ4eWAI5EDH62VtPoW8iey4pzHPy2aMEtlnUbN1IKxHXZ4H8U6HXXA+tSp
BjkqZWIzJWnaPwzdTH8Z9+Gnw7e2dvor3bkJ17/xMNhEtbImNTAp+QZn8SkXkJy1
kCtiRGlvxM/fj6KTEQf0HCntJcnl75eULxgW8evlI581r9mV1ZUPnZRYDImfw7mr
ZMhVyPbWVYgRONFThuEYsP6A8uMvK9Rf1SfJpIiKPFBtEJQ9PXtSAFvEvK9kpVJ6
Rzf8zpoHF2cLVMQRaIwSxsO7pmLPfsh4JpkvQy/8IeQeSkquTgBmFCEHO6lxeODK
tLingMYEBDSISZ4iUHO7cxgDbtYaY7+M8ckei61mAi+02kqDKqXg8ypi926F5Zfk
1XqqN7+JqrDBwrdugI5KcRKj9ge8Gc5KIVC6dAa1Q98brGViqTffl0wLjzDmqNjT
NqjDoa8Ju/islikgt5lsl5HLlInn2D1WsPZzAsYjmU+atyexIu7238ijjPhNLE3v
QtuiSkps3+J6yrW16+83fnoTasS4MlpmYTcf2Qbh0XrT07XbJj3kkH7I6PDiCeL9
61wOasJnIozKMq6RzF7j/LxiWBzrTEQLKT4FEHqBJW5+1NStvpRZNXNBvjC9XdgD
e6zc+AmqroWgES1cHg3hSv80DuPmv/ifwbftPGVsFruiH+/G6nsR8UL0AEFXNYEC
0MHeESLDg8fRUkpfru2PGXFMF4qF5CKinrTgW1XpY3T3owBmDrpGOWyBvP5+Xkwx
6/w1SY/84ZRHYsFTWv3fNuumioYj5W8RvbYYHWcDFvM3PaWjZjI9hJYHQGVH/OY9
SKHOmOYn4IQvEeiVQ7j0qHyE72xgLo7wXkg0MIZ7LnjbLeVCtje6dtR1cfpP28+K
DsG+fqd+uMvW2cpUT7x4EuupzRzQHCVlq43eKWdDPdMJbJZg49ZfvWFy7PdCw9yl
wmPxdn+qBJ46xT3y8/fu25Rswq4fNCUhYzs1UXEFWB14zSVbCi1lmBIAuo0Flv//
gHyAbDRTQu/rEDF1cOXL8gFVcdEia56TSGNRuIn0U/L/JAMkOOhGBG9Gki+tOco2
wSIzukxoFVxbWPegRcU3UniQZpdu3ltX/v6XK7d/uwgN4/IwS2Fhg8tQfOXAt/Mz
bLMDmIJbnjsGGqt7zSOcSRF8nAlbwf/pjLwb/GhtEIUgn2qdco9oha1lMGMIRgDh
GRwerkINuDO4kLE8k6xLO3ZC6cxVGRjfgW8YfmzCc/1tYLsp5rqoI4DJcr4yk7q0
qeQSZNvNIf7H9E4Yk9q7HXh2u3dO9Ze/pK+BWimMoq5DrbMiObgaQ25Os6KI/Vkl
wb85DDuTCiD7cLzHc+5v46Hd0Sq9MWKvkj5ErgzPYoaOZKiR9ZlTaDaGaP6I0Ji+
/2ADVO5bWDIHReeR7j8vIxUBdg4iPofD+ppknh8kCDiX1hx9br9o/XMZoREIEKR4
ngI7s6bhneaxVTYQOn6nahFNba4/3V/C/Gx9Al4T/zWlMTuLc+qLHAy1MXnYyvW5
oZaHstkGVAyR8qE6tJYp3eioMFnMCkfUVReGGGKP5b6k0V739FvcPncR0XhG6ttY
JIls7HiLsVydK/N+osPvB+DDPEQx7GLrrE/c1uJ0U6VwMFeRbr6rTbCumE4wkDGS
UGa9daM/osxep1ShDnZJSE/lLl0KeFVGC3BTsTf/EDSe275En/MvM7U2BlplUESz
DwjMMTlSAHxOltTubVHyy5a/h+ToZBNktpE41d9mtD61SfZPR/VAR2+AWAJNP6oT
dpvWAW+gIwxIbk92MhBG+O74qzyAeiqfuzRP0txH4ARbydlGpXjXrS3eiRLLTmvJ
X16K003qbLbN27cfD9tIiiU86cvvgstGNg/wDqVvIs7EBmgBCa3k8sUGFPcJ5IqQ
siqBTuS5Jy+09uabEozsor6IrZuo6q7paC6skYVTYKmFMQo+qcxEPHtja0UgrplN
mNtYrqbKZZIFql7H8ne4+orcWJKnc7nT+p1hdxUcwfsz08QGlPV1v4Veb9dSZw6T
KRcal8HmXRfUrqo4vwNaaIzbJqExaFUm17J83ry/RbrSUtSHZc7+s+QbAgtvGGNT
kalUexyozsSSXzb3nXvGHmRK4DV76E24HvkhoA2FWiNKcSdOll6sX738bIo238Sh
4d1MPkpp67mw6LgFogQGm+8am5jv1O2QBB3MfApk/W2WOxwrwL9MjzRN+75+H3oU
Iz1QaNm2etVCcjzrx0ubncrwmSztH/6zkMux1XNF26N9aWb/GucdbXBfD4Tl4QJm
BvHOacDrwkbKgnrrbXUfRomsk3++RCWADx2AduPVVs/kkg8OytanUGpqaJUlgoAF
RU7HLV3lElqlNlP5guBtxakzdJpCwjUiB2v+4eLCdy6Ozv8GdWjJNm8eW3BSOIsk
zwj74fB4WvNt8yP2XRiu+4Qkg1S/INIiTq17TkyIDB2zimzrTc1EBXAss5f1v84X
vffy+RVCZNnIdKIniIZ7mg2Ocqxo4IBZZe5Cpxv/QM7GNf2MqCt+60Y/d36UvkNx
sReTEpqgdWVKKxBJUJQxnPG40rvrBrxjvQjX7LZQ2Vz3hZhraXBby/amftms0tJC
ogEiQpIJLHWoHer1fAZ6ZTdaDswGJGkqZufglBrk8o8l7M2rumZKBSwjWweq3V4j
q1X8QaSKSCnUvZNBo3uqEt7K+if30bKVWgl+S4CPHZxSRs6A8PLqi+iJHjmaArDD
g8+harMxDQGBRT2eKugWLDzBLpzKaZwQ7GmY9ecCdzKoN7O1bBdmMafI1aP7JnjP
e4eg3FSPsHGcXKHLU93KJUi9y4rgY/M6O4P0aqn2nId0nDP4LoP0BFZGyvoS1Ywt
wsw1j5MujGBqHFI9hnpthgUckWimr9hJ0VLX5BHwkKPPsSYPpHtn+3dBs06w07oL
UNqR9XPytipbm4MC/tOYn3HNpc45Aju/u5TKsIJht0uxOTMUxk5hckUyV0judc1P
gYJrm7eTwvlW9EnnTLGC9wd8nx41OACawE0ygbo+pyaEgleLZefmAUbPY2TAgVvI
8OFeiJCeSEXJvjG9boMtGyd8vwVDDctR0puJVSJThhGB75DF3TNKYVTzfIHkQcmm
is7yfQaLR/jI81YEhmM9kCYn+IxuFe+YdkAnQ91qgR49KY/sNy+g9UFJ8IhCaXK6
D/TMzO3WB+/ybbthf8w8kaRXtiSRpwx6fyt+xWZmNfpr2f5RSGw3IhRzFuijtRFF
6PZFHVwW+04tZvvAyqVqdOrtC+zjumUrEW8y1/ooq8RF9vXD7nqBy8P7JTRv0J6H
E20vyVmwu0bsxeH6upMjIWHQEVCRmFovRkTVY/hQ0QYJyYR5pcYqgh9zRf+d0/JG
NEuKXPu21Vom2QAUN1MsyqIp+FJ5vJlnZIb+UpMtewUmdPRJX/eopSigVNH1vlwU
zfQijM/r5nAtBCzCH31/aug+FUXxxbcFwSRBUr2G0lM/VR0nOqIZwwYGiScVNPYH
7/p1JSK1ppKF81KPvek4iaeZxgojL9zmPE/dSkkXCfhRNa3vvr8hSPQClDtYtplc
RUjPwtUv1zA081c5TtAjLxqSJdj6MGEDUQN1S9+em56g0UElIeXe7nz/o0zYn45A
gDqWntQi8C94703g+Sx2aI2opAtq/JYFDI6Ls3KhrH0G1QlHSKpcGHCNZsJNFq7d
6PopOQ2lXmCoOnjAPuG5nli3EPg6aVR9WLvSIuRaVkpotUdWfCeeEJoqB//WR7MJ
FwWrpN+8fXyg7cujTCa4l4QjD6oZAtCExjvWyxQFEwOObutHiQ0rD6Iy1FRyj8i1
U/G2lxbn2ux8YzQ1RZKMq2ywxIogY72eHDQss/Eb7xSsHuaT1T9ulsI5rWTZDxQU
RH+CtIigqg8xjIWe4tSRVWZ7wD7HAuwBqqHW/RiqHLk2Q1s9HI+PUkIC6JRvVhts
TmAyg6fWSVuS+Wvwf8Zw/d6BH+IcBal7sIpoCslvGHXO5uBmbrSb6tBebMIFdz9c
RvDlo/47yuXb3PkO2INFnAtC8SrU4pKHElxgAqEGFbdbDS9kV8VGNE07YUhF6y/h
abeTuUOQjbgdmKcbVnxc9ZEJXVH/KfnOIIr+AgDoJCs3FLoI38+krL4Z2r85Y9OD
hdlKV5f8Btx6H/7PWVKsPK/J2UQiIJNzeLSVBWx5oydhT5eF2qdl2rGxHANhN7oa
ThfMymw2mluJA5BJfl8u1TLBfIGLDzhdEUcqzrClOY1OLMHvPuEvN21ZGUJlhpHW
C0EGGR+bNmE3TT8q0lG7SYQYfZcOOrsd+DCYLr9OK7doxYmCiEIoP1911f3AbBC5
Tv7cVSV9K+bDXY8blkTUHaJ0CLAfBwsh/nuGyru9Jcf1rCLHvKhmlV+ZEaAAVvzM
JpQMGoGrfLnRmfKVEVuBm/dBf5ekg/znZD4iNAJTdKdLOiyC7v2xEHYArLvSLBnT
vaXT9U8XoIr/FUjvMd/sML4E48y4dhgq0ZKxDOoCmECJBFhXBLDsEMp3bCRHrDSt
YP3Q2snGMGxFYDYhc17mFl6Q7wMCtFCY4w+gHRbP3efDlTjpFBuwk0iD6Q84tpTh
C9idbhg6PC1u/8yCHWrR0hOSIfTRDF3ljgEdQnd6VmwWxXhwxZrg1wEXRhqVqL82
eij/nzOPoi19CW6da+QYMygkq4QGDnx5WBuRVKPXFKvwKTHxrcGxMYNftF/SWyRw
nUK4BjtQEfFX1fKzULkCkbjOnUOVgLh9cgtuLXT9zEMw+kCNyYfEcA2mj0TP7Cyq
LyDmhfBDFwRXr/0xW8qrkEfd2c0HlYdOHsBHCcax5uMUwoFNzAq1xcx0oiwNZS3X
Inqevfk5qWeaUrfT8Zx591NkxfOOWDEYnwXCB8h49DIEbLeDmZVndOVORxByYBWq
bDdNGbLu+eH5f5a5gt+Pb/h1SP7Z9V/dCv8pE12k62GWPfuIPiJnLwJNRwt5G16Y
WoZ6K4Xmez1KZAeyx5+QM2d/MzDznpcjtvwLDRMegU8BekPSB5mF7eZfgHwPXtVA
dA+5N8LDW45x4XtlGFPE9CiToVfT8QunNY8HzpwTUmhRccjbkq8fcLjno50D1ZVe
UuSPrWYlf6av5paNw1rJici5UFK6LV7FyziPpWfrvwbF/PvZQHjW/yrs+3TsLEkV
wI5dMmX7awIcAQscRWFGvviOSy+uL+tRFpjiXZW9xL/dpUTWTYZSj19Qt6GP3ucD
szLG89oVyhKMyHEyDe21Eksj+AQ2Bc6mRTgxPiTlCF5uTJC3N13e6LNnVTAl4Q5e
PHiyN9ygaZzyp23Ph+rPeGNp9c8s8ST+rDrX8J2wz17eJXZnUZb/9oFDXOk8kx58
Mz8GVqWr2aOSdESLcrCSzsIQtFhRsNC/MhxeI+8wifFOG8vCuDsxDYVlHPe1s8aV
e+sO5bj5W7KINtM4z9VtoS8CqCPvAAyqqaGgOlTN3n3+J29UyKByM5WDtxXZZ+oS
lUIFpNskjsqsqcB5YfIjqfBxAEbI5aQYlRLm9G6v7V3j5/nxuyh/vfyPKya6Hc+t
uOrbLgWCIvTK42woOW7fjL3cFngx69heElD5S+eRW268X3mqxIg9WMj8C+YsNgFW
+pNsPbXUK9QrD7l/rDYBUtoQM51noEri8DzsjWHBD/B9nOeAYnsXA6INFabMIORR
kFdWgH44z7H7UzDom1FAK8PPf7kA9E6yT2/EOa26hV8cfLcST2voddQpl8mWe71A
snAp6W3XWgBoV4h0VIwqCXTJHm5hMIjPSiGIkU07uJ+Gx0OkUqEo9o2MFXgy074o
UKfJGy4Z6Kx1At6mAYbeW2MZGBxrea0XQ9vphfa0P+elUi1TI9BSUQMcXJYP1e/y
GV1n0mNz87x5q14PEFqp8dgwk1NkU1cbWzAoq7yfyDqeV9hJMsp3tT1k/3tY3FJl
oDojTgnrhu98Yij5gbJjUGY/yX9bSYrdPUVECG6PuyttJVsK33bcJa+WvBCDv62M
jFz9OgwOw4OvcNjutYLkdnb0s/DV4SwHAQpGT2HpM8TT08WIpj0k2CymYXtesKn3
sNQhF9KVXLYlq9F/eP8bV21TF/AZiWLqv20GLESQ8ltccDFWdIenrV87kU5aveUa
nJVR4cw4LxmXKbLctGoA0/WFRP0aW1pZ2KXgMyRZcdNjFI4Cp3V/KoM7mFMvwKxD
iNC87WbTEvsQ0oOZYTgyOLHms6iLIu+N5pwS84SnTATQg0j0EXSHzh6H0zqiuDpn
Q1iEEw14IOs5dne7RdEnKSUYeaLtgC8DQUhIlav8qgKsOGk3uu0JQXFXP7/3lWWn
l02kG2DnGx0aryvEXD5K1CusI3sLCbSw8Wn/XmIurQjYHTnDS2pxqVT4L3a8cqln
CD6Kqg0Tq/MyZzTzn+fM/rRys7GGODgGnHqBdQKPcdmBPFh04qLj+kNe0KFFpE5z
aA6O2Yzg3vXLmMnFJwrlbOrbevgqjKZW39iCRpfTNNMW7aO/TrPb/482eWUoiG9c
WljDIzUFGbuFnwX75gxWStsWG3z2Kilu38v7pXPOg2IfcRZ+LVqPKvNwC/H0uB0C
sN0qG5nTS9oM5ne/NKsN0WyXMSKzEMhfwMcQGD4fkdKFY5weK6+73iNZ3eZhRlLx
39B748HhfkZfcjjVsSFza7PgHVY2nVYkxPmnuW0CytMYEu0XRYgi4TE2cAmhRnvc
mkQF42WT6a4tc6AJshXZmJ1Orc+8STekSNFUTsfWV5CiTLnJJJtCf/IcwcdblSWT
bzb1T1TgFMyKLVgVh46KFotjHBdghf0J3TTjmnvNOR7kVGY6/lJNlHMYS9C1y6FW
RIqH8B4n/37eHtfajML5yI4aLPxsVsRK0fODIVb6tD5d04wapi4V6UtEx0R85T5M
zGmX9uUfRO+zpvN5Z9YhF8Sos0CA4gJDezZ7c5yt+Tk3qNWDUmSD6qb6PM1EKvNx
MzwD6Zmyf6FMWau2CVVq1We4hlgs0tvpHyEmzFMduG2XcivjAJkkKggtQorKYvkj
5W46cRjR4okkOOiQ6o7ChdQtX1VJWwRiAb9NAaYJP6Mof73jLelwMLN4P3DLO9pj
U3cGyKc5O1+tTJXFXVGguCwghJGwxlyu+Twrh3epil2OoGQFxTFpdLw3sOwNMYO8
a7SRPCWVAntjcVqbtY8PPnKeU+uQT6vfOJLIBrWHDVM9Q6z6dMotIL1weBewD6Mx
S4j0480rkCkf9p5iKoLZqY/iIGhF9L0xk44nW56iKLaVIIkUf5J9sxte3lUlU+Zq
2JM94uBLMreVhec6T0HoSejwGQUTRh1H97Ioz1QbNm40USh6b/lWJYiVK5lZIN2I
q/XQvN7IyBPMvnRWvn01LVYbAgMw2JUSv9xjAOQV+RlDqByUfRof6kiBPM1MIg36
lHtOCPNXxLeXTWt0/AaIh37+fRvWWmx51xp5FzEnUsb3R6LSzvIDZJoIRugScpfi
GjuxRe5rQDJSKbb1uDKzR6hFzQWman7jK/7zhPPD+4EfgSL6AH9oD/71V+T3/Hqx
JYoNm2QXqDsIs0vTo5eAFNLGSK0gs2o/7ChWKXQnleFN4J8QUsWJQDop4dBf538u
WMfuN3/sTcJwynK0pTWU+dMPPHk87Rjia7YW9dBXv7SOr8cl6lHLlzuR/QcWWAV1
fZCFcHnS7E3PdnMJk6YM7d5X0A4xu9vMtyIqCi5rMSSanKRdX5Pm7aRgnttSxv2h
38PiIqf/MG9t41BuX99met6ToXl59b/Zxypc7ZkkAeuYm8iDuGjpUi3WiIcgOhGo
ZH/lPo/ntlCJbYJAqsAXZKU9Ww2HTotrEKexqQrxqGxmWbTIVuUOlbsdOwuecqKZ
ehsuH15Qe+AGQH6XhKTXha749jOP+kRFa47tBrT8cxwthWCU5x3UITPyAtl5pl2d
aZ/wT1NCHCXPlB71Px6Xn0xLMg2SwMqm+c08rNRj4Iox23PUm+K09kl6P0GNk/em
OMTQcCwgKGYMiljOu22qgHhXDqQxjHS2lxuenYyG1ZYi1po9GuDpfE2gmBqNoaxH
tiwbltuAse85pWOqWSoB8u9Ngfa389fIHDaBDRfkFkOaFAkSmEFrkHtrBCeOaW8v
hW2IsBI4p4Os4+q1TWIGhHWaYb/EkZoINPIaaagstI22H2vuZeVkXtMSK2kNmov/
laLa/bUr0MGSDfN473/0Df33scrlK/p1Dsz9oOOkIpYsoVoCj+2g5dryVLZQNhDr
3LHZP/QpBSg2GqAfrJg0uAJwzGVE7CBtUas0pz9Bj0LEt2qCy+4HnyWslfEALbMB
UzzfziLHfoi5bqoKQ58DMQ6tngN8Y3u8gtdnj1fAdYgC0VySboKkFL/GLfAysN5t
SIKIyt0mzYyMbG+tM/FlKwt8hQYwyiD6Xgp1uI42VAyEMQFGe8/VhqtBr599gVIc
J4nKre1u2GLZ53ME8+hMvUHyUt099xl3gJc6bdnx6OJpgbqVflSEMa1jovdcMKU2
kY64dSXntOysRoAnLwnpxqilzCfCAy0iB0wtsaHqODKbjamXsY/12Hg/BJcalEBn
bvIqX2FvY0Jbi00XpoKD8LWd4tucfBFRTLRN793GFwevKJbX9rzBtxXO2bejP+Bt
zN42GLObcclDcPBZ8YQSfUZ8pWBBX0Tl3MfICaH3mKM6o5laJOUxNx+OGCACdmhf
k+ADpjmWvfLOQqh8vJTvqUyqlbHfut8FIB+3CVtL+/YQFWG4+A98NCsbje0kIdIm
ZA+bQO6ZnLwS07vDRPIKjkAG5fWP8zyIuq8XBupBwFbMipHBZZ9gxD9epv/bt7TK
Hgl20fGBEy0sOCe/c3HQN0JRz/GpoN6pUi4xtf4J4G3sWvHOttgkg5cD4zEeVf4N
1leDo5kJarjvoDDIH1ITJqwZVPyg2YSBGK31XY+dTVQsLpUiZh9KvxD6THR2zGal
DGHr2G3QuJMo1FK6OjhSV7Y/gRB+d2K3SigILWXkUR/jOspoNd6YSqBPxpbnlt52
uamZxrkoVBxvcCiZY/JZY6tgukYwTnNsZjyvCOs7TrS8JK2b1GPiOWp3VF4zifLz
izZ2T+v3XMLlcz17tNncxrw0ZY3TdDEntR2QLFH913ubiEHj5qQgIUb+jMhCF+hw
CG87gl+0YghxLstMJDIDvPcv8Og8VZizXXQJlde657y/xgS5IVAN6Wm6yVMdQLSy
jOW2iMQAJHqf3foJtQy2Vtro91ZF9RQRDTDGCLeaR0igx+85HU1VKSqBpUzcoID6
cK1QWSd3lR+FbISAgmaGYBMVwZvQfeHYYpyIzENoEMjb8aDghIGTW1hDC9DWD9l4
5F9uru/ChX06CcJGLBoe4MluSnJKAQQRqKqdWEmWG2+RcPw3dtElOR/ivYvV9kt+
FiUdEWxeu86tch7L0qLom6Ct/IoDq8tnbEGKd+Pl5E2Fi0dOsPbo0PV65dpvV291
ggI8I6bCsdiHAjXWRl6iVBsEmxwsfIx+e+j8kcUo4Ri+4Iele4ysBspd1+TOsobC
VAxJt5Iw36ovsS6FyGr3VK9I+dTFwq6/bHTtf/qcZMxThK3vdvFoIX1CrNO1r+N0
zQr2+YfYXCzxxRH+cAFgBOMI2MOtL43Mkz2r/4KNHe+jMKzFks5Zb+j5ZkzuQLVI
9ja5l70g5ppL4v2arXTVZgRoUlHtfGdLOszJ76HW3lWB3ABpL5Wfk7NajPRggKOI
1OhRdjtTm/jKwmDQ0pLZOspPx7QfvZmBqMRORWjbbXnE6YkDdOVO96KKqT4uVRF1
1H1Pkdig5t0eH3KJny3KweyKYvCeB01SSG5/OyR/e7Ghd18WIRahf8p3SdxuT4La
oiXgEXIv1DvafMFbAh9ABkeWDkcJeHcqvxSooG9/h5ABnpo5TQOxVtjrAmQnHsF4
g/8wcZCOBzTrpIc/oiICNXidEcjOyC4EIncQO73+wSIU6Liga42DQlLHJgnHCsNa
UBR5oyk5XfypHiuGNBVN6zY/7Rrpr6FHmw4t2z+YanWA0rGkj9PV98YV4l2epE3T
vYUZw3BU83iMCdlXmGildxDLF0VNF9mwG2Pl/B9hcifrc8F8k2qq1DGiMVeyc9OR
JcEMA/YC+8gzVMJLYdoC+i0he8Q7aADMu+aXiZNzRxIUbxLiib94f4WmgVM95Lq6
YTZpZEplfWl/5eLZkGf5nX7bUvQ8TqqUhphYjCRK8fE8+CK0GZe2SOukffXlgV2U
+y1hG9o1kIi6SneffxqIB0ZVO/JbizJXMmqH9xHHxuJdyXZfyX8IIhPICkLCk8/0
R+xWFH/qZNOEDoGP29dpgoatQ4CO598Q+tD/Ass1wiFRn31Fnmsz1IFji/cLHwXq
W/ZvS6aTjJQCQ2PlUwz9nqJJbEub6/EU8NEwivKvniqrgdPcYrYq+rA5IB1jjRC1
KwuXmhoBaylPv/O5mPl/m7lgMJ0E0R2TSVNHqBPIWCH50D8dGOJfWUXcW22ecF+j
iDAy1JNREEP0kGs3MTEV19+Fm0ooObnajv6COTC+l9ORxGQ7MQGxGRHxs8n2gNCu
PLYzhTNXUWdMACaPobIcpbPP/tu7lbkjfHaBzNPP+vtYa9/21pS+X4yUrcESIUeB
c8RGl9hD7xJJjZmlHml1Fuk7ML2hH0jac4RKb7Xtvtrfg1gnFdt7HuH7W1SPFBTk
cTf/9LIOASG9TwhQCavLeItOKSiCOpS9Owxy1ZWc+5F+yOYb7kFnFLmyusjjkIoJ
xN72jfmQV7D/g+xrK5p4TxwC0dSkCJqoORMprXjn06+vTypZm7vjdEGXqnD+lLcJ
anIkiGn6M4Ia8dmLV7MLwBjyqIL3+ttcMV3cdrPIR7r6JOwU8crgBdmGbP+4RYwx
7TFwU3nWisXGUiPLOLreLrSUxJF/t6CO4OI3KZEI5W3jLQ4vX0bMAv4/Rud0D4Lv
NGdxBoKbVbDzrgqRD4p8Caz+U7JoltvwveFP64/Nf3hKNxOWln2F0ZjWuWLE+Fvm
T77QnKr5QFXq9xMbC4GjnlwcKD31sA4quiRdA+MV5xQaFFh/g5F33GEuN8NmyPRM
t96zDwxRkmXHAanhW227lSUoDBqDFgqCc2Jygh6guPc7jAMuZAKG3tzICd4oyRFR
bQ3dwsdyMDXcqar1Qw2s4Fna2n28DMIAFsBUw43zXwSPVHq8nx3vYmMUO3ybpZWU
+JGa2rmirgPsjid2CINsNOcDECeFpWegZZr+/o9eGYU4Qzu4hg6/SOewgj+IMYTU
jb4XCfVrmanTaQzjOrMbaHJk7MXG3SspAVF5ZuJXiKU5W8EgYlnu40CHo0YhD53h
HSSYrUcpg3ZQVM1Y7gBrhENB/mIjXJ0t8yq6iDR1N5SIumC//nj2m/7ymBDQVzo8
E99phEkJpNh0lpIp6TWF7Rl5uPy17GytOgPmfcA6Mhb31WEfWeSJ8tux/NJ/cjPi
tTqtTM0Tu/4wJ9tm3dx/dB1IVsmy2xXYHntrbtT9vyAxW2Ddff9vI08d1PZGzoy2
suFWl4U6kznFuI1fP1Wqs1k2dnDcJG9bT5UnNt2iIrXviHNSUJfqaysX+FDm7jxo
DAgWRcJRvTqwtrkPxhTRHrwCqppLsh5k98BoyoOBIYDaQ+Zq6yQZjUQC+NspFuSs
H8Kylo3XVExRcM8uOGQuTVAEoQITmmoCluygMn1tiLaR6TgnDCNcQ5m6cyxsBCrA
l99/YG7p+DLQT1lkZSjx6wcj3pBCPMvZ7t9NmMYFSMJNuq1GKc8nDcVeMPer8n8o
enuTS+35+3K27CAkq8lNShYryLWLrdcFUC+084U/Mh6kElYuyfWKpXQKnbXQkRb4
ClArHk13uIBJxSf2KqklibLvleF3MAxSD8EC20Cxyack2ivhnl/WQ2gRUymJeEZU
T13F56wHa6i2ZTNQSt1gwoUkxC4B3hyTt+pHbdyF1c25c94ResxSd+LPmJxO9cNS
HoUlxXxl8Pbcfjq8IwcoHuT6D4YKFo36NgSP2Yo6DPmGsby+q50J/PCTzP7X2R7S
YNtO8WI1wu0XnGYyg/i8Eofv9G5Lzi1ezNws8R5nHF6/iBv4dtdtlIGMq6E7p+VV
fCkWd2Hiw9uyDWYfmtzgtSHTKWUuyyaFVBQ/hNVksbHjV0zYMzW8tyRgJ7zoeVYf
3uz/R6ji8NwiE1YG1nfiopYAT2SL+7QTnT0XVyeqzQS4qLCCCB4LnASmze4mwOkd
AgW868sgBrn2fo2TvAzFLygIb6RsYR7ehDgPq1U3SaXWTNzjk0Bo80i13w8+MVG/
vEw4lmCwdTnySsnypl5ZZl30O4rOn4FtvQV52P3RRRygabKuFyG/dScz40ittjVY
NwXqZx6pymxx0AkbLFiSD3633vjLMoJ3DxNigfbB40JPfx0vVzsVDeu+Yj4W0qfW
44u8fAkVrhfQTSoIpGYQ/NfLtg1d3wnmTNUiTAq+Xu+n1FDsX1lvRTDd2EOA9DjN
r+vdFOVipgiC1AYup3/ppz4s8HCvLzxkYKfxpmK8+o+FIKLJ3oaCOb3qi2wVZ19P
3zkXFd1Cu62vORPlpzmeW8Cp7wdenpEOesvevqTT21o30qDUDGL1Y0MqZYtvHGxF
B5zqBhJboAmTFYqudxz+YyZl3jtZyKgoikmGbAMPjxDDNObmntB4UjRzkOMyghHC
cUx+dz2sj1j2rDFDQoGjz8HSlEnevCvBWv8Qe0B+PEZzwT04yb/7Cqjz6qm9mHjN
a66T9Oga4RbksYNilHiUseSiRWwAlQ+yQbtC8Y4yRUa0w2B2Y+9IVbRpOGAVF1w+
7/TGYwCAUC5kxX3mCunAEKTxkkTckxs9OWx4RnxIokZmKoAPlMvLWM8ijbN+zMdO
uuGIUnyJ3CCZi7rPVDfQ9N88E2JrCITon4jRdzNjW/b3GgiHnFMEu5K+2h1/5vhO
QwC/gxVBNcOeu8iuDjzff8hLINVEJNQyvOAy106UhGUmewNL7nQCQzuhnox/lyHy
SZ3ScpXuIGEe8SUxBijYA9GS/Qd7l9scDjp5Q+WWhl4y1z5FoOG8UV+hsy1+vcyM
KQcGKQwaPjrZ7axkmjfnfA2/fcSqbAPjq2dydUth/9AfBlR6guauozUxjwUndnu4
436RrCfUa1Oi3uE5GdmO+OTxHoYV4hiuF3dGX4fp59GP4mClUopFCl7Ax10OlPL4
rxRqs4Mkf9A/nG4tpq6gU4besRqJQNjUP4AhpeyzyEopzN6/Y4MgPdYl/b1PuKwb
2Ak3XxJFJYlBOfx4BWzSFvbsjuOOMz8pmAPWvuimLuAgXqZ0+xfjYwKdRLjWAk+Q
seHiKlniTJIS3Y1fKn+vQmMjsAJvprDSRplV0/ttLPxxOcdu9Fc6My/4Uw+IpVbn
UjrzMs/Yurh6JNGtDbsD4Kzpo1hpLCDZ6uEPP9dTFaoFlFmK51EEoHPJ45PZirxr
Dj62VZM3fj4KMYyEavV7wcAM/uRW1Ie9o0kh7pn9dAw7JzJOf+pCYq9OzLC7zQ8i
LSV2PuBBWgWmwyKkkkZnQBQZ3R5LjJIXngayReHWSAtK7loTOcS1bxV1qTrjRUfQ
iMOUpQM2LcCK/ypgXRfgH3P/WACowHW0xL0oNEmKMlQ5jou4kQEo/DCmyy+ct9kI
yCJH579fUDYyuFkBmOuLgFQMMvF5ePHg4+U9BI4vkgQ3Z+jPWtOAsdFdotfXi4Oj
wB8sN8wh80XmyIw6wCE92a33iaFDkA09uUsPjHI5LghGvwQtPN7gTXB1lBVa8G1r
H31/hYw0CyywBZOhmMNcCGSHg6EbVnt6m66tUS6BSh1kgJKpWR2L3+MxoVkyX9AI
lO+Lh4WzSceEuXX22qQMkrGHtdFbHF5XZlQEtozamY8gr7twCJhKZxf0sxW4Nrmz
FZBFZWei1+A5lKdsbmXQdc0AZGWwaeyh8+pDiEkL8eVKAl4/J/1Nd9yQjnJ1UoGZ
JO3SsVQabXsTACnoPLt7x3Gjhh549lvZ4AHrvdX+g/M2XLD+nen9YK+v4s7F8OFu
yhX4K+iXgk+sktciNDHLWDIyo9M2AktULGdvxVSCQaMAYWvQFvrDHKKLyt0J+Gkn
QgILoMWr0XWPa0BElNbcpWORXuhmW1mQ0DYxM1G91343sC/KhMnlJS43AwgrfZuZ
E5OTEbkb9NMpeCOSJJpcMeCS4UxlNBMhRUniwvJZ6X5Lzfo2O9Ft4CI0xT3i207c
ilK5bVYfVMB48m1pzXl9LQI1Joth/HMefgPxzkJou/5yvwNArgGhq5caV76kJSf5
RKNLyQwylHgnyoX2OfANsOmr7HTt6C6bCKnqNUYqfiaFiWScPeDmWp5Alc2b8neU
kQQpFbTAUNrIQSB3zNbFIPN5OmeVrx6kdaNQFcXi7HOmmLxDGH8WHgxfLXZV33HB
O637rLrac3RvH7Go+ojH4VlCEvXLeVnKVYLbGh3D+rV/6VCobgipLJLyivnlyGaF
iH7Jkj0JbTxNzv6mL2WZgDqccRWLXwPKvjNqEDB5NY08w2aZ3+YtAsrbD7J9BHKW
Mava7o1VGZJNNySfN+E7TlXC3jbdQBQY8HnUxzzf/cwRTMDnPoeGrvKl4PN3Bziz
9Azr9JX7DITu5y8MXA/hlBZcg9jqzBzT+QmdZWIdqnt5YRJmIFm1wMOnmAvgYeKC
RlDte9WMs+tvtLYVAX7EUMQK6mjSu+acjZZNqBzdqd151jqO0ht2SxLJtHQTmJcq
kjuXSYz1kxefCrAOhiqLljdH/tbnT6oTf/qt1JDokAbSC5fPK1g68cGaq5eXfzLC
bppCDD/Pp6x8Yvk+d+8pxkfGJpKHarMipFBGpVZJmTCB5Oe99imesIh5rlWdC5X4
Jw9+Lz48u5gqz3c+y9Ff0XuCG4OUoJHvpNDxgPqcvV4+axpd7wpJEYUhTESF8gBH
G+vPg+2lxmbe6QUoJskPbjO8H1hoGsJW6M9N1hGzIfMV8IDXR67nVKt9OMpj5As+
5ZiX2GIsk7Fg9XV/TtUohw8eF34dr0WVYtajl508G/RPfiDFWRfTNPhBEZlSjN0l
aaCiGQDxgQoWJRbqE3XRIgLT+jjMpe2k+2d/nnoWNPh2Z2mof57PG9TQZPKvT7IY
3UcDXNjy30YhPgE5XcrrAvQvBndrtJU7VCIcolOeg9D+rWYutjajwp4HsvxxyqGP
L1TljDgRtGHB61XLQiA2rqz/HKdm/nwWwqpo/ccJ3oBUIIu6uLAoyHkvDnTamZYO
p64KwzGZrxpiFNPWxxXHF/xI9aAtrrFRm3Zov+wHPKNa7+LOhBQJyLIRzbtJVUz2
+cl3t3yVU5LpwAKOMfvL8bpg0AuDRtNgmnvnIv+rv2LTU8EW/W4xTku+rj3kD85h
W7rhaz5XiswAsq3eXna/Qvaem2G8UkpZ7/5KOKFrMhLc4dJRlS5MKHmIDCIJnUsF
Tp1usKHacn77b7e8o2wVMA9QKz7s7i8YhMZ6TFr0JEZM1wGAvK2SHSVzeFqdo+BY
pliyWBOFldK029n+qByhtQbjqAb9mx0cAiF+gYO2G5+lPJcXMmnmbT/0WDU0pOll
J1BlKZy8SJMjptdwaqSgKpbY4KcIbsVLvZt3htHeYAhWeoks/jI+XLlwZdk7GpcW
KAUtbE9JmVjDD1OE52+cLaEHy0rVEohMSsVDdVgS9KNOSEhHsvrRnIHKL0tdiz1U
UlNed2T0F/y0RNHIJ/KgtsK9UWbQKbxzi+k4/p8LgUHeq92pcAwKr8V4EfJL0lBA
eGvKRYV5+aVAv+Mwn8mIMw89HRjvnCi/K51SzHqe+S4A2+2shFVtMLY7OJBGz8qC
6kundZYds2Prvhe/elsK9BjWsoxcvojXDl2HdYdjcSufu+kgk/O5+CHzJhuDwsZS
L/BEqdUTL6Hj+bCiwCGzEGEMcPfv1YuiGzpmKS5Edj1ZWqUDP/zKYxQLS1TOUjuw
w4doFdq9mzMvbZBNyzKDBkc3Cap3DJDYFYbTSY0zRaBzi14B0laDo5XKBDZOM2ZD
lk2V4xkuIPV2bwt1DYuHkxuPnWM/T5BzvuJdSi9aBVOpCk2hbhdYm+Qu+aSAhol9
oRz2W962OHzIIgpOYHaYvNiH95JNOZzDhPnau3qxnr4TFs2Ds9YdOxiUXWiCjcMu
oGGQ17hGBokXwcLeAUJOAu0vQG9nPcYMZFSc0PJVsWySe+6vNhlQAyhiBK4yGiaR
pMi4+on2C1yTmI/W8v9Ue5qkEvRKyO6tNnqtJXWCbe2m/YtaXjgkhMiIh2PC12eF
E7LZCbK18U+hFCOtt8MauUVlO5IHfFUgOCXpHQ2gUsFDRYeH3nt1zSRPjjb1eiRx
GPUyaHRjeCFQCaw4WMpdwpcFACBr6Bw/1JW/8buHgNKWOKXntIJzSWxZ+iP5TZT0
2Phn1XFzEg48/302Wuny68UYO8zITFTRNa5vYezEO4C+jDswiQUrhWyKatTXBUck
+3s9rlEcUIdUtje5ApXJDjMyn46vbDda7Go1Zdhleq0dulxmotUIp+KCioF/uki9
Z46DH9kLjs4/VIqgSC40KgZKZcWB/XObGMkJqqCZn3GxtD4e1fXr+6UjYVotcFll
o35jX8zuxRSBYFjHk6CWSqCKobixdvVaQ1lX34WZFdhdqgzlYSqfXesxND6YFOUW
rWAhKTVvjHR8o7Crj2VoosEtp3juhUUzqpRQiiB3VEyyBdVx9YQ0XkhuC3OIBtlu
DBw0HUwAyh2FFAJUA+XB7LUUvFpqKWj+PUzX2EB9sIUNfBiH9Q1gXmuyx5/sIiFN
a9t8+GAj0j9Xnc7jHwUNTWytRXenZRT4E+LsuKkdsSM222ULZ2c8wOutwu3JkzQQ
Gsxqms4Haek0bfz5G/3XTaNf+zkTcAteCBbiJ0402BxR6ONgs0Ex5H4VVzL7dtz6
pFJj0BKAb12V5Q4p9t/7gNs4PemiQ1SK9JHEZ+C6wDjeb+FlstjyM9T1p+WBq8UA
ZEgtbahSqO5mwycy7TW/JLQdfc7b7QP6Lg5027ZcrUhvhp6fEZtmkcP3BxwQm2Xf
r4q3E2SxfKVrKxwxn7oIAJcDW91eu3U+0UfKE0L+V115W1qSSfqh86rchKebN7KI
tliM53gwYZgg2IQPUtqc5T/2pvJ+UP/OslIlnBlW4U/KTm8ytcAsRbD4j0Yp9HEy
F8VWrxbTFtzuy894BijSo6sFsUorO8TwenR2v4vv+LM6zqhbWynAvl1NoqbRbukI
SksSo2xwPkStEFbW7QlQTQWK2zcjCfGmg944QlnCcMkmBu55eXliFi7pqOq4SiZ2
b8lW/Oxmvq9s7i1jkJCtZxmG2vgoQ+oOlfnNIGk128qapLcW6Nm3bI4EFbVkRBPc
aS2drbgeiX1xgoGKxlB36OIh5JbyRgxRi/iRuZTj1wI8bQMhDFk6yBq1ri5ZCuX3
g7f7kHsl8RH8Veltb46bxPsBcMfkZmdsOvOEGFnMvq5xd4V6H6kEGq/VoscYo6pB
dOUSjKsmBnHujcp5sjllaNhglmaspb6Wk5n5kJ4hZ9TfpYCzgAzbbnecwmH3zc6x
uKJI04MG80AHAeYovXSpHbtHD02EvJgTg/DlapZ7xllk1XJSqBWBlZ+vhqbKLrP7
9QAFIeE16G1ghUU0JkNH/VuId8kIK309eWN0SnVGvqFH2NNw+788rSI6OkOTty13
5x2Q6g9jrOy5Tgzb503dmU4LaXYUktlDQApzjqTzDHKSzsvIzioCcacFoIdFMXzv
q98loKtg9BXhrnEyVd3dZ0AXc7Fxt/164ivcF2gcjzhwOpoaNpvIUOD3HLOpkqNy
RwgouYEuE170v3wrwl5GyBzcbbRiOypQVAbOKHshud0JOqkAe1ouCl0jRCalln7f
Z/DkOKXI6ruI0tk32N82Ew9u+BATgstyBleRQIcK0x4gYnsx4S5S9R7yjYR5EzEr
C317beH/JxtrjUPwXLIYMz2Ey4aYNMgofgb62QnOBdiTFZkTWnEoBXlTMWpKOPKd
3QVabWE+biyYO7mHHzFfOYGizJphDc3bETHhCJzfzdzokQTclnsxZzgBXhQIKjk0
ySV6er1zr4axzSejHLA293c/5rdB9xn6DbQU68H0i1aCirZMTR3TPfRwmOIh3P2v
A16Kk+TSTO5E1TJe1cY5gAd/gMwmf7/dIPl77oFOkep3c+E6k1RyBLo6WTwO8Ptt
8XIpdaXtmZ3Hdoy986jX5w9XEERKOcRCYUq78SRyr2YuKj+70z823AtlylpfqfyU
6OLVvzpattPixnoBhcVunq9zI0afCjbpVR2HQeZkEzPKZOqiIDU4JQv9+n5yjX1Y
xK5V1HoQ63F77wR0Bi4UdXumr0Tk69XsRfIfXxW/Oj3YTktzGrkU/R3vSmqIL5bS
CjgYCCGN9ZMhU/XiNG9RAqBdFBOEAo03x4//CHU3vDs2Z+u22wPtRAwHQS2Ruws/
BcsBCVOvMvVFe8Dlb+123GXutmILsnY1j0eUpa34Sy9j2WgNDeTDlT+NryKcLA/2
q4iNm3e66AVAzHSyu3iKKzZ+ifGCUiDYqBvH/vVKxsXk35Hlr4obQ+3b+42YCNp+
CBbGt2sWrFQ7/4/n8LxrCUFsTq5gZ6VHqpY/OFeRkV6pV/tZwUwT3bGRhStnGYXQ
G66qSmMCeEnRPD0xrHUyK+ZZQpEnaxQLQI6+VhWORHkw0nv1KGcs1cXFT+4M5kao
YA/EPIws3TAc1DA++BIZxAPq2V3jrDmfJy4mpsysZIzjol80R/RqDqncFcZZn9+a
SWGl/zmOZBsmbkpXT/MS8Ir/woCPaxGYkgBvPrK2xkbbnoYKAgKqqZB1HRNoWExZ
LWNhThjgo8GiuAbfvsXfW0jRa8MWmtsEqTcXG8cbKifwUb8B/2lHw0KdtKOI5Fdo
BLbD0KWmf26qmd7Mm2Vl3Otd9As8FAqOzFaEwle9fKPZ4gtZvWU0eiEUCpqiKwwS
9VvtwdDUT3G4QufcPHTcJmCc9gJ6IOvCFFsl9ICEZJYldGnpviF66BMz34VcOM1N
Fq7mUG2gGlgk4pSdiwatIzapHfZ0pwRGKOa+BW/z9l0N/dav2YWVPn6K3uNFQDit
XWNNjEYwByota2fj7XsPHzrOPYLJZjez/vt7nt/ZO2WzZuM6WNVrTkcdyfUHO7gS
KKwtNsobkCLPpanbKKHX+28XIlKNlwCWmVYL7fF0UWzkUinrFVeLC0vXjIwI9HyX
/v2mNLFkoDuPVHnFwuuXJCuPb0w3D7MSItfuApf4TMivfPfJ2zkXnfsjfPAPxy39
hbQPjbqIhsrT7RDc/l2mwp556Y5EF46ioc32i+WiiUNTPEzqhj4Ircqs5dwUQQ1+
ZVJxVX//dV26+634Ny/dJM1tqRXEW2kqKFYJiMWJcHu6vtf4WJeVY9ldzEED5l3l
fo/XN2y5bKA+JzC9soSI5XW9CEqi3plrRl4yRzF13x6jvEa0/zKZ8LlJKM9zmiq2
s9jM+Q2S8GHpvZIKzT7ltTtWQsMHg6eerVXgXvpSWmnwy57yFv03mLbmEuwT/Qx0
ubkklzTqrRhIiyRfQY3K2d+NlFrGERdQNMGumKQ0t4r8SQnjsLu+Y/PyB6g3gfLz
WWS/Tw/vpRLT1OlNL+s29+uqX0GGwyf+k/8M0jspN+Lx7F2EiGIorbii1PbMgMh1
qKTwH7dTlOqr4qPBFKG4y9sLjH0j93pqJS2URV0xhAzwirbyCQ9k3HZo/Sk7thcw
d2qECphiVBO0OzMBc90DYoUwpnrXQWH4NWBDKgFOR1IWoOdzH3Yx8VdeTwr2vkJr
NyiPtv6U0grz9oLQSfrqBJibUxWxR43LU2MyUrHIK/b+9qKQsJyujqJ12EzWYVdH
OSXZQ2j9RDSajoj6ivHbE+aVUXXPELBebys9UGJKhPID71sqN8BRjWjp4mze1x1U
ZG84JUr4sgXZnyA4QIz/MkDIAgxTwLXsaZM+uRZ3KAKewPnsVYhHpd6W6YeRbdIW
ALvQxFEQXVuBA4YkCQ28lvlm1YIt41/66WFZvxuV7lYBW3MnqHe4yj6oND2G2QQ1
+L7ijgDMuU8Zgt2ml5owZD+zMbSL2jHNPZfie7l71UzNDjaFnDQU/zkqrkWLMFTu
GVosR+zw9tAyiz5oeRBsIYZKlxxTV83W/g/P4q2OaIAy6FhOoHf6mOnFDcDCT+su
2JMa2ftLTYQZ3VFdd0KnX+TR86jjgY7rKhjq+xMvQS7z4yPhGIvY0wKRG5Mdupkx
mo74XOOXQS0aJlkb6WK40c90CI2RsK9gPNBeHhj7AlkomDoBkFzc3aiGSj2gnOMe
fKZdUpnhZo4w+vlDZcKPx1FxLaByiiqRBEK1esFjdOSamLtPNJ5WusRbDuot/CjE
K31SzwULeca020cfuWSxLuIguNfAAWf9xFy6dxgFoAbybJv8QOtGWO0FW+bX7H/m
UkwMslYEF/IAZqlarn9DN/1rcqcM/H0QqEWtKWLewJ6KvtobAmHa2KA7l/C90A+f
RN+nPcBfrugU6hgxYyRXSuhyv+NhHznfVPd+HUDRi2szzSc7vlu+mlYnQvAE8rgB
UsQraGqp2QMbeswLogmp/NLKmgk83yJ4gvDCGMsocgD067uHXx2SEhAoEhH3wAji
B7717yhvEdQ/Z+V8eHsFNiyfyCtR5PlLxqx/8bjb8iDBMTKkniQ4UaNskVZ+SlYq
eNC74kjmDRkHVQbLj5eCYC+0MgNonvyRpnId9zd4+PoleS3yiMRPwOVMy6Fm9NSn
CO0mjgby0TZEWKX3zkdzYZGZuuvKjjmKB+jA0mr4nh7jaQbyk7sq4qcG3VbPR+P4
zeSKKlcsZJ682PEdFOEYiz9ckP6VNky4GlyeHU4mjPW6USVVl1amfRoU9+7/Iblj
ctAfJEKVp1lQTAcFlyp8olncDRK50mvisQETqEqpDyDoUV4jP3Q/k5KMO4+ZIIgL
Cu55RgVJhlbqcLnXSrizeeyT4WP+RaLpO7b2Ba+tnX2sChmZVDfzS6NzEnSyCq8Z
0GsBXRnBbk+S90ZvNGqEVEWFgUPL+pjIbZ+qhdywBV+7oqlMPIzrTx6wn9qef3JH
UQ70FJ6GWzDe+CXgtNYaef/XCn5IH4B42XuwgzP57u2/jwmPicIhWKAVINST7Kgy
JaGyc+ukMmG3hhZPjBC/Aw+8KNNMr1xAaIng6g4auW6ZhncjQvWE97x3MzT5URrO
4MLRAsbYSD8RaTBnulgzQ2QbFDCCDjN6uffL0IImctwweoCPy4j3+6IV2Px5MptE
LjIyJQzdYMUnX5b+HYo3PxeOaY9BMoa0hWSKeYUMKlJm+yj2Kp3Q1yxSyS89ZHQL
WCP5j+zkkEzLkKVUl+4580pcXFMEFzb7SE+KIPklTiR/ZTc/l1yFPBLPT9+mAM/d
pwkbNbalDu8oiWWn2dOtJgSmw6yzqRByhB5/V2kIbUF3f94dFKUdrDuLGlN7ZLEs
ULv8FfrI5Pk2edR7leWAJlIZBqz9I6IM88mzIQi9xrkPuT2JFoamHhNKh6aWttCn
n/7xpDoMR4B7FbNfWDG+Hagw21YxcpGHLgBsJshWftMWRYA9eDTGOLPKpCcNzYXL
izcROZvHC19kupJdb9fXA0xjr2McMdlIq1oCe7cJv/C8i8azTQpIiifGR/ZPTdQx
cCIaG5mmqQkZ5B4Gqo3lIhrh7TS08dYV/CwNq34e5zQsc5b/ujhtImhD8R6zFk9p
nFKL7ShJP0uJVsO2h5oqHmVEay9YlWiMttSGMs3wjT6M7hGwXYmXZCjMC10dhtOq
G84ZVVtMSOtebmmXPn48xAkP9+2TEXH8Udza1E1KClhMLNSOFRYIfEtbD9GsyRpK
unz2PQri0ebmcBDZa4fZ8BlI5sSdpNNtKK4pa7RG7Nry5owbXV1JLUlLpVdwaL5H
uoeN3RD97vr1o0AQnJl4mJ/aeErztvb1FA3orKrDFR8yyvIhG7T2IG6dKQmMEO9R
vBQkcbgheoHhKYaw80nWi4TDOEeEfth4E/oZ+cZSBsZOGk4WEp5PKp9lbNtMIaCz
A8Mc/pQF4PO54AR5Ka6QBMlLjBS+mv62xZsQo+xBI6tYmPmx3TN5ZauG2Wxvqemc
fcxx+f51MRZ2AvBR8PLuICG9Un8PxR5gOyUMVDwMepIOQC1jdmT9W4R8cL7IIneZ
oKcDafvJETw9NoR8D/1HUfA7IYflAnvPyo2xLnYnCk1JUNtAVkrlk5Q686q+z6uj
CXVLkTQtu9CQPHUnVBLYVAtG7UA15Uz1ztWC4lvwwmm/uKgalLiW0+7I+QBbahIX
Mb7gBJ+Qqw53d6c20QxuNWmDXSXYp+L8J+IiCR1K1NjAr5ahuJhvwz2t5H6YcIEA
oC1wRzUrScVKsxVNzdRCYz3nWz59EFkXSvAHB6BRtHj5Z640LlnSdY0jItJVjpZ2
ybo6dUCpaIqPSzATWGBI4moUWa3QJ42Tu1JKjKxy66CfoUR84Qn8pMTKIOU30vyq
Fcrwtjw9vhhTHNIvnNVDvDuro4Vz1yVjKIqKTzf58ljUW5+8yFUYN5OM77zGoPYa
pP+V83aeDODntXvtWx4O7C8zGfypIM//MWFWzbSK+MocEfGkYs5BvMorpI54ST8a
SzMstg387j5gM+PNXzQkMIS3MgHW6u6Lq8Gh8VO/DWeysWBKQFVTIJ69hLzkh/Bp
clbelrO1Ft+E8Gnf6Q0PvpPcaQnIajC8yrCOK4BErLaINAD5UTPk1gKXTX9mNq4P
zjHxiGUuNfroYjwnnwVZNQ4nqQFDUeNvz+aJ9cGQ8Bw/46Nd46ZSKUlzOMzbStc2
FWguNAzaL3xbBnQt0lwtDtFBNYoAfM2Eog71x7IPPHyXCTRUvFcDESDV5lxXQEuR
4/arpYQ2zsizZSlWaupQhszBbYb8quU5A6AdkZsWCIj42S2jFLkgJPg70WRafMT7
z8PEiasGDHJROpYdL/GvCkVJktv4j83f46ML5YopdExUZE1BlpqrZAY5SzT8LsoF
NtWl4OQybH8bAPPcfYaxEESOvDNfMi3yQCEh5i1mwjPSrHplxiHsgoL6FAe5DkHI
JPTuzCpBT7i/y57TJ2rR6idT3+lKXcp8MeIw2RdL5n5DeQH7E9QA1XindTOUYhCH
tOugHX+YyB7iT7G6Ily/fGEk0uNKtzVZaAqNFVGrYr4nfAIv+f4RPIOY6nDPxQrN
rzcMgIkMR3eFxRD6+9J1M8lN7l1+DKm6cOPki2Phpo4/aqLC0ATl+wlPljBNrudA
x+w1vNBU7blORexRPHdqxE5Rv4afBoO9vVaRTiydaozM35vs+UqjuZlkoc6quT+O
K1hHcknRJDlxCJbqIEW2wqBNgGwX+Ehka4MkYHwif9SdLqmCZjS5kY1mgVp+/TJ6
tX+LJGlLzAdfFl9AR4b3JOm+6txbIk9zigPSygYnsGIJNSDgxaGrB2vkXyPQOdsS
AU0lmbJelFttON5G2PTIcMMiKY99MfmaIOcNMKR5T/3Qo+MFjuUOiDik6u5gWbr1
qTa5aMsEjCMEoCbkUZG1VooZRP7ArpOtn0sG4H9vSmMWx8wQ8soj+eogpc0WSDbz
b1OeyvFHhVnVbp8zYGE27LgnN9pBulxbN1JJ/s36b4RU7d4OPt+qetVBVVBuEQ+I
CWMDxejzt2P2atDMygji9wicYHz6wGlZRppuPbZs15Ep8FRLtN7V1OzWPBONY0s5
3Oo2dlOZ4qUJjSEJf9YF0wsD2AjHupx7d3XTAJoOUPkPBsFzsJ2NmTLASZSelfJ6
fOIqsf+Swz2QP6ldKmAh3WbwbMuPFicxAos5om2+kAZCwCnjlzS30o32PmsdSLNT
RWW00qURShyh6uFp58tX4K00pG/4bZHeVyKwA+tnnfRXBv9BJRjozgCz56XKZ7g1
xBE3di3HzgqUc3N/8+pKEGOGM8JZj3DOhkvNZtec8tJ3zyvLXGFI8NwcJs8EP0wb
WvsEYc2T20biI6NkHfXSb04IZFW9e/su/xDlUAgSMZdaYWOvLQ9ljg/tpoHjnfU2
KeCy5CsWz4cthDmnekpJQqTXzNIu1jKoQjNFRdSeC39h6fgayq2MPct0sxYr8vui
ImLt5XNlerzY+Mjcb6xR1PF3bNdWDtrn3Qv45Fv/ML15mAUHzg+p3YKPgoIryT0X
gTFbvC3R+F9luDHiut6y4HpnoQPv6xsnRjQZ72nptAYWKzigmHp4EeXpbWRLavRQ
uA2istILf1dmR8mqKSl3cd+GbwWs5pO/4PCVPgJfTqGOQ3oeRDSr3pjNCRI2MXlB
Gcm8F1TnTtc1jRbW7rDXUlquLtsrEWuzxt4Wk2B+yI5MdS/bC0OJlK1mp0/DGt7u
Vszoenjl3E1aCCheeRly/3UvpmPhCJBwMojJOeFe+znrNNA2OykzBy94H9uoI+nj
WqC1A6r0Hrcrx6GaczHiyik+jKxieo9gGb+f+wEfWiZs+bbeue1IRUMpZToEL1FZ
/8ftK+gWV66L8+XR84o1b6CvSnS6u8t23Zjo6kw34z9K4Nus1YCnEuStk9e384aL
Ot99/lEN+fulXHPC3eT0tJE8PVvLBG0cbNNZKRsc1KAySwx5dDKAJoNP2DCj01SY
n4Ng3rDB84Z5hfKkXmT669bse6d8VxP9eQFoX4Fg+QJuNhH6gjPyv2YPtICaNylY
kZU3T6mX/R6AnNJ9tshEZKTndejw2JHqUuRMODJWBaYR0cwPXkY7zr236v8SqGy+
VKEtvCNOcb9mujtqi98xJ+getQ1JWCpA3QNcKfzRNfsrHajjeRLloPonXBZFq+Mx
2bU4PST7jYN5I3Ml+PXWK0Uxn3rby5tZJ1dHHSX6NArGp0wAu496iE4vLIFfaQap
oomlFklVNWGtrTCtoM7nH7ZExOpDzboIBS7oq7RnsDOitdaoBVWNhALcXKulk/F8
ft+Z3GyFBOhncBhH87Ky6xtvaZr7MpK6XEUDZ6rGiRdLGx56Y1GZRZ8S62HP8NVb
7W3zVRad3chl2Sm00dLqlupSQRepsNuoyACsoGQjQcjFkTl7wI/QG9wXyV/ex/mI
ChP+V6omOyMXm1Iu/D+qf8cNlitz8imNG0WopEw/qdBFPaSfbv2j79X2TBrjD0QU
RcEtdRZoe00k00xPirswS/8rnUdwPVL5UfS5nkpHqC3GNy0Dv6Z3vwPEdHfEWBsd
J2kYcvyAnCOWImpQfWqUuwp4ZD03xPyA90QvIF4PBDJcc62Lxf2yV37RA3LA6Riq
I4t3Duz0/vvs26aBQ+prVDK0+XTgIXMCawQCWYpm5ytXUnvJccJImbPGsuOmGlOm
iCbyTc2sMOOPDDmuqgMYzyEfhTTj9kwABvusTPcatsKRI65HLQJN+hz+9EYvHEQ2
KsL98uNNHAVKRJg3Ez9cxcZ6JmZwHACDWyNV/NDEe5A9E5GF4tSZuOI8FoyjHyST
iQped8S+HInAb/VUYeGASsiCdc9G1Iqu3N0DtcThzY4CroJ4JZda2A20RNVkA+lu
czq2K8e0KvILgNG2UG5KPfH6LktQI5uK2rpZwbre0AQ6wZO8BdGc9zBebpfYTni3
2C2fExKgOAQDhnr/FndsYuphr/dGwmHn56tKlPOKlFsy8KhwDSvkLxr9cAFAlTHW
sHkN0Bra9rXhPyV1cGwk6ZWMShkVccxbl1GTL+KPZp2v6XIpOeElbQjAjh6CHIAR
cnt9H23dcvvj9ronxA3r94FeukVZgpYD+EGbcuGnAzJrOhC+HWeNNtjiqkjPO0fA
lKfxqxDS4AsLf6s8D2csG7sfg6VPQc6BMSkqvguIQyf8dbio0KXEczzb8J9a/JEV
Hn/tdAFRre+OGGkA7eL6eiDBT9AqnuY7y5gBPJZoYKZbeaDopiExjeudFYyFTKeP
O+9hXECf+kMGs/PL0bsHYVP4+rXoNH09/q3LaTJm2XJ74G4GZ7wfeTFMw+I1yS+i
Fem/MSHHm4yA8ndhWQNBWkwDlU3CKGm8t/x76tmWSbZxp1G/ATdHvcBveo9ONS/j
JbRXYK9LNq1exXq1EMS44c7oNkEb5hTVV/3TLP6BRjqTRbq0QwIY0OhVCncaClF+
n9tJwXFXcl/BggyNj0AKdX/IRrR46GCa8n0gVjXvlUq9OH6YgPwWlQs9h0+AbWXx
ttnBnTy081WTh3gxWJYcblgniDRZPXq+iuvTbrXrjTFk+QvtIze2Jd6b9Ehms9kz
CezVjXVBNpODHy2MlTnKEnLfGUxhOhQwcbbjucHtz/vWi94XS4WAXHCNWSXVrMhU
NElH9XFkff6tQ+j9dMqT9eBu171UfLwVI1R5raFXiWs3QWqUPTwbzZH+0BRfo6tz
hAa4N70CfgDuYldkbQdztvfh1c/nLFuBj+Q0GMGZfY1gcQeDz8h96nRkqG6pKosJ
+WR6pX2ciALdO88yK5pFWYsJCtPw1YM7mHu8jbHGbkOvNNmMVUi38avaki1vhe2X
0CxvAxR6I7toUffE0xa5tYFW3zX32igI8Gc75mqakK7o/sPKKjLUVsix8uIeOezP
GMQqqNr85PdA89/1NIbc/n5A55U20WtvG2kEKtRqmMGXiC8nCJzR5dcMjpAzr4yI
G99CxS+kDtVnWr1DlpUryjjfgn2G9MqW/SngPrrO+udIVb9NpqwIppJ+a0cOLZqd
IwusnnZsSN0WXe6YjI5qXSpAGSnz1X/OBeFrfRR0UNhXE/LYiOnjMgkvskx/NH1s
x30f6uQiDpZ0f+aWCnDebefC6Rtg4cvApcASjtNzobqeWWSoqQsNtkK9eW5Gg8u5
mqShjsbvXn9wzOTBLIja209/wlxY26Kpl95zbdZuXt2Zz+hamBcu7f+Wrgca+8UJ
rorOHNoNfFARsYJW6SjGn0h6LF7jaX3ltF+Jy9ovLRElqJ8/1v9QhhCtztjIwpcd
M8Gq/xcGFiubL9PZ3+ZLSsZw/VLWWwOy0y+sSbqtuDu/fy/ssmYmjfo8hnuhbngL
bcwOBPIcAMe23LQaSmHh/u2SDf6h+RBcgCUJZ+5Ad8+Y4PsPiYZQXb9NlYT7NyiB
gqwWbelUk0Q09ISunlsfNxpIICh4iHmwnAysClD3zjhQzQ6C3H9WBDS2FPre8cqA
wnokRaiiWL0A7ldXkGc1JL4iG6k0cbe4iSN30wwM33cuRNppe9L/av5luhmfZA9g
CK1MGVMbd8p8D67PRDKPPXuhuzhbQo5N+pf56F3wGwUBsInDM0RO3cqSm+JRHw6F
bg9DR9YLbvU1hGwezp0d5xmgP4AwRaTxwzNnjp7yK/QEMIKtTavYXcv/BC3/Uxov
joOn8tb7zgLpYEKwsPdYvlfhN8pvt2P1WjL+taAKn1b8V2ZobCIDQk5Ffz72DcVO
nDvcB/T9ZTUN1qt0Ga3nd20JZ1dbMW1BSfo7Vwe88OuwL5WqL1/QmT9neq79qqQe
tkkJPWny3zqeMdByd403MbvAV95imhAdnUl/ooIFPbkFXYSanaLl+olECGbiOij1
6JPRYtOAEqaaoug2WuOJ4dcLpT7nQDIN1uXorbZ2CEMCY7+Ck4wNQEsBGrF534ug
a1tMcyMDqln55ay6+sJPzG03xsfm/BZ8DxewfGKhYt2tBTPFXN4fFAX1zbTNbKkh
HeTgWsriCGSKMs421tIncgzaXwT37BNbkD1BxfC0odRdDEthHAcm6FBEGDMv/rB1
t/PyPxJUOE3ByIIMFcuHtIkDtTP7inZ7Nt+vfHt4tECQAaRXf46op53KkMtI5jHg
JNbGFOcJD0u6Re9FSu0+aRPyqemf39ABPcQbYhu5df0gFdsEu/ZMBgxhAIA9kz8P
45d8+LKeDwcHUHZmkUVKBZfMfT3mLCu8CuhfKCvqbIB+R/lfMEL9Sx/zoYm5yj+y
YRaar3jBKqS+hatTlqU8OKUJ8rnmMubJhX1PoasW80fPz3pRPRHNO7to0TZGl11M
P2MbM90eLSTDYwZ7WT/LjZMXesmOCKOJNHh3VMtQeyevSOQVfS/NZ4LhArwqknua
R03mzJWcyCPt4ixan+FHQVoDfzcBnls04FWpgCHqNBuVSfP/jcmjPH2KafQ/HZG4
A2gtwp8sL/7Y6GHwJeSMgEJYoTxktFM0/CRhNhCegHxS0tJDoMnubxXEvYnov9w8
uqsJZ0qh6nAi0REK+BuvkJPJH1BLD9lO6CfvwXCObCTnmXFgqwIy+e2odj9ZwUD8
Xk4gKuy5vbqFMQJSAVuW0fNItkJ/lmTzb/1E81/aechmHAuXtodfxWWCgQbTpgPf
kmnK3rfFb8a68qQC97RkbqnCUMedm85GQBQlKz6/0zuBKrVbq9FU2qt0FK8FH0yU
d579W7t024M+epdA74W3JoPPsHpiHGlqw0KLouCHTAsCrmG/rbxQ/fhIuBrPw05D
sFPCBMe5fNE1SFaNM+l9d5lrSJ2zoCpNIrpEX+QwYL84mlmgMiGb5ffGdttxU7Yh
rCx4jWj0u2Q+u188sl1Ezd5D9nBFIPSHIBdgZXsY80o83EmRBHRtptFQOkKn2jsK
inGFKpmBCzIpdiU9E3C7dSOIIV+1dgK4vRbR0j/GvGt/NZbPq2M9sDTmfKtanG5X
lJMlfr7ZE7wOrTRpwndU0FJygmGP2hZvhoPsGgf2yhTMsykcVIrnakSamWY3R/AJ
X5S0jNAg5PgXQCfhLBgrM+cHmqTLFVkMXQwX2dHSIKXSGhZrXzUHYTTymOOQZJlM
E2n3jDW7WzyOlNegUryYgLSPZD9Kf6ijZzM6m00kBeThjZQwqTYwO5MOmW5f3hT0
olcq3awiwhWeFulRL/bBrLvfkTWViAt14kFKaAYKGTK83Nel4RDDL66suIFskMPY
qK/tHZcHcXJCfLVOPynNewS3YhKiWhT0dFzsMCWtZTmWMMiW7Lb1pstfvIOi4vSF
cQUjrMNoHHMDB9cpA7MSzyC5+0KT4KXTpuSfuNJBlqsadxqv1AHfdz6QqYcGcWfM
MmknLPsbZJe0bPpRxlSo5kFnIFTxSyXaO4Gi5AofuNLz39LMk/fP8JaGUtol5ZEm
aJy4Xc7LA6OGltxAqjvCKN++Oq6EMTEYuU2+XWypbXsU/e+Oxkcztd2Q0qwN4fVR
wemLhs7Y94HU2CLlZe13ZXvGpFAp0aEFNDYJXmjioMbEPH7p2fRYuFX5uWP3nE56
uykwxj62ceic95gUTaCJBxHjgbEYTuobkvjAe+EJEUiWXASWcZ56fcO3FYolzGUt
HHdgV4LLrilUSkVSWMCGZwqmqCtUrwf5DvMlNjal09ATbx1xKc+0eoBiLqZnkNW8
tS9i9aR71eRo8fS7dyJirnmtpGrk9Dd4tkSTKMBNkDTUPHHOGi2fIGnLuKUCBJF3
PKbQeoBadb+x8Km7utsY4qgyurzJCrck78fRf0QTWhxZOoRtQ4cao7QZfRAsdq4R
5kA/q+tzP4a+nVwYoZPr/iWVcbOzwCcF80IUFeITu4pobnkv/oQQpw0hbj1dzcdx
E1411scksN9lMgypiQU4/8tahotVu+VGCZpmaC3EuJbKF1HB6NdXO3FL8TjrAwUp
zcxr0fA7P1ztzyC1T5jwc22K3/9ic0S0zdoNLVvV/CaN5NGGBKX6RdlebTY4Ond3
XjO6KkHJHjhaW8ff90OGJi+LUAXoWa+Q+eKPr5Bqo3xFhG3ppiNeJgzAx3N28Gz0
VRU+jjpqw98wbSGOnA/uRjz1x9CmPFxNMRNtFrsn151A+iNrmS+jmIYKlj+Z8J83
VHT0TZOLNz+gIH/zf4W0wHvo3cWelJeN3iHVIswTGDx433RuPCYtMOFgIezHNBy6
NaDz1aeU/hjEfJDOw5XP9AmMRV8Exx13hBGSoc4krj2XOTNu14liGA+PsW3exfJK
UD1Rsm89x5hnH++gWlykIFO0nsOVW//7klgFdstjD5ZQKtLOe9uM4qOxSOiOGTL8
LjK8+DFRxfIbbWloKKaM9EQjZpKHjb1KEmaWhGGV4dIFUQ3/a5eGg1d/2pT8cZ5P
djJ1USalEmNMHR/m3xpY17WYCGwrJuNmmgZ52sXiQPOC/RruWnKVlw/mBD6KtMdv
o2aoV6sLIOnu8dwLpFj0QyVSFWZB+mamab3HA064NA+2uI/cGXOWiy9sWk8TnNOr
pzA7eaxW/UEEaV3+MjwQfDLP3VqZ0BtRM8u5gtfTfAY9B3Hw+oLo/yeXTCglnsCE
bcGYnNgWwDVUNxqXAa3YemrB96X+F1l3d4I4J4iMCtEcbFCOAG9hfrSrWQRpUhni
IHGr4EQUG999QlYhwAy2POpW3XwA205xV60BQvZwE3daATYhFqKYeYHKe99CryUL
eurxSOwDFXZWDLM0Y3J9sGbrRe7eygd8iALP/5tAREMeNjwlHXOr4JpZ7l7PdDYZ
INvzuFHgqa+xT4D03am1TiyTAsRA+xyoNQL/vBfde2ibnNNLoBRFrQ2jGpl6DgHn
3gtkIY6zToOyKpFZDdMz5nVCedXySmYR41tdJg88QRp+v6ODAJib9p4pD55uAdLw
Vck7y0HTvTFtcTPZ/aSYPYHxlnGZUBUI1qukVGKC6thSLx5Rui9U9yIxskrUkGir
6DK1OYlh1HzXpDMPxSB7NCv9xmcL0wv0GtY6oe4+5ThYaxf2bEVu0X1/rcSJFIvY
x5mxew6nNCRNfqG+MggpqhzwS8+5BaiTeXqoLjMs2A4DZD+FWsqzTd2T8Btd5y+A
Fu3Gi2zdUNmj53ehBrr5FFr0nSEvTgMuBBiEYuRF+J14nVl7k5Q5/P5U38q88RL7
p8U8r+jgc3ZRLTuTUDPmOMwNL6VSLh0IRp3eqhUDfzr95cNZoJKvGTctGEfgUrBg
kWJ2Cf9bN/wUuDFTUuXWIdptWQfsvu+mWSTI9ugc92Ch1LzH1+ABmlEtbTgFG/vX
f3Sr0gNSnlhZrEVwin+0MBVcbcTfzUPa7TOyHmhyJ/na1C6NnfkM3sU+Brp5Qq9z
J8YpB2kn7CbGR2qTwL6o2cmafev2YZjIONFS4UCuLL2/X4UAccOEhB4tCRLRQJyc
KS1hWcjEwVcDPQwjLUcUxeOl7jDFFWLGFxzYijhNhPPUhmL2HBP/tVz0HDAEWl/m
j48ZcyfQKdLH0RtKoGVMtkZWKPo60ARxdTtkvDH7QDHEJ10KLdQ94lSmgpom1NHB
N76n2WMm7bcHgbRVSzjraQQ/WGoX78YCUK4IkVR1bNpi+KEhfbgfuA/XAgJMCVQr
2dePGfHo2sqambmICWAF+sJJXg4+h2rKLNYLSd8d+VvNyExisUsviA5CWEM5y8kE
UlZ8gKpe+8Qdewd9l2OrQqLJm0tr56aNcofJCS8/+ednGrXXnlzaXHXeWt/mWItk
X3YRKl6zH2w0AAnZjbVh2berFruAzPrbtcO0HH3CcdoyipNkKsOBq+fs8IUQ4KzG
RsRdMhNFgswZlrowD/XYSqIlOVjrBXm2spEMeYkAHninTenrp91dweFApOiIfPsH
VeYJ1UMaDPK7u0AATsdgzcY1TQN4oUAXc8n35d9x1iwK8FeiNEIDjuq6iILrxkPy
pD+6tpWUjYuD8syZhW/irz8/OSCeCoB14HWZveApR6P3tG32LhuLB0UmlcE6fK3x
4qHqfSxa5YTzENTOcLMhNp/IerDeO3CluDSb+bLIzS0Wv869MP3GyjyNlv/ZYLPC
omp8ubaVLaxvn22B5kIBiItkvDEyngsjPrASJO3FGrCJkzGcqJiajBR8ZejqAuRX
LI1QmvTVa2KmOvln3A9wlEqQ27lvT0mPqjtQoW886UomJ+TeQCCVcXpU7Uja91PC
sjcajyC/kVuMXDpWOxP6P8b5mmuXMzoZeXR2DrGBwnmnYoNa+uBzMsbuC7td/fva
J56wQ81Uo56uDOomJlKoYreOsEPz5kt/uYIdA5pyT1oyeqihPhVFfvYPQ/+8L/ad
gQ5TJD+He56D6EGbITi3t/8FEm7BtBfcgnbS+Eu1Oo8YKMDQf2KNHtF1WLLhOCt9
6BkNwfz0UBEzqyzLk/eEPDuzkW5vruWUMzmpVZerp6EdofOXNtWEp5YtnHWK5hNh
82w+nrmqxtgBK/QHBtrXvDqdleFJWFfgmQhxHF4Jet475cY3oYaINcjYheYjjCpN
nyva31dAveF83/wdQPMR/mkJq7S69cj1ECsKaD5kCd3TtfzlM2GX4+N9l/Q/9ZPP
dFQLVSgWhn/MpoX5CEYNUf/1guoDHQK9H99NDhpq8VdBXjmDrDiPZuNhBOr34Bid
A9YbBTh6KUYKSQZsrvve1TWAVjp2OldZMuNPG8LWMLSlOvU0r5eCP2uoZMDlhzQx
6mhko1iLT5MQR7JOnRDr1+0Vl8cqfnc8KeW0BLE+1ihsj1idbmXOcV1/Zph5kXDZ
t1H0wnEEQjjoNkSIZgw//gkgM4M2+bopq3RGmPmn59rUUaeOUS2f1XwsB79YKEXf
nkLL9AHRH5zUeAMqR8WBiIuXWg7jXSk+v3QeX2D7S/SN4zAi9Qtup7gjkk3nLGzB
yMkcgg1gqhpRyhdVi9ImCjav65CRX/I95O91a2ARmaaEtDmnw7RFp1cxzoe0l/9Z
wEJuORmu1j2KkBazYuJ5As79adIxl2RubP+xT5goSC61R3P5zZonm4p/zn0I+Q6f
N2QOJ5pSjzsxlXvYGOjPSwgfm4iaWRbqvyCLtn6U9GfcPVbCMGTEEqTnKj+84IXj
zCK4a9A6yr09eLl9Ntpxxe/ierTTlSKfPtNWIpQdz8eoN9APnKiuMJebwNrEFyOG
cpKo9ApEJzT1LFw6FXpEjpHtLk6bo2l61+p+GQ0iXQl8suUTni1yRp4jEoMYMSJg
KGeh1oRe1nSwFKiWxSkgo5f21hiAVU0uRRscEVtX7RVoZRJdJSlXKw7viH7rzdN2
KoHxuxEAA3qeqxSPliwsuKEaWxhWXeTEZPcV+HR5g/sq26mMwtXLOI7mWZ2TDCpg
qau1kMLJyhGs7i9TeN4UGq5h8lOg7WsrQmuAJHmRvEwVQ1ehWuoZqonnyVfmqlIK
/13xcIoiWaNYbtMSWipQkEg5Au/DDFXx/ClAjrP44KKeJLxuC6Oai87hV77RxfrQ
DWXIyTWRHQ3CXqADkMMHMPDX6iWL/ICKuw12AVSH/QQ21aPQPBLYMJ7To38AXtWw
zB/c+Sqs8H10PYJ13+RDxU8jsgA03Du3YUuFVZR0D78lKipg0ANhj24VXbmRpyFr
XfxjqKVtbPNPJKvececVvOQ7JYtQXo6foxFVHPatR7cJIe9NxxsIqxqxZCK2qQKG
48X09cNhQqDWatWmDQ1hS704aV4o6avpcnntiW0xymOx5cS6pQP2myPKq0F1Bvto
uTN9wJpxvanWZ+zLgh0rtl6luDj6J7EB6G+gONANZEI2tfdOdkgSvi/9e/ZZuul0
LDOv7oU95zr+HEaYIiBR5gX2K5qnL5a5fsg77j5Y1ztW7BymkXGCk9S+HK7bxsxN
npUGmBKhyUjQx64g5Htnxg/QGDcxSrAO6uOQc77asn2+SDN8AZnTUVKCxzk9ZHxY
Vm4bCTVe//zIzrcBgebhG522eP0uw58WKCb8aJ53XGHNDEReNAEPzktICZ0oKvFj
DvQvbWbQDqbApasWFq9r2etGmg3zOk3d6FGsQ1o+Ei5BN1enqqfMXmjOMHFyk1FR
ngHDnyRLex5piNu3ZFjfDjb+6AJ17uRMWU0zKAn/kOPY0jFJv8UzXTn2eIambzqt
bik6mODazqDglGkNsvMqHt2s1YXzg705klVReKCbuCPgB3LQPGZy8LmHym8COAQV
iscd/EB8c6xLHZi7TKNLhWTW6GWsjCb+NWN+POqo7BJCixFFeyay8tLV21t0rNHl
SMEJ16XHbBmrDCfENcBuu5HcpfZYvn2H4D63YgmUbuhbwjdeFmzN0FCBh8rEZto5
cB7FT5pEA+JfSGWOc9IvjoJnshz44n7YC2UdwfEGMZZjHU1e0buaebb7xLXKB3Y3
MdmPGduvReAaTfqHQc5c4Y4YIum2MTi6cgVABLd0JtaFbu39Sdwb3YUv2zoNvrD8
R1/zQih6A54gKf5/wy4QX3xobnYZ6EG8XRdyp3fDIzQUoBsOTEiqIn4XXjno9slq
MpOcmTENVEaXEodRlTlpg4pfbTIj+aPtAv66YQ98p2j9fo5jCkhrboABgXg7U15s
TAkhhQcFXAFjuu5o5w4fzYDvvReimfhjqU7o34CzR46flCFukmmOFbVqV9HwgxpZ
ICbA6QoQ7caDLqqLDRuV+njXnVB4YhCOw8K32OxzKHWQJnYY8AXmORhK7Oyzbd3f
dRwyFr7FW+iX9mfZW1/e/lOg6JgqG9BdXWKFGfjJRsVZG8MSfmD9MlF5VOucm92g
/zlMAUkaCV0wntsQAYm/TJsa7e/FxlbiAQqSyrL1lvU/21Nk0vEazSAc25A1yyTQ
Z+GSx/VnD71MSevYgWl2ZlqgnTSKRpqvI7VWJk7YosxSEvcy0qmjNhGq08YXZT/w
t449lDmyL4Kb6zqVQNS+B4lAGdXLWEOjLBF4u+NfB6SoZjHQ3FwDYvZoBVeYgqiS
Js2tOaePQkoE7Li/hOVgbqjRZaN5SsPVrQhn6WjUr9F9IClyWBgswDyqtT8Wu4kJ
y1lfB2D7dgGcCMpgDdtxTEdz27dYf6/cCu7UbXRFFCXZ87LX1vwAmfi/zc1gKVtL
Jpa2YqYLE8KRDn/nqXyt6+qvUYgfXnzwm8HnIMZLtCpTXTK7qj+nmSFqxIv2CnoZ
UHxXJ8LxWGRIVitjBRfmBe6gugFQngTxrFhmsr7sRj4D6r6V5APUro2syRf2DIEA
yEoiCnNEgR3utxh7jyv59LUD5ObH04DJ/MLAwkXdAuJIuc8K3AEzbngz0lZtZyzT
83CniFKNXscN+jIJ+Ko5UOM4ZNDsekPQGlrNf9bnMzu5LXSlcLC4fpem6lcVUASJ
aA1owqpTuWWHdVPcMIUT5zZPw/LUvhEoIW7wSLtao80tDlqWyIitG74KFUqlW1yG
LfQqBUyx3GYWxK5R00zM1vno2mHjrS1EekOP+dJA+rmFI4Vkf/cfo32UxrnMVf8i
2ru9eGLaII+7QM+2VuZ1XVHwLVHAM86g/gnLnXrbuxCtnNz2w13u54E91RvA3GxY
z0T4KfTn5cPuOu+TLgF+2ShRIRlu3I9H8QgLCzAThz6SuuyxURBE8lLA7DhujVEc
reKbgETomEdqKnKUFt5zsFpVi1uZdHeAWuFeOAWsVMj7Uk7N7JxKErq4FkB8VOxD
E68F599z0ZDikcn7sF9rHWwqaRS5MhpoqPAx07fp2dXdhgtEG7RigOq1CyLwjKDM
goDktOlQzcP0yCz6KfOgx9/ZCXX2NY45hdiKOgOlNDLAyWK2nh7N1P5vXh8VBeIU
JY7VoNYsbw2CrUAT75uV0JV9iT9fUos/XChM2ZlGEIsFJopqfeZd4W3PVPPX33Cl
p4abEhJZwgCwhbyOp5nwhKi8LJ9NjWUksL6a8gLS1WNszo7sI0FaUjHtVk3UulHq
0fKpUaJCCUIoYmgPKOzCY0hPVP7+bOjqlgv/N8SnfcuIG4NA7ooiWt9aQDoib5li
f+3+t4MVdqXevWRAZR6CSbwc49edn1inhdXRThNDz3PwGK3xMgCmzszV+uZWyurN
drQPGTbc026KMz4b+nmaghlDKuqibvjG2QjIuaHBIDEWIBvaNqJrh738oL6+nC6/
ydJep3ASgs5coNeod+bNpotYtTfX13ypCcyTYaE/7/jfoMoempkRRGhT/ZSTxcay
eyTTlqgQp4dGdV9bmKg7/qi10gi8cqIR3jpvJxWdwnkCMxssw1QUz2fsOekvAtx/
kY6nG0+/WtnrHDu8/SUusXFDWmi29tJ/zmIqyLedzanx0UR0M12PiHd44zugj9wS
qcmm+mad9XtEY5Vjr2PLg1AQ0+v3tKk8SyvE4hn5MeN2oY6DM3SJw1QfDR+GqAtt
LNlFbSSs7NQBpWPhfgxPkiWOqObnbh45fx/PFBhmsY/HJUCraTTcSms/CWpvnjRt
AiB2v0mfl4vuBQW0t0NxNGgqXfdD47eoccVWVGw7CC0tv29+Rh/N7msn2o6TOY9Q
NpAez+lmHo9N/7Vb6KaajpNQj28qaFW0UQKOAHsf5fG4w4YJ7DUpbMr0DIfhDUTQ
YEJ7MogAUdB1drvnWZJCI6Tq2/4mSAHNmGerR2F9/tnlNlkZwdpJ2bHwV6mNWOwy
mnS/1mM03c5/u3UUY+YBocafqe/wYUXUnQy/B/mo+fJI9WMH1xBjQ+Bhtf7BEcq5
yWf5CIaI08o0wX+31kuYm+m28iGROH4Np7NA/WiCzD/cKIRSNtjh1i5BPvVJYUp8
6xsmA6USoBExl96Pu3VEeC6ZnV/A68Tc+W9OaOi3ZMdn3ITDHFNlHiCZCzAl3rdT
8tjb8d5/0HewAPsXxVI0Y9bzC1BPUVRW3WWq6Sz/GOPFPeZGJFlxg7NhkLl9FkIV
PMcGxrsLuJNtAWcD6vRSbat4s4YkZP9x4h7y0lOxFOUz9IPXI5Qbl0BJBzx20DB3
Ge8mCgibrRUt36603Xjq7GrJopSZHCbY1YOX62Af4fQ15zU/OMZ+KC0DDIgCOLzp
GuLafXsU9EC508XMCISve10sRwlpJtxUoScnWBfvN+8sNSnzAUnaJGJvD3it6E9e
nAy8s8XM5fzqQtXi5J5XFcEgBVJrxVD606ZkcB4mYRufp1KKrEn3dNV6qRsHTSFV
H9yAhvr50K0PYpr0UYZH20jcN8SqyLctgY2kRu6OUMb0m98LhE86AEfUoQDddNpm
veTPej56i/9hDwVcL7hdkEGPu82iuxjekuqAWyGmRBMXNNgzcHcwUeiT7QFpiLqX
EvJ03nORvH5EO5E0Mcc/RiwbZFQhTr+r9mPP09P2t7uVMGPsS5vMOg6FBB7s/b2x
CTe8DHGqjXqaXmBCUv/PUgqZXAGNa/2RXpV1GjOcRLPS4W1j3bsCzzGvSrs3mkZy
19lkpyzxPxzlQyuMgK4RAD5m4qxi3wiiN/IHRAlpSrZ7XaU12Ov8XsGH/RPMNxjm
Y35vpSFOqlA6PxTin14qnYOCvgehExLg20BykTI+X2Gd0T6ROMEPkKGteKfwvPzI
OwGmtl11y7xhBMyoaXBxhG2qRBBZ/xXTl0blCQ+GGUbSROvYSa6wUu/XfKPrypFl
t8rYmXQx2u65Z/5tyFLpaG5bFPynH5Jj+Bw7Vu0iJDcl2mK3rQnfu6ARzidUS0as
D1bLEaDV7TMNnRYvqNOl5jU0aEI/uknuQqbS0NiwplrzZ0UQXQqnP3+gNMcmcynb
cwoN74cCR2uJ7IeNar20+W/q/eu3R16C7DKnfZ78bp24oMOnlcx8Bqj9m15Oemr2
F3vCECEiAqzti4NagrZgJA17wK3F465nrbIpCZiGWuTqZeABRZAF2jslIJ38NmXj
ctds6PJhLGLHFUlvljIFVp6MukuEEQCTe0vp0eHxX6tdR8U6IopQxJY3omAxsYtC
biOJL2YmWPhP4xw8y9fE1BMHEYrq8jt8BwMTX3adST4QkA8xs/ttR7q8Xj0X723A
l3frl5ke8Robo3liUWIeL9aO5z84Ppl3fPSxs0bYlG+Z7DmmmlScz/2cImtWaluK
Nc0vmN7f/1pgrR1GMKQ4AxC0n4Zi1S+vIqE/FKSvVm/ZEAmTZnl1hjTM21Qu2DEZ
26Kud5LSkjDdilVEER9nAg7F00oS64yPWlc0CHvpCHapnYctma/HTqqFQUNv81QM
mY54w/oNjWLmTODZpxc3GrhXsTvBGyw7M40K0IKL51VdG7Rzd6ppFzVqm1/Jl01g
qlyhmXqt/as2puPpQ0YP5ByyT9oncq3u2KcoR28prIz+N1s8jZmV75//UI2sWuk7
C7I2E/qbKcOmnTsvE0cU6k/jjzLcShSk/Es/I+gXqRQu5aYVOT95Z9onUSDtg1FQ
UQrSDekPBjXAWBt3MsNYvTQPHMy06kUrCCl3C9m9jfq6RIrIDC8lkXw4Ej5Uzcgd
6thRv9AoCMv9s3N+lMvlr7rJf19H/K7j7j5lwuIwsnDm6YUup7BFEVmUav1pLJzH
t+tjfoW6T3zYJYpgEeRq6pA50+TeLCbtp60J5iMTo5iP4uUylXivoNyILM/SKDAq
FkktkCz9spOc/+HwbSuoAk6IeFujru4/jtN0fXYN9Z4K+1Shm3PtFvBwJeQ7gdVD
e7EBVAUbUTuR8ityQ9DXwmXQqrZl8F/m6LK3hmfymFBwvnyKMXPIxllAa5Ka8sVl
jTt+X0VvOnMKWXwcrlnZG7oS3+vDXIfAL6qBgXaAd6qutFLr2/GlG+qHHY6rtue1
9X5nqgSfazyoRqoMDf0LkHprfyTuyfnrOTqhVP/XKFlirQGxSuuWcVOSSCD3WH3l
G+HwMGWLq92ADNBs+3vCZngyMYI0I8aT36BLdGOkT+5BDv/3HDn8qtlGujnRVOQE
XXIvYZE0BSbrXW0kF3OXW1BT9lj+Dz2gbiDOyUS2AwPp6M3EsBIxAsUNRxTKdr9n
oC0V/MIklfZwFINVvvke2Us3IFmhjtxZ71Wjn/hiIo7AwZdrTIzvBBVDPEqCarMv
4pMSRz8INBbLoxoiul9o8bqYn+V/GDRi7iXWAQ6KAQQ/e+JcXxcwuX0SPp/UUPFC
ijL/lLbxmcUfpc6wMN9fQ7/eAHqetCR2wNi0a7rOftlZ9jbqEL4xzkxL7Zu4re1A
imPKwpmEiPt8kROAHH+YlwT4CIvd0Y7C5E3SXV4C2WemwxLUpolV0uzLlWmPsSGC
gsMybyd/mXEG1je2Go5qs9mapx6wB4I0JtvYilgsPlPyGyLgRR6B+LSn0ZC9nl6z
jnBKMWAePliO66rUmkcI7P/rtTq9g2wO0H9YEk6oiceWOygDJ9fuiSFDBZtO/d/O
NUFABiCW/COrWJddKDtwVl6HH3vzszw3zcnFrqJpA7IAXkYybmLkSb/vTMRazj37
EunOU35XGEjHtbb1cWH0E5anXSzy1ncFsTL77I1hoibPph9xetQbButYdzCZSqVG
cwLLVKAcLOcU0PbtxdWweDOVFIdh+BLyLAoDg3YNI89Upy452z6nV9tCUC+v+5RK
vNDswK08D5HtO42FUNudahfRYGyudSW7Tv2EpcKXvpC16afE3djpUbgDTU/tmM/j
WDsPkSfLaMi6c+fscqBgSpgG/FRK21sS1r42pkWiN3MmsqBf1UnbMq18va9d6AWd
ErognQ3FpMi0a4Z3mJTkT+Ig4OZU5xnj1KJHU7gauCLBRrDVTpzpmFOUhQqYBktu
OhGs6vdrO/tTp5p7d3/J+n355VRU2MRuhr1JXou2PRFawqdCebCJ5gWkya/Zuo5l
PuwVF0eqpxZ/ukNYY2ZxsLtk2NPKgdojhkoWMHBsRKbHTwS3e42TsWEC2cPPFlnJ
5gp1AZ8ruTm+743A8lvccxPZrcG+VjbfgqNhEWYzcw3v4EWFPnAZNZcgYVdVXUBc
gQ0uxpGhHLL8R2RSovFOiAgVqN8nereSK1HPjrp9rnGQKmDkA1qfHsWn3sW8vmUn
Dd4vczMTx8+58ge/SBOj8FP4RvAcGGkcq+GUvwClSl5Ky8Qk2tc9czAwxfUUs+4p
X2CfQM/U8PHt9EIG8k7CDChOJF8/V+GIzQAiuTyNwmVOthQ7CO7194fdosyOkaV6
x1s9SwdE0PwXXx4Bvex3SpfDrLqZUfU5kljBzrsyAlFxxRVSxuTtmRQ5G6Jtqzc+
QYrSTGLZeEqzSqJtfTOraGAH0dvx+Wxpm8vzDlva2/C4VFTr724SAeK915YSUTY4
Rxyd3sRlvVnWFa0jJ9NR+VvUifRM9amAn0kRFayytiS2IK1gTvmWDp6n3qZmOGCS
Z+AF7pAUUUdDKZuCp0ewyxLmL/XLIApfY18+37xppgJP14S8+DiQV/BDH/9JEbYs
Ep5+LJ1CYFHLnAMrweqkH0Mxe1ig4Q5fOfy3iEIQS4X4WPR20t9mtulagU6+OiCR
bW1KDLmKd3s9VDcjekiRm+Hx3F3LAQXfrybKMgyr6YMVzU/qIGMZ078VtwxoYN8X
WOgeQteF7a7ki5ooWJrF1RrBChTKnOB3IxekIl8GJ55cVYclq6QUQA0CDMcpPR7e
WtqXnQDVNMEbsuogX2zrTzXKhbexE3BFJdMJTjCRK9D4GLqaNDEPwp0TaJ0BW1uG
HQG31JtKfoxO7a007kFe+WUlHZO/PqGTUMbsLm9BKOCriacayjH7Ogexk4uJil25
sLP9fBYf930zizBRhCL9XFHzE+QJ/90DCqo1pXsNuMxdSOZq3Rq+LicD81XKc99B
CZk2ZbP1zWp1FUoTjC6+tlG/gK1Y7Z7g1CiOtbkbFxHv/AAwGjxzgFz+CMx79MSX
yKcElrUjszJTBedInPTb1RyqfGkVT8Fb9Qq8/AmoH0DmdYC8+OuS7w9XOlth/6We
HjIWQhdEUFxfzihvDWSTazVVTjHeDnmWC44zEeWrMvp8uH0a1WduUf1+LAfqrxUq
ms8AyWjaj16w3nlpmIHVptbazM4qLNXBGbMl1XTJywbfXzlFItkYvw8YtFW+hilH
g35OYIIWKbI9XGRVgZRkyHC1K762mLp3VzlWfUKdK4DvNVaFCZdN/7XHBZBjL8qg
EN2TRDA+j5pPJ20jOIXIEORBZqZ3JtlNSSxICUFaI4aEd9RDgN8MIxebdW0R9qvB
g+DfPkl1Sq0dLvSMCJ20QaWIYzb239RuzOhN74c7KMLcBQOriuryTz2hhdJXqPmS
OFKiPzuhYyNiFK11QYK7bdErVH+yERYP5db8CWv/vFdzGES+1VE0uzMJZSji5ovG
UhfouUpa8c32yYeDpRbS8bd3gRPg/RrweWnC1Bt2ivc2HcR8eLgqZS5Ua2+20Evc
eJY6zTHqsOynrZL0xDfZflm+Q7O7nuKs8eN6WUusHuCBGUdKZe0RHO9BZGsBUduN
xTFSUnv3yXK/fpMvFMYlKy2zqd2pUxUw4WkImMx7ym+Ft+NumAY5DpteMfaDEvEc
iAS25SNDmxqEnGzvPv98rRArUxsCqvFKuPbJc8COr5od1bMsuNqiliTHvZ1P5hQF
QMYA5e0/0Vc0Tt3zcqjkZCJxMm4971HfRk5yEeKTo6Vk6VrBAIlu5ceUfybDc9PH
3h95+O8IOfjz93mEJof2+pKF57GREGV3XV+modWV5EOK2+YNoZcZfS880UhdtQdf
5bPsQT7JE4ibeiI14za17nwULz2YqtkPkW+DGCI905rPcbRn0PiaOcZw6Fzs+UmF
wS5thiqt6DAeAw6pEbW/V/vGKfSS1q0tHiw7zMQcQYBK7NeXeZgjo/bjSO0+FrXB
Sytjn9+2ebA8k4P7Mz/GsSMjL1puYR3KNdgVitdzncij+LWWuYRzO1cDQrzldPPF
kf5Kjvjd3FNGeESbEEwNMJVdLPh3a3L6pTxM/Pjtu56vWETYSzmxkowZLHRDvZYX
c+Lj+ibch9SD35kPJsCKLlvTwN4LtubG5yUrLiJWuG+2Xcwfr7ZnvdGBjGB2pj2i
JqBiKelkzu8DBUQg8/INf9LVSdd7d7TmGjyigj9snj3H3Dw4pMACIytbDO97e/O7
6MmgQk41PpXpBtp/cn6fgm9zK6YFPQHHJ4V0IyYqAD+61QNHcdVnj3VIhowfoskJ
23frisKW7f6uldNrqTB6Y2c2K9+n23KX1rz9e8pmk8MreN2P+5j0Dz/XA6b78W07
50OkKCVMKP9jX0eslek2/g55b9kqSZ1poJOLJfhWOdNDZRSihuvg2/9A/co3htTP
hrsieho7gMUq8/sLtZkY3Mf77SLrthRwx5SMqi8N+TLGhh81/mo2o53/APxHV5S8
IBxkhjqBcCMd2bVqEoEc7jCBG1HmUHjoTPP6DZg9hcFnmXdy4tseicXo/Ho8chFz
0+S0mm52DKjlIKCARnS8/KAZLXimwcMk7vbaTFJVE0KLzn7kD9ThkltlBGlPzIGI
tXBGPbuxkH2eS05/+7dkZOKtKaS57YPskRYlQiuq+vrQXh5FWbIbhm1vusYE0q6P
Fs274Z4tH2YtrCZYLIB6S33uDUNl+O/L3rbsTtx5N2O12UTiMV5xEu/lokFYNVnh
vO7g+eYWMlwNbLVp8MElK7GsZsJ16/CIiBAddxT6ivFsGPTUdX6vkK3L19e/vhfT
DyiE8fYADDheBiWljLHXHTlNMySmJFFtb9B4fk70OJ3cOK6BAafnMR83ONbafjaW
RRTxrOun0boeUIsnfp379AwCtYghfniBWDwUmm0GqBrLIcjzw4qlNP7QgAjwT2+m
iY2TSQkpMD96pToV/noJ/O9q839VFc2JyYAOe6SEDr/qZBk4pPpICYiR/tr71QA7
Mlz0sqaXehjIhil5ZaAnr3GWa3zWgMY4FLrz8+9Hfj0uAUePaZEdvDUQnMhDZ/Ix
uBfPtHzoZwlK6vbp+CWmkgtkil1P8Q+BTwHbtfpb5HYXPXUnkvLZBluEjuKbJYvD
ZmCmfttTdAKkTPNosMLllujAxf9j/yU8WGvuK3dilTbeVh8BBlUh92dTZH2tEqLH
6O8usOK6qvEcl1c8eUS0ifE24BX+xI6B3VCApuL9Hl4v1eZ9xPKsK9boHWR3Ee3K
Ei2WxYTG4K886RFgl8icCOKQC9hoxY3GIaaB4aYf71YoOegYOHVX/Zrf+ExWNdFE
4u7NhjoWcTdKY06pjHzNqpKNfdCiL2Zl8J6VAzIfjG4gnOyjPe9x/Tfk20/gA4dQ
4fCSgnvgWZjjVaz70QXvHYxeYn8m7OGeHwxwlMMYePTZlMHif7Y9yE2dXCOLCFSP
Jvq9qAlFq8F4wbX9x5VxlM0OLO+viFAEbVMyTG3wdJoQm+r7DbXIIA//iRVrPeO1
ZGtwPdMJkF5+6hjF4OzD7YGEsud+5v1zi5LVhfvQYBqAh//tg+RjcDba8L7HH+9E
bBcnh2BpKz321p6WGSbfigP/v6DIgiYf4cNs1c+AC28U1POFadKqSlFwomOOH4WI
ujE8reWgVb2a3KIWtqdzkNNjINV0Pfq944e/OS/N/L8lNXOTYj56dfYEY+qDKfA7
pPz/jpa4y4ZpmCny4lsPLOR+kvILfxack/Zp4q6OIWUQrEpAtdEc3kTvtpYpPhrb
3jhsQy1rfpFtqhlwX8frmxUWe+IYUlt9fBj/bzZCFpYq0CR8JrhrXhHLmMqfFM3P
fgNF9mADIarrpLJdG05K5WVgcV/q0iYuXOyowShd3AVpBTSZaLMIlehFpCNyy3EU
DltAxPp+tT64xro4I58E7UYgdmABs9nuKZb13HcmThF5zsNE54kf3IWoZUFvRas0
VhRaIDMRcywbfUkUPi25FzMBWq2pABq7ppJEaoux59X17ldl4+Y9+Q7c+UhPw6Dg
iLQu+0+hnIkMc1tZ2KCRTNg9Jo0rDSKLuvOWYh0cs06oM8f5mX5NNY88PGKFTidl
0ftQnmm2+D2eVne8rFl8jtYQNpCzmH01+DaJByR4Eo/7yl1i9vYNKKQIsJkDWvMB
GKMoM7BS5EFjwzPHfF7UOV/XfhZgsI+GgAVNp/rT9XHBzWc1p2Hx2m2RAXvaFiTF
prf1aXdaDbWuGhjENXzinkAwiMMBfIH0mkxxiCZEWj1dXTJT9lfkt2riYMnlPWPM
YLWz4d5DeZ2Dluq6FVrGMgD8Ju3RAZIuP+XOuwClF3z/na6bHVWXU6fFyvjAS+Jo
JEtWqNUWDW70gmO3JoxvHqc5BoAPHA387m6eR6qTOwpnAoD9nMUlWzwbvbggYfn8
NKGWEs5HKwd6K2AFkot8LEumTTvtWD5zdGVH/mhOMhtFs0Sdwf5BymvRgbKjfoyP
DM9xEAsiplN1j9Tzow5/KRutMSYdz8URt1jz1yyh1tIiPjQRdUK/Ker/iFt2O7Y0
qK/jw76jnrHhT7LjrOXgkjCEPj9YmniIXTPDyKhE+qzdW0LvJnKCGgfZPHTvWrOM
yUFhPrd0OzLWpQwRb4YOmdv7fP6HrwUijOslW7CCagL3mYV7PBvsceVHNhGlIn6m
L5YjT/rxmRzuOZEtwAp+Te14taGOxo0MBGI3DQxy0cTx0Hx7TEfqgJ+YVrtn6jsK
e56Ac+D7IYcwHvU+jYHLW9m9YSN2aT/W3XFLrynKqUimunBbK+hyVcjxEPgMutlx
gvZ9EtYOvuv08kMYvw6pQ2CuWA64kq7mhBkV89WGdKcq2MsQu6hm4ynh/htk4rb9
P2RtBapPZWnKF8q3sgIqXkdmvvCJzTYUu9cuRxfuHf5XlAqdJt5NfAB+jEvRsBzM
JobzJt3CWsyxzTYjaDdROfOkk+ES+OsyzBxvSY9rtBd/O3iTntvBByN/c0Bn+fte
ijd7K1id+ScQZSGrdeo1+MsL94erz9+EdjXIP9Sw73C3K/ThguzVHZ37uHGbVwC2
waHiYE2O8Nk4HqxZubk6KrMg73IDQNu+n51upKZb/cywpjABtykU6ZmztxCpDh9w
mzjBI/emtgrflGOs4ejuvSRS2UD8sN+UPSDYd1lCpsiMDuh6iQ+5vPe+j5hubY9Q
ZDaXnukU00byV6781VKkfKAxiacJiAlZbz1hdKwN6I4xwBBYxKb5flIX6p9Qdlez
yG0YS+lalunRE6InmtmOWOSLBkz4Gp/VnayFaTgnhQ5SZUXdm0hWoq4/Jfp0/srY
PKGCejjt7WuSL3yPpnfUKG4S+gdjbRlkNIA+eaKKSzTXlWr5efol5zO+DvOkw2M1
Xhhrubc4RnJ3wv/5RVHy8X33tDWXWOAP315a9myZqYateM01njVdWBm8TAoFEsyJ
hwn4XRFY1RJhbK0IC48dNsxbZOg3p0tfIU9LMlffyeuXfAYLJIR9+dD2Kl7zhFSA
s6GM0h/Q7ezJYmmYOfhp8VPoOVs90gUf/XpzUTtSFmrIoM+rbz77wbKgX8q1Ujq6
/6m3RVgD9CVHjpG1BNB4v6a4MXabQ0L1yG3qUNgqXqiOY91z3c0IIeQ9Bi1LrZ1i
INhnYrosp+/rSUbGcAakOd79iHAP4cnrDDhlft3PBQlfJR2oVxXl6oy1oavysrlX
qeAIpl1XeNPGAZtwNwnr32W/7U6DP9P2kft4KdyST/bgFtrCRQYUMwbpUeTaa1pE
m8CDxDd9pAcaUlCa6HuPXqq7DYEsrtTBPUZwt4iqj9yPRF65tn9TfqXBzUbkNrD9
OSgm5bwABDIlUqbrm+anCTph+atm/3h/qNEEodWubvcVoEEFFMHHgCMpAnYiU6UJ
L3S7IWLC4aVI8weDUdBcqhztafssJeuMUMaxQ+6Z4xPD8yeO1fH39yIsdts1Dfzh
GW1SRVEQrf1i1CI1fw3gZ/yNaT7qgND28ykLLi2uQlQKge0VW5AIWXJ0TrR/tSD2
B5uv0Moow3celSXyAUSAoBsxx7L15rHJRfwzYkbGhQO9Gg0wQlioPC8aRHGGIoDK
Z7sueQxWNtSm84xvc4PnAS6oqRg+vEVTDoeahWx66nBx86d/HuI5PjInN9cnkxY8
OtIlM7zr1kfQanGjUdRPu2sGxH3WkAOz4hncGwQrF9xOZnT/V+eI3F9afwLrKSLk
DP5oJWN1z70HkVOuVMkKq+yZvqrwkQnjuJRoMXQElNE4eIEux6v9G3H6uFxDjUci
PT2uS8fR9B4kuHekomFfE9AfjAT0iIGzk4S/6Qg6CvTLv2EbNNbA/nAm7NydlSIr
KSSv5RpcqJTp5KLltXtp0sBksM3OrZgrdzWUOQ4pWILgDVn0kTlz62xfVkYfHIzK
C1NEpw8+xPKNz/CTXN/JCLQpzKiuB6mjNdDEVvxyaNN4R951c68uyTxBkJ2iJnlw
5UUDaR1P4QWghFK2kIlQCWpEkE8IVziXqSQgOfjMtRK/N4MyeRDWqJEwa2DJ2xJb
v6Dc6s/J576c5X7BclwJgGl8VITwPWlxtGZACJ4l9ussbXot1pUQze+k5X0cSzcK
1Z8ydhUqDTWvVAWgMOOPVabrDvuxaaehghIPm07XzPj8Zt3pRsHPLyTjBrb5VrR4
HmN5hDG26wtljRAmWNP3QtplfM6TKKN/3AgI9dq3HF087kFBNhvNVvt39nv104ly
0NQ0phS50AEU/seVDtUjbv29trpSAZBXqNVZj59LXuuOw99zQAqfn1V7HyYBBRVo
frIuSKarghBFdP3HzYct30tu1oOtFWTQph+VL6jp8OszzJCu6HYhuCvuwtjiATY6
ZkUSmlufztSBIw32HJED/4VkSBNVmon/HZ2MJjz6OtTZLzgMoFubEBDHFemrAree
rHteNW9jOp7F8Eu8JRO0+ldx4IOD/S045tnsFiVsX5wR3niUr35sYdMVTVA+tXLy
NPhYPhgszZ+XMcK5CpgMDzF1V0d89Mx1JPH0CIC47J5QvM1smkHXLzvOOo5cvR3G
aN+CwtqaPIo5dYNg3eZecMexmFOC3/iE0IPOFoN2/aFqllRVjl2sScGKeFcTu2R1
K6xDur4HoiHnYEsO5AEF4JJikG8AmtD6BRHnr6DnkA0E3CIGxF3rlJy+l6mpLp37
exTcxmCIdyLfLI0JVJ4SjEjoFcLwQlcbwcmcQi6zTxUQVsl68udM2QmJsxR85lml
1vDHku8qTuax/Y9lpBcVrzMD8I3BOUJP0ld9p3bkV1DWPcqEQaTADYINtx8u0txf
EbxGPTDKnLS1Afw83kz8S62ATQmikEOAJoMvSW7P/X9sNyydKp2doK34G9O+fD+O
c3TdvZkAK3hqR3Ihyq1Bkv9JmCBQtMyOuxpS26m8xyNQOFW5X7caog742RgP2XNF
9unXt9O6DxNGsguyuXgqt3nNjAJ8f1oOK/SEdP0STvxAyL8V7Qycflf55lhlaEX3
vPGx+jd6zdfAOCWwBZh8sfOLXnfO3oh2a2VpjTLPPsXazrAqYB91v1IindDN7PGl
GcFx+9xuhIIKHLfH4rh60Xggo8m4rZghv9FEVWyvOq4Nt76w22AtPVOmddv+SEV3
hpDIEBXe+N6sM5VjZKxJ29zAJcnZ4NgZSodT9QqBCrSSnZwWg1S2RCSkjeHU4JtJ
owaMvS/GLFOAI3FQZs6+AN7HNaw1Y8QLH1mnQQksjsia7fLCbjD5nvaSiPdhM5PV
WYLDgJje1DZ62GgGashC1JwTML/Ngy2Q8bYPZPxEWYjtHSibcp45Ikicg2StzEou
gBXTgEQulGDfk9tYHdwZLcKx70hbUVxpjmlxIFDiwYJ6uPHMSROGxECz3jw38ncq
z3hyGHvpFIzKnnxxOprkO25hhDuSVveX29hCp0V9MwBV8llS0X6tfnVjtgDGAvp5
OqkIQLF9qrmXVAmlIku+4hpLNDfQvP1y0ZVKKDO/N28z4TYvdH0/7+YTuSDwAFJa
sElm3fOn6VlHf5WvHZOOgWcdw5PLm282klqvu+Iw+n+r4UZFo/9tbf0rPvY9oXaW
S3YBrPlKPLGLO4idszTC4pWNGWpDBvSal7uNQzX/7OU/RDJOfl3CYvyQJnYUmOOD
RfRSJrAiZnT1sCNUVQJZkMjZxzgDDW46LuLPIW30KQ1uvQtXmJCJLaMZrluubZ9A
b+zGXEprcnwq+bs8PEypp4s4kuXK0x/gopEsIVPl2BZGsYD9RpsBgF3sfSaWIanm
dMnNGheRVb/uI5wM3q6FITdIZDsic4iWQ1Vejdkuq9R43fHNSKwuAkiexDPp70IS
3O3C9l7yUrUp2Uz5DvqT30YDYiDJ4Sm5MLlk45nbA5TqRBQLOlGh53wEixASGReE
HWxx7sNkVsD3e99cwvInIYM2SyTmQyfud/0YOh+iQjeU5Py+fZw5YGglk3gEFCPs
tvUt0RcmAVk+S6mZCSgIDuVAuFALKMrmfTVgs/bRBSRD2jtFlCcya1iZDEbIO3T8
XO4C2LWk23Wb58CZh5T6vlejRFh/R3NrXIikPcUWWzS4DZ05ebSmohFaAwbQ8zHv
l/UxNLizU0KnhWqEMqPhaRX84hzQmVwKEYtXiqnu0AXIiiaqJeN2NmwY4tJUDig4
K+U4/KJC8p62n1EX/DSOAJUm4EEKLew/Zh2GmA8stMxx4Y18q64QPfIC3eTUx7b2
Iv/X4yCkxyfxP0sLjx4/CBIrN1LSvWBhKzQWeVR1JGRNVwnQrjHoD2jurtfyTigK
86p2HKEHmtjh3fRHdpqZUrewxNJHBXyMKLy3gxD2eHZfmkNReKlzANJM6Dwl/SNU
Rp72j8pgyLXGylEtiya9/G6VyUzPov+NJ3h+Ibw+yYm0KbYK9rwEDU/A00Bm81wK
5/GeNWLGDSILzulkp1i1XBr2Pt0NK21fnqEPNUHPsGGSLGUiZo9WM3MlcLnm2vpH
03Q20fccNcgemmkT/4l6pdFxeaUuvi/RxqM+FrwmCfLiTL0Be47Jb/0UNu1M+N8P
X9nK8v6WuqY5WIuA+8/qc6yNpgrcFJsVlLdKuzT/IAPvZCdu9uM6u06xqYc9vHGy
uZC2K+uF6Uozwc4LLO1Q2D9XHWCGf4E64u40m/z+8RwZaF44Fnv7tjkln+rhSNIO
C2vie1Sf54Y7e/4cK0yX/1goQjAUNFkyu1u9rHAWasoSgldz5DnwMl25UyYjERz+
eMWdOXKnB+fqAlMesKLsphuAsSolSSRc+LWdlYdaCquBxW2f4scCy4IQ7BCoSlSg
Gz7BXWasEIX4+5EUDXUDl3qSPjEKhuxBM4Tn47nhTPxpjZ9Gz4HplAPS/QORgsIb
rnl6cGFPha3/tr9k1Aq1yfCAo231tZz+I5mtbuAf7hM06IxMhmJv+00871/nnLbD
rZR3DGgmVTXZRxWhTNwH6PIQsSGQ83OGpSOXbBmL3B8Vddasp27K0bUHagj/L9HE
AzDqKnlpyjEqO6QIpiNcphXX6xXEicDApO09KI+yhSv0AIJTs4QxTkWWTgLAF0z4
IC/H4Jx03NjC8wrTIoJP8fRlU4tdUqKRIfvWfZTawn8QkwDCsrjNp9/ryPeFE2dc
HlE20ZTfMA3ycKv+5KGOMWIPuJkwzAXKDBU4P14MyQ3q/X6aOcfAzEVTgHlZJAGj
wFxfUIZbHS1zztEC1C9D74/TxYdkq1cqK649MqX+ysN5iTU4/NnvvM3h0CPH0/uw
akh9waJjm8+Orp472oudHK7n4yFcUI8WGnKdIrTIkuoBJV9NYIPH/0E22I0cavZr
2+22A4VuGI3raL2B4HfB+Ccye5hY6HWjJSDwPmiDAj8Qt6KbmPeUEKYw+kExOB4b
dWzE6ndEkEhiIdQ++IMeaqAAc+/nKhQxxAXe41Sey77QwkjyvV31Z7bzPNDOy4fs
uE4Cb7P2qe62c+FNIem7brSkhFzyWgn5FhKJ7dVubfA9Bs7wazrUoTCxtK652opa
/6FWpC9gOqxkvTCVRVk/jw9nPDmIpVc+hTu6q1cfc0ITx5TH8A5wdnKuPWEYGpYz
LZsnHs0XUO2VJ0X0gx8uY+O73w5uErTJ+DQxjsdFAJY8fW0UP8Kz4/VzzW9MMfiU
vof6oWDySBJH2LK0G4Cnn0SbNwGmPQRwLGaUd7t+hpoZOeV68MbQ2AlpdwQtwIQX
xTtmZQSUIudiGMS9QxMKLhnv2ic79TtKQCeZ9ijGtu7TceeS5K8kWaI5IZtVnzY8
IHAGrT+46L8bGRKdgiuspXoQ4AWFtv4xvxEvKnBdyzwQBZ1O9Vpcp/2CpRr+WzJ6
J50dd3LJNN7iey88LmBUjE4kReTf4PfEJMCI1psO3j3PL+W4YKFVX+7QeTifCYya
ld+WQ9ma2QlcT0lHiksDlqJu0n1/hQ4fHEE2ZwPLoeTdiahQEcif/Ivxq4GPn/iD
mxieyR/55YGo3PayHKvC0W/xG4+zQ7pXWfSpcs/5LD4oxEnB7fKeARiclAH1667y
6zVsp+MFJyEYwNsXVl3Bh8go7e3pZu9ia2V7YcBlqKlWzVfBj+gTmjIUXi5u/Jux
chGOsYbRRzqdrOBk1hdpYKdJhIG/UvbRdfAZ6LVSemFUk4ygN36Q/eL4G3L1lpsc
hGyVahApjafYcahhE81zzhF3A/iNxpoks5Ro2lSuyIWijk+jeRnGO/JJGrKcwR2l
dORtlr25/NxPe1J2IsjJTFskbGFDEVd7w7T+RbFIOSBuCKEHwiJIzT2yNiPrXuug
0SGFm3A9QGaSx2E1g3Img5GRBDyWPU0uI0H1XGdXepDFSF2KiCPZKbrGmB5Ty5Jm
OhcimNvZOigre2rpNKdyc5Tqt147z8FWfmJNWraza+SQgnE3xI4z6zLW/2E5qr9R
Qp3soC4QweHHYeiJjVFKGZ7gISIZkDCW1pAyxhTxAe91YR17C4otdR1bMAKaaKyt
ZYO1DLTJfpsmRk0dpl+vTYqmaTyVPMjZUaoQf1DEd6H9ZqtfwfP43Hp38olEQqdb
axnp6OeHb9ksGc2EaOmMKKEr1H8+NV4VJ5PGGCJgGwqvo+eITbQs4BVZuhP/8LLz
oUrkgSuevy9hYUtksHrjfSrAeUKgMA+aOPt7r+mxpCBJuNJTcyXEbWuDnmwHxVhE
Hfar5I/j1fWXRBNqjA/LM7T8tM/UoCkuH3+HnrrRm16QexIzLvsn16OOCk49u9h+
oY9MTkA+Mt8JHyBFFupNjyMCCjSUpuazQb5B3eyEfTqDdHMlEZIdXrAlNHE3Vle2
IvEjvZzYhM83IQHcwx0YFJ3/JA4XEYcoXP2RYt1e43qAxbPOPKPGufUpaYDqS2VX
Hs9CTSdiFuoJuOBsgPc/ck15aC7vUblU2J8gFmLy51RgUfZmGYNzq2e2Qw+82/Im
duGPRsw/cbGmJoLOoiFLozxXhCY7VzTrKGjwcMpS1KB1aWxKF8DgpglOYIrGx6tj
FNHjyJujHIvuYz4SxyIOydEAxNBs4LsFcVQ5oSfXso4wAAPIpKLZCSderU1/Ide/
QCc46dHAOl6LYZU+g+clG9UR2EMPFYaryN9IGjYuueF+Ob6je8bk/AdVKCa/zMOt
WZIepn0wbRN9dsanvt7WMDNyR2AMK9DPXzZe2VtHROgeT3ktQ+o5LX41cu2UEv0c
ti1lu0jIv/nIc8xSxaj7GOiwLtf6bQwVlURl+HGztVNthfikfj0xz4CP33uEVGB7
tzNKM4wW7PetqgpQiPIFLcPRUAOGRUo0iNPm8JQu1ck4Iu6jsVbhMoedG3TPk2/o
r167w0qpkvcZ9i16lmKXv5ie6JxiA+r0OXKfj4eqn8ojHOEB/BAaRgnubjyl887b
XEMLRPlAH+n65SmGZwBemk1fL+ADkT/crubTK0mmdPxOLuGT6XYPr5/vmnuieEqo
4oGJdsNeKHQT56ymzrdwGZsGuXreVeUYr9+AXrlmrF6DfAPAbN+MbStla15OC5ZO
mO/+dRndr2TDJV+NeAehiFNwwtvymcjKY5KFcmRlegHjG4fpmc9a+5gQ22449t/2
Tcu916jikDKXMfwZU1XJXAinsUZ0Jl4tjujLsTfMYJdBZHStj+NMSgQ6qQ4Y041z
hj7Q0bFkLCdF80dcBPC7onp43OfRCQnMDhdrcyzWeh6o3F2RHvW3A1RhZGswNR2p
/6+0XaCXXpPoc74D2oweH/i6BLaUoHzrhQv06rOtFSc7RycyGBBREnGZMFydGTM6
uyu80R9bijWFsDuyRSFA8T9ezuc8rAP46oWI9euocV2Jvv49pjsUIdpw7qJfc5Wt
+M78A67oDohKH7zYtnvZoTea8vjv5CFlDqO7bEpCCw4Z56UkeIwF5BndisNEVMe4
cE0Crw6VFMaq2HRzx6cuXPPjj4H5t68PusxWGdNRrNOXhW02MnlCgxkTatOk1cYx
D75z2HeO9ubFckp82Ny3WkuXb8MHE0CnWM+3XU4lAogi9F/xdx/o7IlzGCO/N2sv
SkuevRfJVhySs1IrgNVfDkwMNAToC5sZ8Bt8X30esZsEM/MY9OEzR58FrYbj5Jd6
hl6RItJd0NjN2fV5h/fndKwp7YDKckDWo51Ha8xppBrlHEimiGAh+3w8WaauUjtW
mwp8Y1c2C1779TAYCTyyG4J+fsYdh2HY+zKv22kf4MlHkNHS4djWtss7GpEfPedZ
aC4KBfD51MucB7Wf2fJjGlc+izj/HhPi1lspVngKzUYbGHWtW4rJZ7akowbSfRwk
b+AXw6/dWdosq6syxcVIiYNYKb0WFkXmkUi653e8S6k3GtuVwTpMolhjU7BNvFY7
vvniFG3h1zMKxpfAByqeO/r3x4MGQpWBg1zV2DPy6zE/egfFKPhn+gl9BpmNgz7K
dxNDLwqXYzM6D4mYSJ0CZKEmjxqSjo0gq4qCZpOtfx2EugnMIrUJnLWLrAjjGFv3
YbvCS+b9P5JBDHS/4aKUCLl+FevUBpox3mqt9H5W2WNX3b7YfJ3UH5VPX6Ym/Lqe
/R3JMcJCfeaRQOPaPrKg1y8d5UrQB/VPWlhwGQRvBEY9+e9znuBLcowdy8ErR+xr
X2aQOiqQpy30SRIQiVHy7s8zwUz3npnMCtC0RDbFO5w0ngDWXOExXVwmVxtEzTc1
YmH30aP+MXj26WGFHA+imvt4LJlZQ/fbD/QusTpm+CLXGSGzDtWaLiw31rkngB3W
sSlor7R/wAYa39WVtgaVXRZsYGH0eyd3s0u1msgettbF72e1DgQvZ8Suy5LAz7TR
uSy4U4DEkC292Mof2vizFdrI/HBepMeiC2aYR1wKzL65xLpgT8V1/bMXLef2jBrh
VLyDYYP2lmrHfYCfze3V6PhtMi11e04LR2p6n/OEBy3cCGlC2dZNkKjvUsGWiU32
gq2uz5fDbvbnCYqUG2kLExX/2CqL3KmQvAxkTp+dSjirHy7fX9cQwHugaYNKRXoM
+UAz8gzDfSqV2xekCcri/OorEkaps19AJ0kdJT7kQlBIzHPDVfxm3UbOE1fDSZhL
3H/VhOt5gV00AUs9P3uIhyy2G8knuFuH7lLOrwz4bF0xYpFh8K3Vm93SHnGpg5xu
qINYxAT3tKz66/uQHfVKhgpfLqnJ8JFEHp4Vp2AhUSGIz7296v3MI6k2aN0uOF6h
DdggaCkqGfTjEP+VXgYPYkJdhXx7R9IBb44Vt8PkHrp610f0bKZZnkJKDNudgYbY
Ui1jnBsGahE7e3UP71BXyjPRZNwENoo8+ilM18qoXYOjk8tpqaZC0bJfX8JtItZw
LXfskIbr1P87CoHB9zjpkM9Oi/SLE+JrxvspQjJ0yOWKGQhUaVKnqv/7Me3zkQXS
9hITjG5CTfMo6wfEK3y9yoosmIx2RoP76S2d78G0tFWboRZOR3Vz+Jkqb/3YTLRv
xfhtI6//RXTW9yBd0Rf1/+HAusglKznKwOfSIzzzh/SSZyZv1cl/Daz58zRKLvw/
9AnViSjptUfD/a8H2vgFEfyGpy1wOmrwROjPKGeOr+eVkchKfGlWbQfb+9gykQXI
t50+S30h+NLEwWgNYuPP/jKLTQotzkY54QJ7HqOfvv4suNurvQg3NQGlgUpdn9G7
v2RpNiSD5w0DTO4rRC0O//0rpXueyU0uQ1q1MaQubwYeaQTlaqxw+PEGywWpq7GP
wlbo6rXZBPSnjEnz+3JoMxqZNRrBWlnbrf/eZukAENnEtyybx2XciQsFBLKSj64j
768d5BF+JNwBtfoss6PcQ5+8AMsE7IjQY9lzAjUc1E1/6BsB+6U7uXIFyej8h2CP
RQJveJCVFg7yVRzJx8JyIexXb58xVzhgDw3xjU4xaxmW1dlrB2r+/3uycjsjmoS8
KXuWm07k7BzUAyP2RvFnhwGWZwPudKwFNC8v7YWa8DJ1A85L4aTK0zW0JExsuO86
7ITRF4qmSVqh0mEJSkrD20qOVyNyo0uISMBC4wkuPGY3zJJxOxRNQUb3dAXiqMhn
rJeykkPHfnyEgk/It09TSwZIxXsRbccIR+KLKfaoNpSGelt4Y0XyJJ4JrvBV0Jir
VrA/3oLyexNAAHJWSDsKNc2oG93O47VTf8MLpkgGpmrdZ8BaFnnVAZQgYECYRQ0c
yDg2M4OrxSdipVu2KMhhgV2VHuRTBHNHDE06JfQKFquXqRJnsuC0ZIUdwXbdXJx7
eNU32AFA9DF7zmD6YlHCvD3y2Sz5uI7zuVJCK9DFRyXBT+/sh0dDSq5E21xSgyt3
pwckYxlXhpUgAQ82xrfCMxe9mJF+KrzDhl5ohM6x4tmNGajx1iQgBFCbPp2mobIt
LvRZByxt54aKwBMttgBb68vi7p5W1x+M3GTu5yzuQ1JwZuVVb5g/dwRwb7+dClFu
VKNojeac/tuDRYDQkXHsoo2QFfqdKx6J+gvTFI5XpK6LYT+H57GqC5UzNptlmX0d
L+WcqM6UOaacYZ1S4pECDqf2cDaqyuLKBrVhM5iZ/nrLQpVlSPkHSNZyyejXwryR
K7CrYlIlXE7zHhuQut4aZ1rk1fQPauA3+8x5cc7/AJkVVmdf1Ad+SMUmngdEodZ5
69l3gCrgydUSsfw3g9DbjKbjR7MhW2Eonotwha7KD82fo1SxJ9lWP7ggZ/9Vdbqj
XYFkSS/ZXFxlgcgKKFxI2RR60A4LZgLreTcao+2MWBYEbxsEh6mELBvSzB6mhKmW
M/Mi8Yh1/7liJUNuBfs2KO5iK+g+eqbEDIzcZ8gHZx/ZML434nhLf3E96C7yO0Ni
q444S/t6AR+aikKuC+CXjc73sBh/zVjg6nscAkWWJfTK7U78sUWM61CtFwtUwCLx
ngajYM6LTb45S1kKSxMEOLzvTYxz5L0wtoEbKw1fRIfRdjbPx/zUzXxs9nVILIa6
LcSR3PYhdBwipG4jVJWxtOgVvtvTfbyS5AVUF43nnp15ooQjCFgkAunEfMGfrwig
f0N8ERuxLmxRvgkO+yxewIG/KKce/6ZdLnd95oba3mtZnep9RUbRwQZWAh0rTmZg
tpJ3+3fFvWOpxbPzSVU3lFg720Z6t/8z6xETimCJjmHY068qQV86aqUaTyrkBk/4
BdfVMjRm+SqANGY+UaZd+UptJzkL9YTbbx0ZDEFRk8R8gv2zJhcqeXdhIZQXrsTe
/bn1vI+k5TEcTgjxfxHguRWPXgoGx8x1ed9RngU0I4Ui1jeaDmam70GXJUKgPalG
joFzInBBBZ7K408ATjlO3qRgwEVurPwXYvBX6zUa18J71ZwCAKCYrwog5fl3XhiF
IVSiLJCWTpYBg4gr9unZUqr8bvfo4UFT0aEU1xVnxwsXxvse2ftcmjXdmcPEPNZt
8AEMln+XQZme9dLfn7UtQP/6paxHM3IhGlYFgoB3CXShY44KCv9Xtnz9NY4Auwmn
P5hlwpi6eznxhIDb6WyXAz5Ar1sT94u5gx4+cQhKf3Ug7mqCkB9TakQkMWp068BK
MqWWN/OlupH1QHeUuL9UQH+WQUIRECiU94sZL3UsTlpXnBRWMhYcOQsdIS5z21VV
EEuvemrhAcb7ldyyZySJsavpRj4fZvNngDKeDrFuULL1WuG6WWpB3FVoLOcUfQf+
5zt3sY00Q+zfnXqKIsMzKMomArRdwlKhr6bR7b+3krsIdUX8fSC0CDC86Y2BOeWB
blyPJ9L4/zv7I4prcGYHkjcxfvI2WDsoOuPurKyAlN1FeAKMUREA0Lx0ERS1omom
Ls8g9ac1heGS9kKD+cBVF0UYulxpsuTW+zoPdpqbj9gYDhb7oWSE1YHgMG8vCYm3
kikIexeMR0oWqlToQSvqI9scoe1TDGvIU+IfPvXH3JTN9Kjf1EC3I5sGeRfrL0+v
/mDZ/Gm8pauFqQ9cBl6JXzTnPCxhXGDBbTxp61CoQjR2EAjd2Y0Qlrt6lvQcIDlp
LUmfIwoECpX9L907ipr86zdPqlUQW9Dnb2mcCOpa33aJZIuhNWS7mtumJxzbbaeu
AtEr0FIGRsPo2HxQbGkeVgOfLH3Z1D6sAACp3RCz0QKfS5HfAl4akR5xDx1lBq3h
n4z84VwM3bfruwGbRX3KaWVma03ay+M8uVtp0xLiUZJhg6xkAfBNXE52nv7PrEHJ
ScLOwXy86dhY0C3hjgdM85sWdUPObVIvcyfNRRT8zcB7jJ6wQz41t9AEqXs0vltN
DblyYR4ayt6gZWMGOU70oaYwB1I2KgTkeytn66g6SiXR1hDLiYpVkpfVxoQNP9fj
5BoPqM7pTigITdCnrq0dF7YrFWayi0ATiX5kdlUE5xM/OF1307F9dHtKoU/W80F3
q01jcGqq+aFjCtuSBuuRen2A4ZuZL7VCApgr8uBEe+6Flw0PDc7Vt0cmTcsiio0Y
X3tmxUpYfrETriR9t7VxeJ3CKPkFU/AxtpFZNTwUoryFA6CYpnhCnim2xmLkXpop
egLBZa4SQzEFuOqEFtDZJbo0f+CCNaiu1OfljY+OUnaXNjkwywlMdR1I3lIzBHW4
4RLtA/CjiyMgWCNkqGxxyAMTBPsdPxPZYCxYI/NvGYiFQxG7Ygo/4+JIduDr8ljr
HvBZdrmwLL+kck8AI4+eJ4mS+9ekaaCq4guywy3TKR3M2gJ4Z40dujAWVXhDsR9L
ZqGPeKRnqyDDrTjRgfuSGNe35ckt2mlccli/v1SI4ff4IFppzr8JpEQ64zcZGrT9
w315oadwfdYTiCeFbl62ojsl6Kkll42IlEd+E10wP4G9iZ4VRqPK1sH9pqe9XDRA
+zjz90JPEXvOwRzXOyb5WDo7kuOTS/C1o7EW7DPUTy2NU41QfWLTGmeMXLRw3z5V
KJydDaqpnd3ftFyFTaTzPnTu0vUjOowynyAFis6Wyt3QOEky0b1F80bFXEqF/2il
UoeCBQG/WPB9558mMjWTSnVt1x+MrKxkuu/dqiEQBiajY3/MAqFGcfuobw3isVIG
tq92+NAuujCVpuv+93oZoNGgxviyZqcAL1Ly60buMoMwmg8P+jbt9kJ+ozD+xjBP
Oxab8y3VxYI4wwu3Dhx/fOh0f5dj/Agyy+gdXMvw08oWyzPNdeyyMKtClFKGpMHF
VAYkcNa9YGlBX1hR0YyzkRx9NBOBk5oCqS1Knskh47snBPbOCmT4/taKWPlEYyxU
npo79+lgUyC+aToW12gma+HKGQ2aO5URmsQxaUMy9G6Wh+Q7IkxQHCXcFT+P2gma
L01//Tpqhp3EUR5MDyHRpIMAsrKcLUKOSwhrO595O8bO4erIPHjuyDzC0UTVMyrW
GjG0P98VDIOfam8GTrUXjZsAojLWz+dFE0iLh/Ivj43vLX62aNZZa1Y5ANXaF1SV
J+M2fwGkBhEEl/WOq5bumlsqilgMuQNqXmRbBz0tcHdgDynZrlpx46+DAS52wJFf
nZR2bNTVGPXHON10TXMPXiOmUesUPvTkudGrxEmPbPjClNjgzYVbsoxnlpOgCY0i
16FR+vAg1JUbCk4VqP7Xw5FJtvPOkshZDGAh3gtQkoadsnQI429bPh6Hye+rnD4V
Qsfx8J4KeE7Qzqh+ZzjhFcqondWTLp1AuuBhdKWsAdQit+CmrY4CbalkYvjoOwC+
s4tWv+VuFmGGEanzBEP6diqTUya6EaizO+db7jTCewhhSUabVpS1Jdl98W5qDcbK
waHGxmOGPxoQMFl06+VdNm8bKsUr+65oEa7XMnxRLEwdezFq4PDiyA+eQDx/hxVk
wJ3s0ZbsIMHJTsup9f/lPJT5Ku8YFLt9EMCRfQHllbeJZad/NS5d2bBFs8P+YQwZ
E7V6PjIvXwHFNV39kNfryHCUadKDlBupYGdHubIV+1BvoW3+e8iaRd1uNZDVcX1I
GBkjD52JxKVFqMWms+Vdr2zewMRRW7yi6RRMpoIQkP/18G78Z+6K3dWTwuVO6Lnx
lgGjl3FN9Abdy8fvri27eLYQyAiz2/ZG6JxeWU7KkFvEk4eCjWqIJo9Rap8RkVPV
uIcm1z6Wt2ODrJQL2rKu0RcEmrOh23VT6vFu6ZGAZFj/w5cFDh1Ew9TaCCuip7YL
BZQRkht02Yrw0RgAzyEVAZlXobIuMZlXE31QpfcRB7h9tCknVCskl+rTO7TiA7e0
VrmB6E8bW3DSGc4M52IPgcgaXdNn9SLcBV4yzz+Fv88okJ7B6FMQUp5Yhcfcq2t+
5qNO0kXWgNDlHXkCIaYNQQ77HJ4xrMg3cUdJk/12D+e0nl4cjERZte9iI5b1Lj5y
CcVKgtE4HQ/KJ/oCZ5I+39x1ACdPZ/lj+F9Z9iObYvEgmpjTMZhIC31ndE+j10uN
8wfXChd0ZX1p8Af/cDGelXIKHxlWtdpDNwrGPDmna0hyPmlRylCALv61vL64Jl5h
BW+mTh+QCczOG5p5Rqov0f7wBMpTbnGCyCge/IV0XhUsGlFDLu88SH6uXVM4f0XT
pybhbYxnJFTx3LXZuXIG10UmNdtWCAfsgHuZmzZ49FgODUAnVXYe8ZHFrMicaWv2
n7kHJhAoHb34aVWgBmXSENMmzhpu/G9cbIyLfFqSNJjcoocNwAPrHpaqzEw4nhqW
RX8ZpdODGtwhMzpDUreROfj8SxInDRE9qtK9N/nuyDTAKGyQ3JVBmB1+l9MUlp6z
rjl0Nb+WdgtwcFLUA7gUoeM8cv0mugBiLzs9lgUwZRAYJosPsbNndYL2ySKGCTUr
6N0L6gjaZuRAKYANlwOT7Ydek7d9QXVPwqbnjZ/zHXyI7qMSEV7CwUi88/bmMGm0
zoIJ84/e+oaHh6s3+UJN88jEUVMVZ8BVLLR/r5iFeb9LAvEZ3xUXxqoU9I+Gq9LN
0lclKBFT7bohVpDUVfRp3W1uIb2sNDh/9Gs+le9h9h08zvnoJzt51wddmf6Bh/e9
qmsYsBdrB1rozcoIdzUmwfgmvi6S52taKxVcgKNVOzyjCAltBcvYPgk8qI4VMR+2
lOGfwL5apCraQXt6esXdUZpN1RB1H5H1E801BLwCqJixuq1GZiZwuw1ikrc0aLIs
MKsO97NSVlFz06WjxKdJ0/myZuCTNW4PCXflSpOfc08Wi7FvO/fKHDQ6ZhhsuM8L
6aXbuFTlvCWspYgkLR6MZaQ5QfSjqQNIggqDkfnS2IPEoWdPKv9h84CUWRRZR86c
GlSNQEaQtyGlEBa/hMoLI21xuVPH4SOd7REdoppKyuiLB9/K8XN7/iJGPMECkVhZ
pD+F9UqdCv4Qv30rmtACh3mnNRhN4J82HuzKz2CbwwDEm4JjsUKSeEFvzj6WafbE
4hYXH9xQiRCHTgbsgZ+lT3VRPL+G/Q4a1k4HZkg15Y72TvtbxjjmY0hPyGxst6Bo
8ge0RycOrkGYYGNMza8mUeKGPoqxpqnVAQbSO+Fja17pcdGQKSHx5u3C7fPG7Se1
uSjKopGsP0K1cMv40K6MW33AcKtgpKb+9QuMidDETEfktd0X26P/gi2XyEPWakt0
4X/Sd10Pl/Mgec7cD1MYyVh0YjaEyfCtoaavcIG33p5svyxo+I11ggmcagjhcVdZ
ssCwWwejHgAfyxhXcFlLk2sMB7zPHf1plJM3Totj2XaxmKOJ0sZQFaL5/+NCF8U/
HB+s+J8Kca7ZN9+LOwvftLIdV+Yz/1eU626YIyishcneXaKf3NqSbWMe5sLEcXZH
JkAGp+Xyr9ScjO5x+edleJBwljBuJCIEkOHSZ3LEZ94PTb7SCPIsUWYRFawbR6gU
joxsnsElhsEtpQBgmT956DwZu3CsCF+xwG6yjRKQNxxdALC8NVNiy7p2w/0vYPRZ
0Dx6U5qIzd5Uy2JFPttdHvTVIqUBxkR+ZrImJHQ+En7Bit+oHn9Ylidb9YHi/gyg
n23kQiVgHd9cG+fqzVtwW255coT1Q/d72kH2Ce/bA7eK2KvYyAzHB7xk7fCpR3FQ
6z8o1bKQ6cIQzOl6dyY86pTXQHzc78usH8BB32n33dR/P0P3zcOU7RibSrqallrE
2aNf9oIrJvYtYYf2SL+EsGLR6zAct6UICSb4cVIY5HJUR3i1jtqVcNfh9z747wfh
6KRCX6k3rmeLMaO6Y//HRK1yz/zs/mv6+khnntc21mnWm0aIaSoJ+jEAaL5JWJu0
K6B2YPU8YNeJ6D99EyHvSjquwBvBYRPiMer7DR/WMMay6wMW2u7e/Z/yshP7el2X
6o9W/dD8nGUNNH5jmI8YxQtwuaF5d+omLZDdnmBM6P/qF54+rUIP3zTIKO0+T7gL
yxCapY9Y8WHH5KbmyVytCZ834ZT/StOh/aJJANuTTvLPogTGrqrorJAnogwTeKOs
L6VSbExb05fy1nf/YPIQ+wP94vVPSK25xN1t5xzdtQjE7zJkO+jaNU6WC2rf/0iH
q9ZDSZGyv5Jut0J5WV7j+/ledhmQKhmJ3FMEN44GUi4K/bkYNSLYCMLqjaikpby/
96Zm1wRFqQKbkD+fxOCTm5EYR2QRNUMhVEeHUcxKDGgGMcAGdRJFnkzJj+pY8ihn
vmxJsKaAHS5arrQ1pk3AYXuI7zsgTFrsHhdackq8vcssJtI3QMzHPArl4AFpjcqX
JrE52+JMq+hTp0wCyPyTCxIi34c3+FAvBgM59Mfa/VwR/mGBxQUJfFzQzt63nzYo
QtxNY2RerrdjCruGSykb2jpgeKRGq/HaZNU9Qw1jguoepyT77Myqo8q4Fturj994
YEsSgg2kDdVpP1HaLdi1AJpp+XblmxQDHFQhQpVYNIG5nm9ZWH1hwaisWSRCDVgX
aqVxsfkS7BEtMvfSI3v02loF1fTFjI+x4AZxNX2KrLzhJ9gM1pBHkyJkFOpqlOtu
Y2YK+brQMswBCA7eKzygRFgY4/wocrWrX5VXGqmsHoRDHTEAS9GZyKpmy0h2QCNy
Ci3gpYvJWg19a1NKC+ALUkR7Ds0nUZGBtfXZTQDfJcTH227HW6o5OAhZH+tCcAZA
mB1Ride5xQCqzAJPSLzZsGUueaess/FEWMA+1fAII3C2QcGMhcXJNPDuqD5NKWXB
hDzQiHnxhacEYJcjz1NjrAaZd3w8iuM6g7oHvfYtsxaHGKqm6UamCSyatYO+Jr3P
rXFb4cbnwDjkayG34gAuzJLEApDn0cVrMvf9f+0FZfZrjdEoknnqY9vbhawwBmgQ
km147jhE5QuQAc0Vp5+nWyCfJJtn5bRvzdPNTuxFbqft+sKh5OKeTR+mWph3aTCq
o7kuEXqwbbc8kAYUpBX1ALyHayUeIXxWRAHfrwvrLDnG2FsGxQtgrUfAVT28hVSn
rOpjRE8/2c94LD/lamHaHsXU1wh8zd6CvSViYf5WQgvwOcLoFu1cD+KWb9W0gHsO
sGrdnIqv2ZGFJswxx2gWaNy1rf9oNV09pVxfapp+sGXc5j/NKcUC5zz6rKGcIzqf
j3sshFxore8j+VBzXoAAb7iZI+VF/HWXmsdx7QlLlkBftoNHfUDW8UtB1KSEjUgN
gjDr+X6y5FXYAGxkpP5kq8dmE18noBokEuGwubv/g6K9PdViXADHppHZXf0InQAF
Ld1fkU6Pl5YpHjdPwctLfaJkem74HaDeVKEpV7+q9Em1yRgkOuCL3cTsuIU/G9pv
ws6rqn90Nzg7lsJGade663afr/u2VrVjnkuNf5oow+2c/xKfkqSSKnYOqQyUqbzo
44ndfpUuN8GU8DCBWkucUO8BxRq9hvg7gKfUg8p5eGNf3LTP3q9mVGu8cOaT5pYP
2zdI2GcRZ8OvpSfj6IZSIB9KaOdBvM6xo5VjBGu/hA6Z7GvZCCfW87AGl9b3BxXx
oLXfZ3fHrOhX1qfEnbRBWE7iltcACct8h6+4/bPWgtpjDZ6YYC1mEq01SmsoyUtU
88QxXyCpcp5aoOWWhmdRpB4iqCaWhuRAQesXS5YaSBdmrTk2ekG37SBN1Md2Xdzf
ES/2BZ6PdBWsIOIeMrjBu4jBS6FmcrY9CeRoqZ+WDVV55AByfwzPtirQOrYDDdiw
HVWk7dUKF14S1bLS21/vS9gVisxOnzozydBs0kHPDdalESfDGH2Xgamsi4IjCOaK
GD0qntHzT95qOAakmfcD32oINx7o6KMdI8QZ2kfvmDqSsfK2SOlCUpei9kx1pE+u
jop/WfEEfdmuuZA3I8Kjc1m7G1R1mBflUVnNuT90csEHh8w9W6eUiqerJWT1SDyb
heUxPiz7iYB+0xMs4+dDkOz1+7k+Uh4BRrFwn02qftmBN30fJLJeR1/bq5bVfYxa
9CoLbNaEkIfaVXJO43gajxaa9IuTaFPaYnxFogzPEPx8zoThWs+o1/7L8HH3+O0R
RfSE0aS6pbHPhVM+/BzTykHrnMeT2qpA4Xxf5WAKht3vXVdCBLjzoGJno+ys6zHO
k1lF852UIxW67ejJh5QiK9N0+e1Xti5GfjEmXbn2Y1k6zPEpDpO/PognOADVzsb8
7UV6ikgnQVZ8Zd5/4N4BvoANZZ5t+7vMz4pgJnaDA2T+pXNm72+L0G4h2LOsK4Ct
x3uEOvHqnMOukXltc74eRdqQBqwB1CZ4IUutlY4/2dgXjKC3CHlls042R9600TQ1
7qWgfxuoDhMOLwdF3VjYHiMHOX5R10qotUtfeyD0yuJinVaUnkkX7FF1WZNCM/WV
54R1e+XEMSjA78aSLfpNb4S1oSkcLFRGBCVI3VCSrd4PJzSBXGeOj9ciO3kgHV8m
RHWwNxAFamzxMo/zGnFyNvdgZk99P/iYtVnQ4OP13QErA7KqZRHwFez16wXcsH3a
5JiUrapmH0jwOwS+27YK0hGjVmq0OBzfKqIBBBM918zT8J42vGiI3xeFPGwFP8b2
7Ibm6NbTrL04PgFYgY/1mp0Hi1SG/MIyjP0/xyFuW8FTMMJ8Ek0br1CNYhnbCRHz
Q09SEGHwPLjJ7zrq22/9Hiu5PAMSMuihVXI1E+wOUf5e97c47I6itYxo0TsEdyoS
DKgS6ZuIwHKKZhphkY5sO4MeTmEnsTJhQQq6ZXQVTZ07436yKJ0GLK6cwQaRN8cU
gV/aqm91kHJ78zHe0uUH7caYVRNLv7R5+bnbylZzmltQeQRKX1HWmz9uU8g1t9y5
67RoePN50SIi0/qwmlt9KsSAJ2qHtK+rAutPhYS+WSAsEOYOZl7FMf+j1Gi5l+GL
Gs0o569mK07GbI6zEvlT2cBlHunRXhlx8sSowzPyIYWAgCYDEg5DJhdtlONOyzV1
YBoqOmIjpGu736MsDNvxz56gqcv5bLuztxwrmImS6IwfjAo6fQ/AJhNPQNtuqX+V
bOkDjVGryPDD1E21kCI2q8WrE/GzdXdwkjJ1V3n/ytXXsLz6P67dJR4tbBQ60kSY
HINMe+UbaDHh888AC3JKf3vDm9mA6BsRblpax7sy/wzHEIz8HZSaq/asFkfphCe+
AuSDi94ptc5sfwep/RNyrE3059qdQeNxfwdOSbeAigSqm9O7C1dBsgXiKSJQwdNT
xRelalY7RLNFEDL6L0yW+qmbeaU6M6vxKlDxfFkLTTIzWkbOwUorzmgZHpKLyUux
DtiqGwO7j/OqlYrAAvMhdAVpUvv96KsDVzV/Wy2lq+TXMsCzN844rDaXdKPLnfhp
Q42hlnxyMS69NOrdGF6rkX0pQkolmm2yGgCR72r8Z8k4ubChcl7vEItgTg467hGN
sZqBt95i0kA0Go7xZqfKRQQrOYL6a1NS/AsJcNAH23zfni/35QsXV/sZ5O1hvYes
/ur4Vk1s0r/GW8G9APuXMe7wPm38qPrBOHNW3Se1hBQEXjphpZ5MTtgHJYbpDU7z
iyoRDv9/7GiKqovDw47mwY66O296sPzM3NQEHgF3z4BPm4YjNizc5RKhuZYAt+21
4EihgLaQqikRLLFCA1KAjWpGy/BtCT0wzkUg88rdwhwgYshw8MZfYHfQ3NErbUJu
DBkexngmI8BNThECQiBAMt8YhYY3tH1veJq2hPc9XiJdze3WrUAYDUdGa/zqzFoR
HG+hOpP+siyWjgO4lBQf6xzcKQxnWwM2cp2cxvY6JVGvXtAKPEVOLth0idbSp7MI
V4fyLm/gNH1pXBlpSLyka/tH30sU/pb63xBL1MkvLpxb5E2dPWGjIh+NIOpmE5DP
6VcRyZXYV3t0FjI+Y3ysb/z6/eaSgYL5z1ogysrPSFKCMUogefalUSE0JsPp3q8G
um6HYYbyz/XuK++CFNjqwTO5XND21nc9WzYgaxzjy2jPffjw69X2RuAwwKcRHCeK
0L7Agr1VUtf2FyMuXaKMtWAqU+VulXz1Xq2tUwj1johRVFr/k+IrQHQf87DP1r47
p4ZUKYYfvKcwtdgeDXhDIlxjPEID8zxm1CuuPqS6oUnT9cQ1rAtDCls5nfkdpHW5
7pKykKRuU/XCZi8Ihua25lF9xNfq5wEhrw+GCEVh28m8HSFXcEGuaQWLvJa0rXxb
+TZ1IPaoHlSUJjfeAHrIpQLJOwjVCcpbAUnEAKztmZFkCWYYtcdgDJXF89c8dI5o
1VOdNr1OEg+9TIPh+/1BG/zbzFeIvfJRZgMfR5F3Y98MZDe3iHWiFn5YOq0H28hk
AueyvIYdkS3x4/yZ8Goe+zlVYmYiIGemyYBPE+L4fwnvu3GGM0kKbioCQANyrf5u
/bQt/1amg1Gwt14hyKpplpyFIKLxU5E2AsGhJzPMhS9BJXfinBQ8Z5JBU51jOQjz
Z5o+ZGcnRLCNtLr7F9C2HP8W5EZ1yDFRQJfYZCq7uX/TKhQTx90U7qn8vw963kv2
4OF3xR10i3Q/kRg0vCBlnfuTmNh3WK0m8IjJGcAlTgr1cCjg+UmV8CPGQpXhtjn2
GkBrwBi6cRiK0WrBOpPdHj7HRspP06D29qSfYKV38tG/ywJpp0nXdseHwWFFQWem
aM0EV9OeLeYEY2ig6BRigRX0RRWLVWYPsGHihg6QsC2Jsrs3fERq8lZ8goOn40pQ
JLleGHCphfLACkIQcniX9aW9rD+FWjgSHosamsnbYAZCWmCiEg2CeCKHwkrP8zMI
FmAFSWy9w1N6M3AR68hXLhsP1YH7r/mrqnBpFyy6SUOU4jR/UEdRefICDmdjrW8J
XD9iZPdGQKCAD5Xw9ablol6kXiv3GUa3mD6zAerIJ+mSlIryLKUOdCokth4gJJty
ZS9BA3ZdxJe0Otpd0Gz6MFBoJzHDzAd0TtICbJUqLuR1SM3e00gThWGLPQmkzRGB
d1y6WhkpGBBQh5q+sk+zXCusWsclFQvjO9lxi3GEcTHnGHQiiWbFQKjEqOl7gHnl
0Z1UQEztME43vtRrgLwKH1aaPkdVUfgeSuDsa2oPxAixKJKVSh4MzVpKaVe9NhRI
504DRb0/+UH/xbXEgQn8+af3J6YQ9H5QB8lo35hA80DWOM32JyHkNCwjIafrd8Vb
FfaFiJ7trRMzU02SajYJEm3h2P46Gm3yuZeMLZnVcqmnpFcSwfkdNlLbbz/x2W4q
7sGDX0li8HrYsn5NO1x/nTi5Y65p2p2eCyaPbd3H0y3dtoxITqdQm3sdRQdgYH0D
R/003LRCZnA5cyxGYw1vY1x9pG92hV28OvCZg51LgP4f/QzXzWIQ6fkWRcnkaH+L
yotNLDkBSsQ+oB4Mt5S5MsxecpQBzYIru8QqJyHulCNi7uqCEhMXxyIx1ZB24ttc
VFJ/kNe+MQOIak2vtLW3r93HMv/AWx+snd6Ep+WaAIiCApjhe6ZejBmUFUqevPOv
IMyMjyauNhbmYTcmeUc3k+f8Vz6vgXn3mOGy9yW3eRRSAJTZCD5Xyj+r8oKWKlcO
DBplfmBPtG2iRx1DGHHUbsusuZyV1cNc4jX0l4zdo4iHnNsZl6BDWdkSM7B2uLA/
LE7J9HCcPm6ZH2LRoNaLgY3+HHPkdHa9MYQBHw1gCVMJNi8ITaeuztktkPMt2dQy
go//Xkv8rrbWUcRBC+HH9mUuYz7zi0PlOtGlpWa9ytgHq3nMpLWC/HaIjoz8tnsq
RWyrdzJwh0ZQm8jvswpIip3npDRSY618WtV9Vga6AiFRdYe/x4jLk3wZIIuCCA97
6k2p+KqRJZ3cbLRrMEqo7YTq817pgpH3J+HqnrMmQb416j2nJZS3TDqa/MaKiOBT
J38MCptcnocMmZ58Ktjqgh2E6OcLreLnj+CDfOi7l5hEVHmksD0CPIC0Ce6RJ/fN
RqY/YVNgK70DDK3JG2vUmxyPQkUtmMfWG9P77nP8FXZDXGhvsAkExXgNf1oE69JE
GrDC4Wd/d0FOAuOaMnTm7ySI2cVTJgf1RmfjsbqqMLDzCi5kwC7vYc+LAJV2T+I4
/TGCgNjie1KzlvKEpTFWJpZbz7zllrEEKstXMI8myU0P1gCiOoV3aL0a1Wwoq4C0
C6lbrXUt09Q+H6QgAzAbalUsYjeBwj9cLPPCyhbJGa2cRwvxsn+8Hbcb+nGCVt66
6Sje+sm17aKhxSdBswcPxVIZWUEmjTrK3fmzG40TTUylFoIUYdMscePKB95P9BXo
fALkErLwyPRTGvL41CkW7/YWVOsdeq1EaclkFpNzWoqTmE2DgPBi9/ChyAKoS45f
yVpPAdszyG/2S8eUDO490NMGFrT636GdmM6kuNJQTM9f0oXi8S19FZdcbzuUe1n+
/I7YdvHW2gGHervlHXhu4XxH+Yap19GsZhiFBAqO+IffAVT5PFr+VAZbeAytEK7+
ClW3YR4sZhUzfzTmYdx75vhkdqz2hcw3DyRr2RyRhyuq7sYeLDFUlVGE/Q3NMLn5
J5E7aUe66fD6PNmoqXL/x5x7JUvuWwhjHwBnsdUpSP1k1hXlSx3P2IY1Q/GrzhiQ
EQAihlpI0/2BcmjaNNcLtqtwplwXQCaZBLdV59LX0+kpdDvWf4GbUlXNZlI8TIlM
OEfIX2Jz324muLh66se8Iv1NuILaBBuC+QIpco/LUeS0+SmfWFFZPDyN+ZdMP+Kp
63G2iSOzTJ63/N1NELGbnyDNVGZ3Li7gC/ul5Kz8ciA8QFPtWdcPDFSTFDPlLnks
6xYj/g9wIQPB1Kdcbiire5MmI3RHaergDzW6Ym9S+76FLnOHtPi8clJwEeQV/9NQ
0p3FqE+TIgL50oP6dcoAIuRtnpzRCrP52HxZUGy+LY+9ZK9HbK6kzGIjwO+Q4yES
4vDMJqA1AopQmZs3zzjFD8XjTzHLRCzzak4dM+jyAGDwSC4tihVVtgbAqI2RinFy
6eg8RVNCONTIt0XbxbXQGjd2BmxQ87qmWuxQbDvKzvV4ic59oSKS5ndAUjkDH/nY
9KJ6c8adbFlj+hgdZz77+eOPwjq6F3b9/QfdFkMux0w6GQ5uPNrq6YfXeRT69ema
PPjpsmbzQH3lL0DsDhU0oufLq2lNmQBQb1orcDEYProDBRsxnm2UZ22YMnjGCJL5
dpDq+V8k+2KPpBy0ifeCSRqUdl231Qx9+pnpwRe5lhKk2BxZcy/apfHybYbMenT0
4WTiJhFuqucru/refUBphmTscH2C9a8Rsy/+dlh6R4YwCQvwagPCNXtpmzGmtz7H
eclnYUiB/gnCo3iMXhttyH4uPnZMzTpScRKTApHIxw+iFLc96LGX5dPVOP0SIkvr
5cKe2pUVUH7vaWOBi0j4103DU09Y1qJxZd6h5TPDe/bht/+vQUn47v/byWP3sAGC
Hm+WEgN0qhF9CfrsqcibwJox59aSAqTO5KzDICEW2LqbZSHVCUIqaub3Fd6ZEFcZ
5FXeuIGrAHgN1SdxcH1Apfx1FtTX29U4Ko0egtsX5ovUWbJTnsNEqFeC4s99FFw5
Qm+b6a2PmsCw5UjN0qR4Y0GFfPNt/bkLabDs+qwEgh9jq5ZRABkqN1ZeGZp4e9Jn
pifyZQK+WsgPVt3DYKrQmmSXkcNHwh2ZniULwRA0gCLqap+pwLx24efXs6yTlPJ7
F6WDhn06YP/3Of+WbMX/j70sRoOp1uG+Eg/TAfXJZ3ISxt/qa4KGi2Jem6mNOaJG
cGTiylxqSSCy0WmpDQ4rOCDAgT6ZZbhGl7NXvcS4rY0+1VbaAde+/GtxnLHK/248
HbW7BVmbDj6NJCAdltDB90niTZY48LEZQr24tSS/Kbx6A5YWljL8zMvtrlRvtOHB
GrXKr2UmmJdOaBpU8WHdYdv5FN4g1VU2/89r0IyjaCF0UWjHJ6fb0cKo9l0qiVez
92u5RgGll85JK8fyE996E6Y5KOFnaf9aRkRy5ozGSEfr4aYHZijylUee47VlkX6O
+h5rR/D4acFpo+TWDEnosZ4aURdkHnl8eWscgm4gwMYTbydOyIp3Seslmob9Z5Kp
3Bnyiwr6SnqEXqft5BT/Ng6En2DSg5yvN4ZaiibEYIHvsSB0ebHv09Y8ed5BE10n
BOZxofz8t+wz1ZrYrFs2SOFK+SMjP7OmSgH1oW7aH1y0S1duW7MaAOXn9riCLje3
qNBtkbVjdO8fKgpwBCjEOQ/22UYYJRk9mWYpfjpV92QoE9Tw+yw+o+fsjOmUh2D2
ugYGumUEgnoZ55Eafj6vh1AFxi5oHMdCmxukqw5T4WEegPPNoTamk1bMsundyA/1
hiF5pqdfY3LjSITzto6jzqMXs9JX4m4OeGYDnAT27N2yfSEsD+IrPtk+sgR2WXpb
3dVh/38IDmhLRRO/kk2BrSjC7Dj+atzVP//xEsbBRd9KkopjhYISW+UjcHlfrme1
KOXIftpPrwmlTNufwBCKJoOQ43lyXujiZYl7opgAQK75YVnqHwpq105SvkwomyVd
iJ6Og2cX67qfHyvMxlpElBJI8GcmPCvWVErw1CeJrK4letCwSa7WCx+S6UIjss4s
4JN23QN9Eij/8xWQQ22PwDJWT7DC+hiFXj5buVElE9SqHjVIKll4ulUCnNIXnIk0
UJAdEUyk/F4SeEjNuPGVT+/4AB2dYE/EGz/FwqAXw/c2PyWSgn0CxzK0Cfbqw86t
f8DueFHXhfjMKKDrbClJ0k9TcQanNA4k7KizuDANdhE3PFQwjcalEB3ukRK0+r98
rkaXIF/i5F1FUkBX7ZogGJuvXS1ESOlOiFKcvN5XsOvmVPrcRC6OLP2qVF/gxr33
51y93rzHg2Qn/puUnE5DkyYqty2SBy03VNW+VYkQ3UQe0oZuar/lrC96EHqSHql9
sEF3SRIIsDchC2NDGdxztJEOKPoMWaJhkxWHi2WEzw1AE88xX0mv+u32PCnPKpo/
c6v41+DW8QovcWa6gXLhvo5plFcnAZcrnN0w1UOpZZ9SY2KVZtOvcjm9t3uJE/8Z
l831E0pc08waRn8sQjLuvXtOYRCBEUqyyvMXjDKjC7HqgqA/cwqJAygFUL/8QrWv
sYPS+490hKgLaE199qVAw1SBSYYinkPVymg0xe/PZaY4c8gT1AY9NBnlkbvSWTKQ
ZXGKLmT1PWOMjQxAyEpRLQE22M+dpPEq+Y5lQw2wSrkhFCjn0l9lH/+oPN0K6dvx
fajI/HKdqsdzCOczOs06W9o0jG9u0xK004Lc+CKvlFCr5uY9GmwJDxgu8lPz1uah
equgrCVBPnxON4HAA+ftKRB13V5oeqIwa+B7F1pCgXPXRzoiRoESXn2mskZ/Ccik
DRwHi/W8RiSV63g5IPMjr81HIyJyhW/NVEG11seu9PvOqgQsI2+xFmhlyQnHzz5F
eIYDLL2f2rnoT35NGIMHYdDcohq93C+EoCNDQbjIdE81RjTz7Dw5Bv6jpCY7dloW
9u4XYAvyRjsg5s4EZy+ALwB1vz5f4Bp8TQCGWtm/xGvmS473rk7kxylTzh3G+q/s
2exDOgPD2BigtOWGQkLzpi+N9dXHpaOBmzqxbb7/wwvXkiGe3xmqConlAehSrso3
4gzxhSztVwz0kDTFOdrcMN52zOQZpDu78zrl5psrUUxp3eU05N3wY+n+Ck8r8Qs6
DMSXayKGQBVvvnXByCNI5p8aIHwaHXYmNFClTKy0r2hqmZYiG8v7r+BHBuEKkJ5C
Sr/rn/mlJZwCMrrUg2lFfXS8++7M+jDihhemf1wVc1nIYVVtR7R2tO0jk26RJaQL
pk+gutH5SjjcNzPvymPAimcslA2RDkR4ZtKxGZpxcfylHYeC01lCZX5LAmszKtbM
M4IgiQF2/gD7rr5lauZqcPtKX5I60HBolTHZ9QYfItN7ihfV9oshsb4yJ+Xyyz0p
x2x4RWUVO2tSVSFQduBTJJjZ9us34ORxBXuLtC4j9bUjvw/lJHJLmJWHGEtzUpVF
QiIV//brIMO/iOjzasEacTySRDtdTvOzv7HIlY9GA2LA4sknfQ7WlLwRNF1AYn5E
Jk4WAbgb6mSfdoINv2+JH+KF0ONSG4clSbK5JpjYrmimFZ5+QNZZCJKqhv9v6PCZ
obqycjZ1EGjeJLkhGuOuL3Yo8NzTM9AlIKsjsOjl0HdnI0yhX3cLzE5bmTBlRMrj
m2FelrKnxGzD1P684cohRdTi99FXhoH3UPS/7Yy/CxExucms9mCKmTUW8bphtUVl
dVN3qr2OsQVo3f7I1az1ZTMEUaMRKA6g4gACE5lM+2P/7CvEX0DXBBrXEISRU1CP
Y5VnkLpy1VLTyeFvJXVzv+X1unx/ORks/wpTOneV7SzAf+84XCy5ksvUR5YhSEkN
98fccfrrWRlmlZ5U2XiWIpHwobn03I1RSBGJk2TCVbVS9JsJQNqHGJbYHcJHB+Eq
Mv0Xjat0qRlnZ/VMRZdkkOgB7TfWHp6AyVWb3AZvj0ymAHB+TS2hzMSNcPJSY7m+
u6vUfHxzfxQL3JzbVeulEVX/duBHiRH7dwDfTkUNRsGIMThx3erQUj6hmj2AmYHl
8L80/NsHHshrdHMq3pP8UI/ad78r8aqHz66g3itEiTm5WQv7CzrFLMyyfztCNJL7
yfNeIdZN4ZXwz7sQwKiSZI4fi5g6xRRpLFCsNNDmvwkQTl2NsOfgb65Z1+qwJDQO
GGSt1rTKhnobKjEc458N2u7KHjmU5BbdW9TmqfWBjBMyFkbikcQN64XoYjGcXm/Y
KfRzTRj4ZBPNvZ6GtB+QP9X7jOIeH2WdYmW5O+S15svv7ADEbMukUVkSBp56Ucbj
CklH8dTfpusn6Qvyvmu0tRHzR3ahCHQ8hIPSLKCYfNW3JvZJ8Vkue1C3RZXbqQA3
/cO+JWEiWNpeI8DrTfdTanYeNYcEeL51kVRdXg2UDYQJmUVd4fpyPORXw/fbISqI
MMWEzblnExQFV9T/PZEZK7vKWqr1BwZtYkeE7ljd0QtI3yLXhl6lHJoUoGbV4k3t
ugCaCWnynLGULgBLMZVZsTUuqPVBhjp+0Dt2DHJLHCOpjjn3SXateiBksxs/NL+N
unvQgllnrTgLp+k1KHDyGh5h2WQUY730Y5iFfDmyTOM/ZMQ7sP2hD3zl1OAEXnS3
iXIsvQ1RWMr4TC00BBxDM209Tg736c/E3WsMcvOoth8wqeZ1kwoXqy/x9VSYU0h9
/pG/x5KIXLRycNCuJk3UORBNCTzr7i9Dc/XQeRm6BUrifZ0LJ35J0WssbBW6V1b3
68XRqJqHhtp8ZHLTBu6Q9ZFYvJugXhwL77TvW0bEi5n3DslK7NLrbqOnlhm0ilrm
dgKs96yGj8TFT3zF31UAOWPx2T6DGmPNTT73BcZDzZXaLJa7zkF6xH9KXIkaqLhf
pzRo5sVbW6wIPpIFIozBrj3pn7M3Db72WC+nMnCcElWD0tXJufMmIWAVP5HAC9UG
2S6wTtqx21hbK/OdVY+OzuMtm440O6MJO3aGqOD6aeOj9ZM22TCwyZ3akvbbJpv4
jmCGBgpD2UnL/Lq+40AV/8T19iu4hnIWghygtsEYgGbrpNRsvgj18SwpI5q3qbzw
WlV8KyiCDOs35+x+dsIx1+vGZbw+yTtJ/CkPLJa7pSL4gf4JGkwERjBE74JHETXq
P4yGMP1Aiewrp+G4pDuGSsCQ2e26Lazl82M+e3kUmcw8CtCmodHLAe5vt9QA8wPW
r6DqoTCfoDhh6Wijlh/SPcMNpMwPpHfbIZXGGanciWcNkeo/R5iowgcrcbGSisGp
EjZQco5upcakSG8CvW0RPiN31T9klCUBwPzfxbbamEY/zqwIa916tq91rFL4gPdT
gu/S8DOncQp/g5ZGdkNZ8vK9DFUKrSrJbfn4NOdt/+NaI5rcqWVAtQ7j98IvNJiu
DbyYj5JJiSkcroMGfh5jFsswR+Gmmp5dWJU86ck8ExIGp5mwn+WD6gyJEX/jh87r
gVGOQg0sJFSiXq7yj5+4S0JKvYASGUN0fW6jaA2ZmcRGAtGq8IENJR523jXFj5ho
nIWm1w+Gzoj3Z1YANriXT5cnOsTeIvvvFoB7WLgryHjvHevajRsxhgGaYm/8sMFx
QNCmrO4xHNdXTHhL8jVNCkcnTpA8HVcWaOXjeKsgnEfJoLVT9hNTKORpJxttjAoj
Ux9WnEMRcvcCSz3KLXUzDhJTxwrQdCoKA53GOlvBi/m9hhMrht60mr0i0XsxqlJB
NSYk98NeYBUhCbqbg1/oU/RHKPxyTS9Jcas6nd/OdfR4YL2IQW9kSuQupCCjGgtt
vDdVJq+NspocdkD+6B6jPG4tYvtobImEHn8T7jiAt2IRTQfhjIP3MtD78DTN3TlT
TIZx8kssX/OKocCtmH9UYkDSG1GXLVOgkolIOiQf3liaoX9Hm95btpxj+BSPaSMs
qNHz1M1wv7/9oI9+9tHUMZ4kQJYJJ6JKxLHn+jBzi6epjlfb33DMw7t6WHDHZOsk
rZJtKuFWZ/lHX1pnLiTLcAKis+gP/AztrhVLocJE9zDXYQWVO6Oo6YXMAeIGnM+9
qnHaoZih7jYz1wzhtorGr/Xw7LUlbt8ZTRxgPRp8z7b/ya9LU7FmkRMoysXM1WFL
RpQ9TngIoBwoEiueMhoKlvggiJMIlxF9+WzkyWk73LkcPZc7YWOrVElAh9YJL0Mb
zP1kkhrkrMcAMadGKL7XVFGNWKcISqNZGtzMkJ82zQIPcdkYkTM5I1V7m+l/y3gG
6YgJZopq+U5Q5QuCUKxjLlXIHDbtAa046jnL+dxng54POgqhLaDUXaLJ6S3E0zcP
F2VqEy9uLNx5UpdE9icZlNIq1Letuk9woh9KArFy6JBZqltorld1Ba1OA0dCeeQQ
TNaIpVD2ZaJFEDWVkZfqB5/iKPlmUGqzsBP1omYmtJZcYSd/3KtoAJD03dOp32kH
4O33EQE1rYJDIEQnZKAb6jXBJ1aOulvf+lbDLl2nO/i4LtBFxcRNMRIYvZb5l/r9
Omm+QdCPPGZsms7LfQQ0cnE3gjA4E0JPogIiJHRcaTKqVDhOxt2bvoPPc87oKe0w
2t0lpSFL4a/lgpvTI2TTQGb4Bo3VESXFYGkeNd0F4qJGx/hQzVFxPqlIeQndQqZN
UFEhqn2Q/E2a0y6swf+V0Etns3jbTsDbI8OIVIqYtf9eK//fhb2ubQAnD1OV5X72
d4oK+aNPyNcNaDo3u8onF+bN9ICYl3wk0AV6MI33yeQO549UQqwX53GcUpslXDkA
WiouqbaoxgXXzFPOmHSgxKXa1bNs/eY4AthlPUuhT7Fx0epdoHhZ38OZcjgPk6aa
h5kv3JGmDhjgEEIxAl4JeGRhMGXL54J0F/Ve3brgm9GrJupdUKMDEa5fHySKH0IN
b1PxYguW7WLtPP3DjyDWY1F7DoIeqiz6rny1134k9d5AAh0inKzqFiaYBan+bUn4
HbmDb2HeetmZitdk8HfpVyvIzp4ISj5HcbxdMcG1enfoQShrmYOrzZod3qnZPrYL
nP+9pQhjSue1E06WbQFJDqB4RBATHB6vD3zIWDBTvGsAdDstPWIRtHUJKmfoS7vh
dhEGRpVT0ireWXKwCcHAsNerGKFtmRS58RI6FWXN04N4Z9VxtcjPhBXm6d3xQt8U
qJK8S4dVc/VzEmDR526z/kTjQ0n3df0IzfG3NtPVav2DKgUEQD6GXf6qBSYeruTE
wc7931mtja0lXlUpgTKJsCaLG3wmG4DaRrda7Mh6j1ZVrQa09dSyvLni9rDjEj0g
NEdnIKSA/QHU9MTy7+o32tQSQVKS1eNsDi0uH6D3kbtc3CGy097jkMLgUhk5QKRs
Sq4AZJjqzAYSoeXI2WAgM19ApjH2yBP/t5afyP6d9qwbaDikF+e7PE+bnF8XcSXG
TdqgI0112vRogGLWdUxWFPqopaIkT6FQAM469l6FfIaIY5h1sn40EjefU+X1Qrat
xCKnruSgbH6TRbTwZdR7rLR83Rh6fm1cLAKUHounBLhkQiUpAECSEE9vKWY4yJSL
yxSAK/nfu5FPIjZCBmCRA9NurgNF0iYj/g2kkTzkQaxSb8F1uT9N1kHD4TFX225G
u/1FpK4F/I/+eRZ6lAAXNMCFm0usTQ6colBzvUp0XEsUgFJXBTF+Gbly4RtxFiWI
GxbLuCup14m5GaznpCeQMJX+g7e4g7yWdoD6jNXn3YPusdZbxTgPp60EOwI1LPB6
m/gcXGoOfD83sr5eTVDcglH2dLvKExJmVnm+tZHiK/bBha+8QAf3q3TyzO4ZzvG1
vZemvsqUotxdVtxvT7uVbGpngdotniV4Jonx9VFXlFiIjCD2PQ8PL4BkAcQZPDHd
aCKMUXIAEFvsGvKDUgzLSCFTBWUAPlil3tUE+9wZiGhU8KMgM/p6MhNl7r9wUvL0
B4a+aSmTqdP/FYAJrAwOh11qO4CaWfallHmKUstBOWRBLqiJi8kbBftahU1krYKI
vIZ7GxfEWt703xsaR8H16sHscFLYZT4nfSMizOQEzbpCBT9g0bA4z4cAWLZt5wd+
d7jMsZT9YKuJOB+D7z7ZbFjw0h83ekfqGYBCWJmlOtiZMzq6EcJyKIe7az1RHjYN
/nlW2EcKHnA9wydutJOd3afAw3F2fB+Wsw41meu0TvcnOLZuSkefssIQnJEu1Hcf
kYWWwNWFLMrIzWMSi12dEcTjqBXUvl8msfpYBubpNJ1YgiQFYhkEG86MMj2N+UXR
1rYj4XwF/9W3vJLb/0lg3AzkDbwpe70QGsoCU2L7794WWikEDDoqMMDj8ToJbQ/1
JUNB+w2bC9URM6AOa0tR1MfwWn/NHgDRVtutCnnpO8nh4ITv+K4ZNgEyW4WHSaor
/casknOPMjFg7cacdJQctlzioAsTfJYlU4lURcSf6PkoDSbBBOqY5dDVWVOZmCjL
RdYbjLvmQCbPUayVkKNDEeJxXy5mKKUcrI8WEw4B9hBrhKcX/9FR7Xu8kMTUQ4zm
cEUVab1tu5qQbotqfn8EeKMRGRxhhDn78q97RyP+v3q+157pM3drvX26hLEEk0CK
JLaiaTtNvl4rsS4KS9AEJScSX/slcOlW8GkVHjgGa8YPMs8IIrUl5++q+1ooIJaB
QtK9g+ZZuekWOyufP972A57BStsbqTUc/ecx/96rcOfGzssjt+Yz57KJYeBI8+po
SGj0vTSVT6Fa8wDhS58+qx8d19ZCzaWmUJdlEqSQPSCZOQJBufRRwPw5Tc1tdMjy
CZlDe8N1UUa0HqFkRGiSMOU+GgdQjPTH57BvUhUcNiTKJa5I4zjvk2NdeeRkJxQ6
tS+18kq3qWQAv6ed3Q6BPwA9vJAUfE5XXFcYpQggO2THvY8RVMf0t3ovvXlcrkoa
3CdgYbInhGZZvXk1hzcHDTciyvDtkvIGXmfDz8otsgTS4ZisD6KolTbCk/kfiJD4
6hBKhb5GEqjkexNaz8xICC2pc5aojyJPyWK+sDFvu4VbrW3li89O3/M8mWBpg/S2
IUtWlaQbhrQMAfRZLcPkHhW8wQd+47GxJK79QDwkj4yt/pvhxbEpcGHFkv2sCsDO
0fr2ytDek9T7IHOahGoemvWk+ZmN93kix2g/fMa9x7P+ncjTEqaRwYXltvs/dBbw
qTmFHbpRtGrOhdxKqg8juEiuNW+R1JDp3DwTcEHfbe0O88c5jSM1nb6SF7dUmzNn
9/GpsYyhoR/ZNbdx9Thd35R4Mk/VtitClv1yM+Eba5Ya+uMQWawP6jhycxo4emL/
ppO0hr4xriu3GKLmXR5tl5bgYJj6+My9XuQSE4WAi5XgOS/GC7tiTF8am7OzSSrc
b+FbH7avyR+pc8q4OLZHL+Z2D83ik2nI1ZiZjnRTip7wPwkMogD+SsGbXqb0NNrj
08xjj9KY5foXY++/IQ1mQM5K90qTERH6uy2g6vOsdJGBZxW/rjU1bCOaE4kmfbHU
y62j4j2noeAe0XyfaNJcQCl8ujhcQgh/sSfklJyX0UIz7BDFe4DfM0wjvF0Yht6A
dcpfusCnwhy/7tYZ7eJl1W/lhWZDBN3pqYrC+qrCx0Ip+wmPk65RU5mg6/udrgod
jusdwEpBISsL7APfRoVgr3WPzAn7urZKbPPJu8mfSRpEeUrlLja+c5/NpStWqC2s
Qx9jg47oqF5bXILM6YzVB0o19UU+LFxXEFpngzDRgat5HoUsu7E/x5/iR2ZoyNIQ
WXNo1mjciXaAT5qDJ9j1HdW+2DNVh9lgXPV5VxasX45DMRwyLHRiFV/dNorIdHMF
iMY5ayCk3M96LhOH+9LyKk1GRALMEk/3NAukIVVxgeINws0AQKWSK+zvstUSglIL
cjmmgVw2l1dDRyXn3gjCkv7HMImqnGc0Ys6y4WqTEDL4S7GVWHAjukShQqCNYHq6
oNyJPctmOnNR/LxeD8VKdqUNZL4S+i59efVKEar8YCY2Kpe/pWHnaG+gK1EK6jJV
S+4ns0HtJfQ8roMGRK/n0Xfg1hjknFnu9QtFuTlh0wm8yABdMxjpKcj6Mk614lE/
hkVCBctiK3WF5EtMDNWVu9UDFBoo/ITp88iwIYq63v9PmfbVJA9DaNZXvLtYKS0R
mJO/b4H4YrrKIZ3bkLuPVZWP1hXdwvFGl55ns9PNaHxdrlngW0ZBuu/RpeoddNrt
5BKwqsy3D8NYhtar2AG61jMw6eceswEkmddd6ubDudTEgYYwBxCHJweoh85Z2qZ0
zSAMcKoxOg+51LdHXj3ovTVMZTOYq2K2HPvaz1NAu1yifELK8HICN6pMT3VIKsVW
Wp/YdzMTvjOZ17eYR8GuXcaMoAMJmsJjMWYR1kGfc0ZvKbgKKnavegxklmoA6Tpv
YW4noG+aoUHCft9fLkfTrtxd0CM+1khjMsGG4yXKQqYyAwl85yTOdyH2+KECZZsz
C4J+mZJcSkDvuLGyy6FYkfmXX5ryijnNBx5DMQaOd5h7JKN1A5gvNzFXomvTMoWG
MYJ3NBsMMIOQ7hhiL0tiHH1bks61dMj7bguTBs5jGHQl/MjtEF0xGeQ4rZ8P5xMO
GDYQRVaehJ6qKRhuwa5t8mdlz7GNA3Sh9eND+4Rhkg/Fp73dLb7QXMvpPWCjfQXi
L6tvXaRJOkRe96Qc9BVcaqa0TZRSelas2NGXJIOkrOHlpYZMsAgGZGUtuNdEmu8S
N6Wb5yhmOkdcWZYCtH4yxAgB6wb+tAPKBDkkdC2+3J4B9bJCuaugGRNmWlhApFar
NZZEOjy7H5Gl9gaPdOEmdQo4WHeFGn/DHOrt58x2VSBsXjrr14+5vgsK7Gz9+ymY
DZDQjNURHBMBcrnobynNZ8WW12N0ROurQLgOXi1hQf9yz2OuzHtEftmjFept2Ncf
fjv1voyGuh4azOTX1EXQw0Ffo/97ZRbHkQlZPHjVz7/0vFv0NQr9K2RXoh6CX7qH
/QMkyoo5TAuG3EGylO7ZSb+pB6pyfUPa5fe6UwOmADiWyPwC9/WB0NXc/3bqn4VL
4359QittbT5AaC3FWO0R5ZG843JTnrnBnYXKE/2nE2rTIHG721Dx3gEDrKtM8J4I
0GefYtUgn+Ali9/GCn6mqMfrqM+kU+9GqJmusVocix+UyfmCB/MfvlTgRmpje65q
sSQDsc9hiSfdSj/lGQeT8rg9aC7AvqMh4vlU8K1fagylwAl7WbKB5DnVL/xGTTv3
1DeFyXcpbBcZjCho8YIcC1Xlx1mFBBBNsKF5CVFA8lyh1B6c2D8fsdPjocJdVxHh
egDNK+tWzSCPcB0zXkK1YuvyER5Oigiq09mSsOe1XM3Ffp6IQJK+967BgMjn7UXR
LbypmvoD022dGV6lGy39CsT9ej5dR3XNc8WOK4gEMoiaKaGJnNOtsnFUAd/NXC6L
ODDwiYS4ZZ//aIkKv6MobWD/GBZ/lEufXjwlpulHhi517j1WHwgeIyaubbE8Jh9e
R0nxGpmJ6vziRLPUYPpqyZWYjRs/XeNmRsj/FLy4I9OVZ0QFF7NfQNJQLlNlIwFA
/Vxn+Qx8jjlTUObVGLyqP+xqEkWczGRcIOxwNy86HsrVjX/Dm854RZtWKqOzmJmx
Bixc4BK0fQXcFI0uQlS44IMZqgIAWM4aop2RWbc3ZJyQC9lfp3EHsWiXRLQKHv26
qoWHsddIz4IQoIAqBAPS7PZAWWSMZ3ESOL6NrnGIaEQV8eRN8+ro6BsjLAdkgKYZ
h8Wnq2XMc+qO8E45syitVqpU0aHSE5jOhAqh3ZvqNaOW9vKgo8QEwtprc0croGld
n0l98WXAM5WxFGiALvirfcaniIMLXbhaMRQEHQAXkdxwF2led1UTah9DkOHNpRaQ
FA9zGVyMsXJL+1HmuhCk7ITF3LnaGZjQGHCx9SGUYf21KIL/fz+iDnahOJWgsume
Q2a0wz38ZvClISDS2Q7FjNnl+AXKjwU17/vbEShUcx7Hygn8gIvjBIsvkodLMwnX
ICisJG54x5NE5wohwTsQQFFhRl6MKdZ929lghctZFZ3bZ6LHmwzARawbAo/KyQ+2
3gv6zYhZzDlOWMa4IoTyb5g2SdmLTSz3R29TUa01Ot3AuewrNKIgK17tNnTtsWxS
rfifGNO9p1VX6cfNlodekvJkT58j0WiXA9kTp3piEkX6/Kn/bDPgIBOMwXeAOXXz
g7b7S0hgOS1VXtO0czG+poyHELfYFLhvtElz2iVSr5KjLQ7oQTGeOX8eCp+cz50V
fZvzPlUi1j/OtcAGX8340BMaLjLStp8ecnDfU6fV1OhK51dw2pc8wIe9YT7VT6WC
8khJ2qaAm5H62YHSnEKX1UZKUmN7EXDnRf+YfWo5aDY8IuBwowCWExcP+I/XWIWc
fftPJRhLXlCWBCq20h65/RvbAfl8WZqLC8kgMU5fDm9tYCfNmei9pvaRSTnFbCxF
uB8UjYDbIpw7fDfxUdv52kMKHxZKe4NGi29wziyHOtj/2nLwi1iGVQEVWut9ggpG
lOzvVH+wx4B07PgK/qiKpuVkSo9amcUmZ31NQLOtYPbx/R0aMjNe+AXuf6tTmf5Z
aPlR/NswCNCFJ+N3KmAt2i/0qD00ZnwjJ6Frl908KOMT+scNdDdPSZa2/naxe0wP
9AxBOp3O2MX0RARVO986FOZPrZrb1omF4RvB9vvhujMU+t3orAEbrgG6ggXTbOqs
WME532vIrWuRNwD60XXCQuNoBRmofX9wVrtxKGAoxGIUhvZtGazfRD8kQbEazboU
b7y4gDnhrDNZ6XEN1TeSosxz1+vniWx3NMsX9Wwwl8/qBzctHzBfXoEL6mPm4J3D
L9MHaEZA0sOk8ilzrFduIB4M3hOgeh/kjbFVpd+pFJsPttnsGTtYbIE/JRbQpwKj
h3YGT49qNmCmXZsRV52ICRhONeL6mYltTaqo5BoO0zpR404QueM/rGZ0qV2egdeJ
ur3/SsXjk7/Td1aaBy805i/oLPnbDl+wIZkg1L4CcD+2z9IPhHxHMC0S+wFKeBfc
25dtqrKi9L043IWg8JLVODyJkERJhcst+BMcMsp/Wx4hqL3hSVDgTGa9Z9ZwEp4z
5ni8uIgdM50bEMAOPSthXXJ+FtxOFgiJbDNPAG4zLKWomcCikMVI2S7VfPs9EyAW
RmxxcLw5wbiKVpxZElxiBdSp97yT4IjhzsBKXe7zrNYcgO+1aJOKW7jK1nAq45Pv
d3a0zbWru7tdpMilFOyqLf7K1POiEkSWKIf72alQMb74MHhTwKHR9QV9CphZQsIj
Wl+aLilP2Ekaw29Knfyxl1OUFBTWpDpEyDA6zOZHbTb/xmj7F0TayurBvdEMLwa+
cX39u9luDvkZYrqsdueMgqjDeEYheH8TI8LbCmhHIf50l0P/whkow4MUJfvoKuLd
pXgQeYrlFY5whxapNFDFqKZ3SfHYbwSTAktJ6//YcndbIieDD/flshT5Qvr4JaCF
GVSD5N65e6jDKEutiCJsSCOVqrWUSGIs97WKWkqDwYXa/YpnKL67a3yhdrxEOuCZ
mW2ebTGdRhegmXpet8KIC032naAXOS3J4pbH8xImGXV96P1qpFEUZPFTChtSUduA
XbcAVeIoKGVtxtjZlTFMI0fUkFgNHkDJfJoMDBvzbebtbXB0t8q4DqdGkep2TV+k
zi0qTcpzZQp3C0augQXJQpgwBEIj+EWk+Hb3mSBtQ0uqD/kcWNTnRyU2rILIWvrd
tVCaew12KtZZFSwtTugPYIA2Dxy6d7QUZJfqsFqXX9wzSJG1yIP2C7j4LvMGzGp8
2N8LTcm0/Fbv1vFXEKJmlEPVL6n0utdhXhFNtv35uoQWzwHwpXdzOhR5jNAVD/vK
JLuDZjnKobfjoYLL3RbgU6AVs9nC/hOs+l2ppdWnXYP3TLMxmGPk4R/f0eszXoD5
vVzvo2o81AzsZuLuJIgho02ZIEIcT8VfFuhCAQ6MhZ2ZNN9bb/v4JkmUzfdYZ1hS
0kzx9yCHq/WEoB5GE0Xa4whnLfJLT560W7wmQGk1HD5SH1gwZt4C8fqTuYCRV5Hz
BrnvaYBmvai81R+B+nhN8+WIyVKTmJIVFoPH0499ZFaMVjzdCHjP6hVjZaytOVSW
dxv034WoZCKyPHVycFX0jMVL3gEKkhGwPvBXGhBesCO257Is47NbUfeWcnS+WmAx
WozGDxgI2DYMqwdPWNAqL4FIEDKaXijScQfhrlj3Kwptq8OAGiQya0g7BEOwaLIl
OpwIsJ9a100QJl5zc/tr3Ph4k70Es5sr//PPFpNXoioJAGa1/1yv2+abFuW6jTeo
k1K9gDoUtmjNkJHTuS1S6WIfTjizFErI+GYF6c8BM0y8X3gbHb9LPs9BB+ZxcxEm
8xZMoRFF9PVnePFp0v6pOYD4rD25WDCU9QssHoVad2K8WZ76a2mHmh63d+xFe7yY
q8/40Cyb/Ko63i4oC+5nKLjisiINXG1nUNYYp1oF42FyjE0onsgBzlsWhvAaC4cC
qC9DjPRsrMnY1WGaOcZCksEIWvXuGlbu7YQJePsdS6J3Erjux9bgXXE0fH9x+694
jKqfqI+bhySeMW6H5Wftuh89glRaRAhaN5brbqVSPWlLlUog34A4Ru7PqtmUDWxj
90+tWUIVlHp5/pRUjcEukl7QxlhB31DpttKn+PiHj6O18dnJeVSpITrovIzVoS19
m2LfYO1pYouR6Wa7LJF9QGmYcxZ7HutbaH5PZPUSh/xfJAR6kOoQjxQ3goGlOT99
IWkJ1XDuqO7gOeqX2hBEzMQH9b+R45rXOUlE/6PH5WNfscHQ+3fTJY09g8PP1qDL
mlfHyKPnzK7CuN6BFoxf4no4SAXQINp6Q0sllD0XABb89AuffKvkDROylrEQVMpK
IvU5+dj0ETmsZdBFN+UC882nxQPRwWH9aPQz2hRsY6Nr4xaXRYyihmmupWFT64d2
paRBDP0W2lSZ7wdf1nBundBX7f+oDosJC2o9Yptd9EHDkBa7KjqwXyQMV125cMKe
4iGcMkvu+TsCU3DYNx39r9cq5kIaB/j45M0xiLf56fnkr/MJ171QXoIO2Y31oVbb
ronBA3ofg9pRSV5tac60nS82qA2f6GEaBnxMXWvfb0DIYOYnPpbfqxZ0s4EedSgd
OuhEAAKdnor6ru7bySedgbF0zLrtn1PO5OyDn7ujRkAo27885agkzXIH8RB0IemJ
Tm0twNHlgBb98uHnLSoyrSiG1V8UKEtYybLQD14CMgiyuJKssY00q44c/12ofO6p
cMUdA0/QSYFqFpjF5OJq+MIlfsFnreyi9OvvXfCgjtmBtsWyM/eRSJZ4ymlCMtA7
XNr5PEgu7xyN59P9vv0dmYooh2KZ1yKCS5hybu9dEBCd3dV3452KvhO2pLk6DOYN
8AMdWa2Jf1JYqWHngotHX3TvnzDsqR7TVc5YiZgBE7AT5+uU+hrXYJ2wR8r7nZYO
56Pj+sNc+Ue6sq/w/LMQVi09TbYatY5MoxeXu+YhxYWmyCGVNHWebUzqpcioOBB8
nR2Dz1bof93HSsETMajsSzkJHWLwnQWmC3y1yQA/NfJKqwwqM0qszc4VkgoDkKBF
HpWcO6cItb1JlBsE6u7WGRcUe3qBJIVJHdeoJ3UbUCI6IiX2XuD2VleQP7pwTw7k
QOQnp3y1CkiA+GsGkcrIaBUyZQnYeJWZRx/LLk1OJlv6rfhYLH7KN77F7Ax17Nvw
wVlOmd/KQati7RTBz6A0cp4DPdQAffMY5s0Kcqf6N5pTOmvHHrJOUzlXa1X+guBU
OTjwQBzMtBFfxy36AWUU0Q/BFpXG0HBP9SsXHRKDq4TEG024SK3Shovx62n/l0vk
UlJLljhpzI3WeK76VkiiGkxv6NBnIphF8dKTfhurJN/CAEEmgnqW+WoRhmfTN2+2
xEH4tZ+TQ7j7IPkRJeis7gRMIQqgA81vg3SU6pfv55gVUKu3aihiiDL5NX5NIW5X
cuWWH/kUCq3gF0c7ycCosojotSulNfN38jZad5wzZasfN2Lb3WWLTwMoFla5WeAl
V+ZqOqm5yb7UYbXZISvcFC4alwPMUoKjQnlIKJF4r5W/OFntr8RIB0KavLr/jdNu
2aPrJxFjZZezr1nbpgTMtPkZ2kja1y+pbyzVSj6j9BzeHllj8WU5KUhBIRJZ5sFw
UMpo9nzI82eROWFUFW5zeFm3fkutvxbIsdFMkn/Z3XDqCzmvv5kyFMJji7RVOQr8
WoJ69oAGYnZpWkXdMn0PuBo3cHKEHHmxebRpzrLAAG1Fu9lKDTdR/BHgtUc31yjV
h6nmuWG9hysqDIIesw8GdbuOFPzGuW6U5w0oztAdfPzSVdNWRm5g3I6GRb5lqs9f
FKA7IBdRZPWEpWxFPSLT66wgtyeNXIrbBrpzABNoWF1tnzXCNh4+ayYc20xCp/uP
SCzR6YzBZMnakPRSkQXf6iHcWODrEhxrxYQSeyAHD78wf0OWEaru5GMCPjSC9/TL
8hthvI7tFirm7aufvGHSHg/AT4kjHJrLdQZEUqEsAuhkGvZIjci/FJlY3PJThc+/
DOv2FWwXRjYT3bh7NLIsIn/gHxjBeEmWG3J0sh8RRDtuPiwv2zbm7zrqfNTVAMM7
E0HJFRmkbJgiA+8REtF6gpjcBnX2E2FKrmb/ycuYS9tf5xLDi02nZtS+HTF+yibU
fL6Akxfjb03n72H7V3Lb88eiBIvq0ksZ+CZtXCoLDhvK6HxhDx7lADWSMkttVdTB
9ZYJ+sZGokr62WM4stRNCsToYAxxhp1tQw59C3L9R83RESa5+2r2/Ktmm5W45pm8
6eM1PGBZE33lPTEpOeYIkfOtkrb5Yb5ShYIYm1UsB33nykCUAPMh+BSOyCMRALkp
NbcCk84s4JA5vIpPbCZqe+AoHiHDT8jPSf9ExVFMVYKe42/sOj0CAmbb0A8DKOFK
RXjj6IATTageFlFPWYwF2V+7NCHCEqbuose9REbBr6DTOR5gB89cli6Qcqg5sJKb
tDmRwufBNspAc0VN6p9G0BxZGAZ9qCy9Lcs5i8cipsQGpRXMPt1GuYYLxRsuMXgz
zeRB1AdHPpHUoUxDOv1vDb/V3hr0BzoB7W0EkNMOtbJ10gRMkvw2jVK9uog5kkOW
QqipHDp7TWLDGMZedZxohYGLP3tGFrXkJRgdSTCbM0dMNvT0ZpUJ4t9emNzw8BVU
rWvv4nupITgcOJciQ6H6yAAziTKCMzchfZNoHph7jLbp+rNdgYi3twOxLtbGmTuF
ipe2ibdu4HEdBens/zQndiQpmrw9J9+7kGHip/A4QfdVlxkW8U8neqexFNDeqeXn
jZ4JIu7iLKJhgp2bnRMMaL6z0CZQMdS6dzH9OX9R/CfUqNqZUUKXW0YzCPgsNJbS
DwqyioWnLfV2Avc450Zt+QVpIcMSfp3lOC8dKQR/GRANYxzOgHbV0uJJF3baTMXu
Nr4noakej1fCJCmPdmO9bIuy/AZSXN9ETjBPrcVIUiegzlVwL2zryTm59Z/sHNsK
jRczJ1cxgEtmBp3ewRb62NxDPYbDssmreXiWRpgDvmZda72D/rzLvPezcbYKSdBG
t4qglsAc8QqEfZQ2CuQxiJa+7Cq+dGMlO7zCquAC1FQ46dQl4H/kWItmn6ESTV3H
dLR9OCbgxzPPs3PoVqWZwys+K3Ian87ppGB5eAxb5SpSZH+Cd7GzlSCXLiNOEKXS
PBcbR3tmakuoqa+ZjeKs295yA6cAYQPRJ1+nVqtknewa0wM+s7peFXiqhSKsY+QV
VBfVmamRKBMcz7Azf6PbVXkucKM7DaMxJEI6Fx9KVkWMnMeYpvfNeK4XR3/J/Vu0
HeLnP7aLLt4RZRt/uBBmbCDHX92TWrZTBcZc397bSuwxpbUpLUqVA+kGCefxi9ad
JDiteuu0Pkjz3FE2MT+V2/GUJm6nRm9P1z5oiFZoLn5NGGkFleOp6syMTqSXO9cS
qp7DOU+H/7plZEVG9tlZBuC9TlQu4HSaLxY2g/DcwGs6q4CYSMqHpcV/6ZK7j8xu
GZso/M/pNbX8KADqnO85aijGMH+E4m+zVjep54RAZBygoPhGnzAVZj/YqnNxf5aM
EzdtcjZv22fePIAl0cN2IYsOZoZRmGkNCvknu3fFyaPUalOCRYMKSYiJk8Kdg09T
KXnnW5249RBCij+WAExFrNlL6WHWTcv1diYmx17SNo4I+zxZ+4PGCT6pA0ACibpL
vOBQEcJ8N+P/rmdaSAR7jg02vhK5J1G10h9attTkaU5BQoFc/TPkg0XcVSEiVHPl
x/wdMD7zTkgg/aNG0liJ8ef7y+a7m5hpaPA4JHlmkrEVHZWRpVogbiDwN2/0nTnW
pQGBEJOrCI7Hllgi9EHXlFY0uIzlBbn0gqh33KtTzR69HY8CFmADunLRd1xPjkbx
LIH4Ney0GySHD5HbV1B94NW5G+ZLPjsGb67sc8C5bxSpAy1FGf6r8q7XnPC7J+Iz
jy4yrI8vlw7x/Dfc4uiZvaDcZQFXqpZbhDx3lIXR+FPU7AFbYqDOrZnvPHnMyMEb
IWevkqxWLbxAfvCLRXphu5U87XwjYTRdqKh/Y0TwWxdivICq6JLgefb9OgRRKQj7
8ue9UylF6hQQS4qzl8ns+S8NRsB4vqRnEQ1PNc6JtmicnhFHRJfsNEc9A7TskBM4
YAoTMbxVR7Lnh3ufX2SkDSSAKYV96iozmRI9YiiQPCGu66w1KbgK7LYhv4FGjMyk
jRcpR8WRTkBMn1ZcVn2P56bXasjyoUVOat3R+1LfyTveJGqNeSBKvwvB0bTF2Pxr
1a9pDVwZk7pHZ5iaa/jqFiJTwE0XPQ9gxWof5YsB+MOiNZ6e5LDPrdSutvYu4Rb/
wjIMouSJR29Ytr1lQ/nX9QtvAk6nAG0iggm2d2UvU8UhttKMWHpqAjwZYc5jDkDl
m+ddwMP6c+j/ge+a+6/YZTzSa7akfdHWiJn9FqZzqHIhgPCA4NhyFu8x7swLG5RG
zh65tpOgqJs4HP2Z2vN5BixgSrJQnXtZEUdto3ok5chyurLHMkCmhTFvL55x+/zf
fT2nkCDuB1f4CBcgTFtalY/cCUfhrie4dll+apt8UgoeE5YP6JxjEJqEbu2ymkZ1
HAoq0MPYGlMizpxRBCtNoxiHYbDsgAnTENNOpznJxGuXO0XNnQQxqe00DN4FOHWK
E+INL1Po8Appu+ay8r3MQeQWx9IltbRF/Ldw+m7gAyns5jNy2jEG5IN7hKuJAaHB
SdmCY5cXXtQgvWGTPeHoAsMHilXVRDufIy6izbKSLqc5kobQ0kaCD+2LxVh26NpE
5VAp2GDQaGV4qByt3WLrxWToeO9DdsqDKwhxPzTffDg0waYyMYoK6BPQMgS4VBM/
dW/8W+jTQ/kgPA2bfdbKf85gYqZNRt/1BQPXUsDn3zNz99hcViLZty4mUJcjmzDv
Xd0KmlYLz4TD4W7dXnfLWEE6gtR76RgneeDkq6WN3pAdi72S5hZbfWVOAIa8415g
eh4mzB6B67qgREkdtlAElX4QqOsoWjXxqE8+iyG4sncwgLBH2/y+2C9V9z2AD0pu
xSe3lVQ8+k/faojBjeFbqC44Mpo0KIVFZ7AfptZZh56L0s+FPaxkRqglWR9ndYaB
m4nquwwUL8iFSsPCOZLfZzsWtZSCPsQpsK1MDAvzfceAEw2bqMD0CywNDm8dAGEY
rfj40ea4dczSQXRBVlUjFpTvWh1UHFCqXe/eiP6IDF273YdJGjn3tNcB3Ck5zlVB
mpunCnj5lSzLNe0msu6gDdqbjttO1qrlKOb94gSxWzMfLtAXl2RD/8ged85lUvw3
qIJyVJa1QDVS/3L0r5K0HlQRfIV0FR9IWMITwkbN/uypa3YVv4H6Za3z5GDERKeE
QcJXyBat1OLD+9zrk9Hn0UiQjqbMcZLE10r3iaYzYNAEqJzqCaFYDGWJZ+YbwvJ7
GylkAxLXsiF05DYtFOYdoIBmi4v/FgIZ3etpFtR8xVAhVS07+gjNrwaIWSGLuUo/
sbP7wKDtaND4k/4AND0yGTtKeVJ4dsoX/YXbCph3pG6H2Wn3nD0HlI4W9GtEtUyV
m27P8hIRRo4HjsgwjIHPWeBWtQOAJ27kTh2P07s1RX9YyJmd3qAG1uMqZaAdFNA1
sWkLeTaoYJ5sXNy8iNrV8EwmWMGGICzwCGp/nDEiyGg3RRqYp8VF1lATQJkI1GvG
3Zg5ejeXdvt1phBJxwycS+pxQMzqzo96+CInXaSyPt2WYF+qu2Api/lvGYEJW9Qn
XPsaxGzl1ieTtJqs4iF2kd6f/Gy8z7BLW7XQ2cS3lbLpZ7LlDL0h4ReE52piZE71
C20+ZDqDXyndt1vsmQFUSnti1eHLshFI+54LAVo8roUxhFoDp6BtQyPaYmsVGc5M
w1qyCSqZcrh88m2H11DtyBToJJI/H6Wgj/FUpFTgv+iO8FhU52e8XqPtZ6wQQCPF
b9t3Tby/JQMR7yiP53m3VR9Vk7T3QOzj3dw/kSkOUB0BYWQAVKH9P1U9g3Stq8EM
APp/ywOXNcqY8JOD5TXjADC9DMG+OTRj1+8wyALuzjXoAFpBAWcmBmdIgz0DDTAV
TQn2ojK2ep71TIPlBJvnvsPcrpZGaas0T2DC511GM4lmN0WXgpzsxIv62TDvDxFT
wsgF35oNcMQzdJpNJnIl2rZ7iV+17CLJ2uYSdjYh2FPp8sZKwLL2nGJOym29gdix
3wZmEJM2uefixXfvtkkmCbJoYRbvkU9FBzx9Jo/XlLKMLtM6BP/6m9cwNbdxW19r
QBPA/5W90oXHua+dg8vdOptlpL9FDNkRkt+WQUftmjhV/Nrdb7EHL0jfpJx59V/R
JR5Yqe/Ne3ShaVtPMSajHTYLDzI3yrGNMqJ9AxecuLNOgjH8SBAa2XW8q5Z/VOXl
eU70Bj07cWxFOCTJ/FbPRAfMRSjsJtztNo72v6MqPa8YbKKR4LiS3A2ZGxWK98KN
ksPXyqixfN8G7yitNQsalLomzopWQ4dPJaanM4JLjx/8eW800wQXlyG/NjjjnNoJ
grgka10DHdH8NzhO+mKHq8FIzD/3Ov5SBQ9JQ5k58YUk0ujZHXJQwD16k6ixpl1c
Uhtt9Q32MhsquCSqW4rRYH+ABCb53iEvLfzy4h6znZHBgKRHdN2FCa8vvY6fZH//
Q2q6fkLm73AtIsOVB9eXxSwISn1A00MXgqFYz/f6OB5F+uuIHwr8b2bM+B8DKHwW
cCJaDWzArHlZUrq9A26MOS3vXsaWZ/EeZGHeskfJpHz9puvDkEkoQOYq82lcIwUy
YMMspXpLux0CkHpTBIR4p29pOgaoKDHBfxv//1lKlqTQyMFqgmfnpeziSCzvhNoA
ESzUTd3lUqHP0ExMFp36lqSqHbuRT0O0Q81kDFmLN9sRPS8j2v8LRgQ0psTJYbZy
fvLIZqznNg0GidSQyd4O/u80c5A8ASzok+oU2RjhRiL7xwtKc7lnPNBJ+GhE+yy6
Ad7Rwdje2TnP7HZy4DOQnRGUzJZXs3Subr83YWyvViNZo97/YFvzGMQjfXUfc49l
L6ynQErd1D5i47sDO/YvzBdrycJ+wnAbOCdelAGzKsOJCGe90+DmPWnEqm8KCSbM
nMeeS/kj7iMGz31hYzGWLkV1MgO9WTf+RnffmxW7oznVW6l4arpzBvdfkOjFDDCG
72ijT9IoJKE9PCwBdrsjUNvLC9bd5SP1CquhQyoiWuQbWY2//PYq8nFLB0qmW8Mu
0dEL3Y9MT65m9jy8Xba9F5TdG5dbAvuJ0HZWz6x+8ytavcDDDxySi6zTe0ZVuV6E
c/LuYDL02bQSjKiVuA2AEWBWcud6OVANg2mh8Snx/HWCuHQkurwHIc1U7fwrI6VQ
HVLscPI7bENV6xi9W3TB705E+ZmgbZuCdpZBQpSFFD+Fp03qFoxAxWJB8CaBO/1n
BbGpWzHRxJpxV7xFzyhoPFgUtaR6O3Pcp4fJAjoX6S46OhqqZOjq9GzmolscBrkQ
TIgTqgchw7kd98VmCSEOPr3fszcnY+TEDcxnraE+lEUKd4mlkoUT2ElHQL4py6Xv
Fr2bYulx8QliMKGhQJ3VBod/gColTicGjd5hz0Fs8+KbjBoqmfRbLNhnFJd9qfST
sIuzMcVt1VXG5mf/jqsolb+E6bCA5UG+lTPWMY+boLwNbgvOnrxW498/ggkpwayi
5/JXloE+3s2bIN6ugZHPrKZA5DQzHYqODzm9qaAwZibO/dJUWkA0Gp+j2z+eCQpI
fp2xOb0lXUXgpyjsBLilvSHbdMsRyl++J2A8bzRlyVoAF2a/MK177ulS+Vp54GWF
/0ojhSgfOOleh6dkVXFIOnmBWt4q9aGIhLzaQPEQrO1dC8nXcb2DRCJOM4tHbZIW
VtcdrkgXMYQHcBfybUSnMEL96e+c3oOPhi4fNOPwtDMYArGqBtxVkOAn53++Am+m
sTqsA+HQv0eXbOZhNPxm0iffNvm0aahdkWZ46o+VNPUQoE764RAyYGaPefGfIvwO
L1PWKI2dyakb3PQZDaKM4NN3M7arKoDMjzxgRamPr/UQurS7DxJLPjd3Gq7mpzIJ
3BjmT4zJhJvDAxvWGa799qgpe0/FIQWxBluBcf9WN2s2zGVCQDdyTKAKUyJtrjRg
cGd6s6d190u9AqsD36ENdwynKrvB7G9oCzjiAhVwaTe/1GOUGWaK64TVeNMhO9re
qOxEimG+I1TqMMVjOT1BeK8DbfdgaIau84bl/G27ShrrpDNMtA3NhOqeQ0tWF+nC
zwdem+ooBtWWNjrhqQ46qtFgStTk8jyOuRS465nymlGC7RztO2uS3Rlbmczl0xvR
Uwpn4hs+oEUHQ9FHkKq0UDN3ZJMwgsyAApIG6o+2y5AuSkgO/222VQqwlfBFt7qd
huNNhp1h4OvfpQGDE9F7gy1kyn3Z6yaCCrUJ235UFKVXaWcL6y37qcvedoTf3gAc
+Km35wj7TepDPugJSJoV4ARlqjvBCPX0+YAFSD+s3WDqLO2/6uOJ+YZTrcL8UHuf
Qz5DfXG333pheyVMLG6yQ2UR4WXHjLegqECmQTmDtBKTXBc+TLQO/hYY2pHTyiWR
d6Mg1DsUazVwfpO3zNDQa64aMbDPbtzt2TAYqEzRbDH611wlOtFcgrglMWAn/n7l
LxaCLuj2mWRQmyWRbm7oIt5sxVuJqOtHxJf3/KWKQ7LQZYGgPL91s+ycVx90N0Yx
9OP4L836w9IvggOMHqhGU0Fnil/lrc7GUG6xtnKO8f6l2Q31AWBDzS0btuUDilPq
9WT3wuR8Ze7mmdC44cun62fsNEQc9rwb7w38ULLRei00fPgy0x6ft3pO8Qcm9VIl
dbCgAngZvS+Z5c2Pq1MaFGpy2kEH719zQXHcLlymDK9h4fgjEdCNLL2xZrbCGKal
7V/uD2b8iNdYQgYcaFldEHaEFe3tFdWlm+8atMq9Vq9rf3PlPFITXher6JFZQhLT
TJAyQmwk6ZhfFceX5v96mmO3mF3STrAnWAwhjBcGZlEVNlBI41Bn8v02mmz/So0X
dz7RWLy/dhgfvPxj8mnodBF0qARaKoQmk/1cWdoqO4agIzzlIHBCBAtezOkNfqi6
sTK8UgaXus9CpNocTpvyebNLibjwE34FYTtbyL7QnG/pDUIV9gtD5NUKTA5iC1z0
uwEr1pFJ50BtZkQrullBasU08M3ezrdXdFcWWTdHtWSqRYpaKvy8ABG/lW4Jkus0
r3vYeETMWjkzKrfWzG5UWwqdezkJcxlbLCjmJqfsSdxWor1999z4/10wVEb2lVC6
jpGQkKovh81jSWWVjyy4zyLs+DQPLMYecTyGyzQVpDBz4s1LQExZ40B1xxiWjYGF
rSv0kWi5XwcXCq1SdqwKZa4pqBdcPa9DhrK8tvgg2RV9eD4AeDxouj4xtpge4yeb
8NFf5quX4feKS7j0UBCByB10Rw7ocLo3rWl1dlClk7hLBXNF5VrnxxoVxgQf6XEo
ghZumkdZcGMpD/CjyHvDdnvUZYF4zLU1A0vyXbkF6fu7hZUwHHyo1JJaZBTiOOSW
MxLvMWetmzwWLBKF8gGgkHOuWcDKeTJftRKTqtfB8lL+dtTW4a2RKVXeCOJRM6kU
BVZUUA6/3COoAFo/TBi4f3OjMm3GAlYMp37tmdNawELLT1+XOYSOlyifY+MrjpBe
3qkBDyC9fVN+pdpk7InBRfZp/6jQ6TCooILATfq62R8k7t9CPvLO0rP/WriXfC9Z
CdbHNcFfnYj5MFRSMHwNUOzHoi4uqd9edpr4xey8CBi+iX4iMFGqxyWX+j3fWQgE
/AEvMEbljyIb2fSORFVKBvxXyn0kolk+7i/YMqEdjk2aZWt83Vmpo7FiM4NQf8GK
5CZaHfJA+Y1RkXYtD0Kre3iScS/qHR6gHAhYraMY6b1m9ZvNygAhWXQHfdcTMliF
Vp7PE3KUHq1sI1f5U4yraZC3jLLI2YQFbql/m7sPqfdPMeesHzVGKxjtVO7fGtA7
nkuY4TeMV+YiMcujojRH1v0fDsa6A4+ePWBDbHtCWPOTSqlk2MzeFL+nN996RTDK
YdCOO3PAd2tnQF2RZinFzNHkxPnfH5hF/6dwMMApEAbw6cdnb3wtPq9LUQsdNexC
WI0R6uvGU2g2w89S7xp/Etc2aUV29HKgjPNXup2+YtqApSrLsEWXkvB16X/h+muU
V2DKWK5avKyHitijkDr07RWVfm35QUmnVyv9Cj68+ERYyHXlSnOasgA9QgPhvYIB
Y2ABR8+N+8XUI4/adm3KN7tPvNYo30JZhtuJu4N05x9Htfv5lnbWv0tvZvD1agWd
RAGK8KcR27D9YXQD6GnhQgxmlH4mL5VFEPNr6gu+cavU89dxEGDEmgPkjV7lUP2d
8ZJnV4/ZO+gKuq3sfmHrbuHux5OuSAsdmwhIPJJFlEftH3ZORu1/4gmqFN1Nzwmo
2GBft/9DKMU26Ftb0fZvaajaK8mL2GQ7T5HINpcQAaWqSa+yOAiSUYj68zn3MSo7
StcLnQkix361ec1ijqAGCMVgLSGjPazLeHwsYa7OXlfJRi7U8ErxiZVdhEhORq0V
cg18CF0g93i9wx6oS4HgRbHAbGk+OdRj/w9DPzVKBa3rd4a6NQIV+5Z2AExUhekr
mWOFyYkBKQLDslZnnXRgaSAowcVJvs8UC+iqLdXYggZw7MkuDiSv7WFwa5FUfxtc
DzsxR2I/RzDnl8lwuLfgJYjEQCAtLwNAkI4s8Bj35/CBKBPgvajb4RApgE1NfV1i
7hn1RTqh0r5+9jVmWqy4YlQiRFMCbvqNjKN7/gEEaKwOpTWHsvgX1dGu9QrXyBhs
ZJaYRxcChcoheEDpR7Zs41zBRRaQj6S18jerVLyzY/+fJZjApez0UJNzmqyEQTFU
FaLx6UDRnCLMvCi14JoVi8fIOoI/rcQTubvZKFMEpfSdyHfjjke4KsLFUD7fyQGo
XwXRPgdkcfv6uMR3duMGNggwAEQSDafXQbi6L7GSgbyYNJdcd16+0qrpfW8sLrOy
3MFT3j4xDQu/Fw1k4eUDDaDbZIaU5eb+RXd8K2V0VzmSTiE/5kqNxXysdEL7XSzv
uxUw0Flm2uU5MdexV3EENR177+hilZcIg3jgbVAqH5ncxQ6Byc4z8AAgDWXdva/d
mUZBaG5RK36Wbp5dHeZWcQ2JKXB2q3Z52gbsZ+d1oy0HT3QwqDKBjEwerIIB23RI
Ol/wxDr8MQ0xgz4b92Gz3TF+WCWW6aoq2/sF5X1iYs2SC4s9Un2iWOJZsvT7lLW9
YcD3V/AvMMdm7rfGx/lcWdc5BzrJn6MTBlj/mjbEjZQd7hVtAXoEpQ38208pUdoJ
TGqOh1myP+LKyEGllUeiLrEbln9Fl+0Pl1OcZARv89n2/LHae6eyUMJyTqZoxGzu
Pa4SvLVveHoj6bLU4dRoDxOT5vupCsk9I3tXzCD7otQPD5vuBr6STQ3JidWRALiS
Sbmewzzrqlfmqzz2lQ3EYHBuSQK1Y68GVZdofHHwY4/o4gRgRsEsK2G/5rt7dtzB
kk4cyyYaNgBiXawrt65Rc53EzhxYqYT4kyA1zef+EMDAE1GWAXt0hyZfv4esYcbI
bLnV6T/bLjBYHYCW5cRCt8n73oWVcvOB3yG/S/qlulNKuf07LYXcmhpkiyIiSwT7
6g1hGYIW7SHCsJXXfLOFBGcAkiA4hJL7i6yzI5+qZ71vUVqBRm/cuKlVGG3ybrp3
BnA9WojHaat6ZdA64ffZwgyfgBOjqgY9hDtIXcHevy59fEdV/N0i6YaTf3Pca7D6
YEjaOovMSl+33o2ewUUIO5BkbFdItjymEIKx9Zc5leLSjtRe4kdDhvoBdjowwXO5
NkztCgdl9zWZNkMcNKuLve37cRqCanZT8rcmkhYbeIrplJPczeO79YdQ5i4BUoaP
VjABgvDZHf/Fvk//LVwBEcPPgg6CyYxqvBJ0V3rsLx3eqgTQ7RJgoil0fyd4C65c
h1b/7YPWRhiI7nzCR7ejPcZHFCbkXIaf9JTJ5+R3RQgcv7c9ukR1trW2r2s1tT4H
VjicRvOxwGWNJd9HKHMJi30blK9rmK1PYAXfTcuqpy8MbDrxmpwSiMn8QDUXXuc0
hWe3pcWUBc5QQoXeHC+nq9RjbudXa98ODV6B3d9zpIXw5JUMgUrpsdulw2PYCLbr
cCpqAWNs2T8aMKhuGiAr10+4mACV6yB27x6mYT5Hhor8eX26TeeoR3hJfFEcjjio
ckGGnAggaNAT6gE33Ks3H9hcF8wgBGH1dsKJF84pHqIg/3F/V2Ib4Yw/XawIaOHU
v6Lw4tSY+CLCIUI9haimwXRYxylbac0GRZMozzbXSLg8M71yEYa/yI9dz3969VUH
JFgFJRadFwi2UCA6GakpRTpKH/Gz1sUNmhrCup9wdyz80NwZGjcYrJOhLLlZ9+jh
fzwGwuFpyw44GE6+ha+vk3NhC0MJdROaUrCv5IyB3DuVgRpw0ncQR9HJZFglJGz9
He3pD5p9O0S1e7UgQvzLJ6Qn7sSJ5o6UKGKH6M4UG6SOCLkqXgy6nhyDvh04ynFe
KyFojhaguZNC52tLOlJkIDGGifQT8tUw/PvtrH847qWLnB4BFj7kReXseQWDYIYP
2mDrWx1GkOyuBm28wMopiXBWQNwr5zzZ0i7a1k1pMR50YhVdx5v4yE6pHvShlUHE
/ZGbtumDTTcEdtUm6EzPGs70FE7qJREGmzR9L0tXOFf+KUeIVTHbvK3xNgRo5myD
AvBaz7rK1a0hsJjbxgWcX0bvP1Levq0jNcYKB2S3R7uCCDk+OXXNCTzpTiI/Xw1y
KPDLTY3loP9nqQQCYRmcZFhW04SYDzz0vYsSS7slaR+6aOcjSJvFpsyNM2LI958k
5rrLYihvlqr26N+6OfTCrvkySIUDF8p6aTnScIYqVflByHvad9H0Q6BKc9CRWkIw
z2wLRNk3r3iVyUHpsH4d2n1VX+DUuqk0EyaqfcYf1CkHuk1nY3ss1CAebYXfazCu
Dp3lfrnqq8qqOLx8O1v+pZyoPZFDxGxP/3DSzuGRtabLzzIyFnuRDKKfRwwloW6K
WkXDmMG9de4eHwf/1NADxULSWhM1iDiUDo+kvRRcYNUzT84fBXYw1M94q5sliySf
b5eYAKVRZvLV10qilJ+gC53vOhp/4dPzMe4kunh1e+OmDRnE64yVA6B8+QJIcpbf
M0NrVsIYOt0DXCZ+kc7BpZMMPX7g0+pYE/hgZU1J/Tyq9y6bnBHzDIvo5lSfvLYK
vY/By+uP1tDYOhwHJkQ4IRXzyxeTvVIm0+tC6TgztKd8cctNpFSEQ6KjwO280GH6
21pUhJqpZZa38w6RKVJwRPOKd0kvoaSoT76QRMyg/X9iG0dcVBNuN50igLx+uS76
Khtfy2XQAGQGsvcwfMb1h11qGonBhjHXVu/bDetrbT9mOx8WblXMgIzeRd85Ptve
wT0BFY2dtr2kC61JNmQBES1AXaH6W/xcwZhy6EKh6hzbHQ04SSTQ00lq7pz8Q/I8
jh88HUent4ynAmufuq77NOEVy6XorqzM8vA+qiOIK0DIKIYD/3dkkUN/TfvLK6f7
MY/8LlbClYsUS8n2lSXU2Nn+2be1NpnkD8SUpW6q65gwHiLmAK6/UcqGfg4+sNyc
8ZQW4EI1mn7i7qZKxzGovr0z+4JXrop3OoINUvAPfILGf5SZvAyQWNRRnmOPq6G5
RGwSK+JQVaWPj6jk6P4Uy7IwseErCRpr/X/pwwXafv2k76+a+4mMbK4WSSM5TqnF
a0edWbRG8MT/PYPSMwvr5XPamvVTcyMwJzLa9TxaLgALqacaF8eXAfJkbA5PItQ8
Bxvd6PonblSTq/l3fSfu9FtIKUAJpKepZkpdjDwLJwIDAFyauDmc9/vppwcOWQoc
utX3WFnbOYegmbYfeJJoWtlcCn7PjuDUxqG5ZRXd3eT43kg3eT1uolW9sQfLph2p
Xi0U+VSHDhzze+rQdeOn9pXHMSh7S6onOVpIKcsqWjHMjIasdZMfi2PbzGTc9Xav
bHgIlLbtdL39gh5vHIOmMbKrckrYxbmpKK8YQvg+7RqVyUUUXfKh7a1JH8gyp64n
zZPiCV46lRuzMDDsW0K5p1HLefY7adu8DsJPqbUIoYQ3qDjlS3fcak7pF3hJhnbu
dG8ykqX1AeDQO9LrgrAwfDsJ2uMFOGVvfnPq/6uoHg1EcqaCXBN7Ts+D2rtBO9Nl
EEinW38sy5VgVFsT/zpN+sLBkvta/Qw684ihMD2Hitf4MBjVK1O4UY+5h+3t3GRc
ikySNbponuvyK0kPeBVOpmRc2Ur9adyupZZL+cjf80EQ2hqPb13zWF7cJhiLSsja
0s42AFHeyQSMMIsYfemxzw/Tk2ZimMClzamNP8GpoIQN6Hz/sTU9+VQ5TyCv1c4+
UP8OqxmtVB/khKrxvDSxZrDaiVf/hB6WxpXkyfRO8ZkW/OR1xXwFCPl/58Mm3qdP
EDZNWrhe79IrlGvXdCU+bRFIS4Lfy3rVtcKJH/QKFXWNTMuNXRXUzZv3qZ5/UtPN
5Qx7q3+qbBb7te0yycBbob/bUNhSSXqiVCu30tR2shBKCN5ZVgQcmrDqygL8hJWg
TX4VjKinTUPd0ZltYniwc64b/4ScYPk858H3Jvmy26BeRzP+2QCsHQgi8r+CqqcG
uKiP5xOwq91OVXtYy5qcOYFgvvI/qEmM81a4MvhEfA3G2n9c8ScUJ+hw6mKx0BYM
rYvAFtVMZImuJLu7u0sdNe7CEk9RWrjpAY4ZYzWVusqLCdqMMrrzNCdDYvAyrrCd
X62BIFWZsTSvUGkBVc8B8wzuMwzc+Cn3l7AOSZblUL70NdAwB+1EHFabyOjOjhFZ
Gb9dMnURr6DuoufT9DxAXYqGgXQuvZc2WZxX1Jar58QWmQdAWNSbIu2S/F8atOqz
zXg+0UfaJX1QDv1le855nI6rxKshB2XgRG5lKEyHx5sAaXQa5AfmTQfS+qG8hz/C
N4jbE46cp26KdHYwQLESSoFcyil9law44ZBqSDW0cpGKB6YbaDyiC/Ee8Qwyra2z
49kFryEZS+FxYoRxubWB/eWvIjOykoZzFpLy0TLefetghLQ3XfZvVLxS/cVnjEQa
E9FV4f/9gpoFNeLhQhEotCDWV2AGfqES8ZA2VI2yCqRyGFtLOP5tPbwtHBNHeZJC
wiK2frdjzxiDGhiyn1Nliujg5Fcd1i+zGEXKCDZGKSJ1H/BmJnV7QJeF5FVRr9YD
/WnnEoqQf+dv4CRBs33k8isQlBfA94fpL73BAlwxaxKPT0P6gHtKYI8On5Oiqppy
zxlJrBd68QkoEmT5/VfwHajcZxJz6X68s7FaP+rQOdEuJu4FmZifF0Uqa2PZjWK/
RLmTIC+9hCAwgmbjYaFG4juBMXCTP77ub0Yi8WloDmnD4Qgv0p9ZsRGn7t0OCPb4
whumomKgaeHJ1FbFUlvYsCA+p5sdduiAgcGdsYekCL2dCSxARI6NS7GpLqEB4u3A
WYcwViDDDAWE9GbBspG8Wuvl9Z/pTjBIUqhPpTyr2GKgPoD5Cr/xn9qgRygrAOxr
Fh50QRhW8A4NLjyRAPZ5p5n6SOlB8gi7zG25+Bh79Jl6v/X6uuDUISKJgna1Xhqq
oR7m0M5auCJWZMd/uOmRwLiI8brdPGS565piixIdAfECepQyUkiLox3KrDKZ2vpO
ao9XH8Eq7zLahr1uzYke8OGGymJJtYyehBlTOBtDmFtFWa6YD689TvRK77ecMUpC
Vpa/qvHiipdW1ZBqkwqJh0uHQPoBsxSws6WY0Tz35pMGEnRSCQ+J+uN3Ng2bzI//
W1pECKc2FY08pK3WMkjuxpy0h6D/EeoYDAT/w/DwoNq/kyKT48WPsRk43a/BDF5z
cjHDPYHqNxDjAmdQOZTpEST89zfAuD4ETv7EBTtk07C5Y2v/Z8HFnZAMCAp7QP4h
M1fsKRojmONZv4dvjCpB5i+Xxm/VU1z6iolS/UB5H5ZxtFRGEaJcMGZ8lNMxnstm
LqO7cebgx9hhypLQUkHaAMytBWS2Z05hmcjvqfnPh91VKd3YQMpldLu5/Dg1eeCm
JOnVWv6rb1k2RkVQVKoRsC2+KbpquCU28qTbFLLvHNSIPPgpPErwwIOF1rSoqz6X
xzecgpte+GDqa4DZ/QEhPJ6At+cTo8WhlqVvCwTajCEd1otCgiXS9b/zjlRzzqy5
vXNlgyGHkfbm2mSxZvFsLgibVej1lBt8cJBmz5snvmKaZ68xHVyb0la3rwn8tvJy
rbOLbWHx59PB6ilVouD2G1And3wQM72g0ck5nk+D0PaQWOp0fYfIBGixpC4YwNfV
3PtPCzrg21cbLppvxCWjOgeyjUUwHwgCCdVZGEwn1DU1WV6Acn3RCI0jw389p/VQ
gTUZCn21+YH1epRgP/zKWSSAOHgTDMeSTx9yvs0psNJ+RCyxOSGwZHfAiXlL9DJK
av5+dv8atJpOf84oio4A+r7XuGNI0v9FqW1hlQv645tJHDI7kgvpyToHVqoqeN8Y
NunBodjhKbPmhhK9mS58X86etVm3c2gnWDCEKgb+u98hOvsg9QUcTbhhwYh+veut
XpxL11q1oPXZk08Q6I7VBwncQ3T9+DP2QbItvR0vPtUWbvlUr3zELaZVDcsw3tel
/QBE3yI2SnXwZu6AXUv8l1IzZBmqbcrv4aORdOcETlLVQT5X0cJbm1aWyhSeZPaT
zoDrEB1apLfpKNEAnrVwzDUGRJUkHuo9zAu8yxEHT/It+yJU82JJdiQgsb0fT8VE
e1LquwHL7rZRzC2uuQLelZ4jRnrt8uOSUATua+wIXiOPvb5Guys4v5cBEuezvoN7
riX59JwyjVEcYffvFd/Gwztjp9M6RRZCrv8KWn7ibYuAgyxPF232yFxnkBu7MV2I
ifpB41z6m++bQskybyKoTyedAmRodgiKkY9vNuPxBw8Mm0ljW4lmsCQptCa47CDj
rmzZJrwzACEvC3UzzqmBksl7uZEtk8ooRd1RttHgUOQDJdQHI9OdpsDKdJpKv1dW
JoN0M8ztD6EaPYc3378R2iDMb9kodSlfQyNbYG55dP9vzazjyN965zrts9cj9cvy
1RLNjkmA/o8VQKtrp3pazUpdJwQ+a7gePcgC2cEDJ9zbYVX7WR5mx7f8uxH5BGqu
LhLRrB3TwlIFr1VaiRRti16t797H9SCjwpOAwalu0sdOOJ8PU1USoTi7zVZIrlBJ
9xqZr/ZFMpgA/owf84ZJOEXw9gXMmYfaGXCVp207Gt2yJD+oltqjRhubUS3XlewT
zoFsIXTE8l6WhLdDvBNcBwHEsjZPjkxHUSNhB0yxWFmiWsVg6wW1QtvuZVC/1RDk
xeKEDy94TMBYtLSWHuzUAzh/6ZVkvMTyJ15Hc5VoOGEYJ3DuG2zqJN9Lu3KYXil6
6KBzdZ9ACsWaBwaD6soC0GqYrne7om1WFl2XYftxaTncqS2brT7qfCxcGrye5WM8
VNEgNfahYPcYPlgFlByVLjAYvv94p5RYjVESFDE6vXsJd94szHnJnTsTKnRzDDKY
ejqgPM0gTGtm55Q9ssPIFFW5eSjnYOKigm7cZ6op7vhE369FBwtrxT/zJlvlVH0u
d7XNpf7o80hQbbZUL+28k5nRW/WUVqi4dxYS9re5Hg4oeDM72lMvsuOM9fjGy97I
YhkgiwOOObhb3YHgNoDsNUX+zGAHLtqfJ04ASernTsoTy5JBtrSwmFA5tvARALCn
JSkfLHRZnnSUdovHd+TiBo/rZLenES4S7MpLm7gBlkcfccFhF4yh0ZprlOKKe8I1
VP1EVUF+vXrjV/pN23ZxgwD+CmNnmYNOuWfKNuUQ+S4Ywttwg6/734u4Qhet4xjc
YJNwa4lCr+7UWSOJCxs4yULluHlXc4gY9e/CgbP9lloAJlL5I7r0EZhpSVmS8LxP
TefU6f79E+CKpKF8VS5ubVzIJFXK0DJaVD5uZs9d1e8QpDk3hREgR8EIqOUpY48H
Mr1idN41zMpese9waud/XFkMv+iFdVjdPPpeinjZEeF4qtCxPRhsEAyneDUa8eBO
ZBsNYgkMB5o/Zd+w8GPe8Ep4GNy5jjW2/KQrftw4HWXoigJqcD/miCPbk1gvCdRq
tacxk7N351UGdEto+euJCh1Z499SE6kh/De2CUSyiUl7oU5Ttw2eqGsEi0tMuDv6
Jkdfk2kpLa1BWIMkYiJHoKbkrXN146EZ/QGiaSVr1kW/7k/IB9xEbrrTJGp4vm9K
E/JB+710UrF6t7+AEmB5NhH/JtbPQ7xH/J0m1lZUYOCHhjYR7/DyDySLkOUCnsSi
r024V/ZWw+6rNgqDGmV5Jfpr7mUG3a0fNZIo5RPGSkbi9JRQFXMBUYeyRDF3MDuY
HQC48nFnBDN8dAbpXB0VcLcBX/19jG1eNnExOyl6/HKvux99z0ycWtmN6uTp7Yrk
Z9a/WH4KNkRX9/ihJO7fxOnXW7PIq426YKn/+ujhq3EPC48Vyk6TM2R8sPOeT8xv
YjNnYePRfo+WtYTLIcRaICtG0pKe4i+O8Rs0AFo5mGl5em0L1r8p5h4aZ+f4bc+y
x4puhC9WJaRMGIUcGtxrc3ANTb8al+GYW2ohpgLV8g1RRmwNlQVTv5Zw291JEhOT
QtxcYXynchfNb0t45UpYsZvCaPEkA+wIfziP5wEudDXKAYxgMNkYlCBSHNAjMErF
crQekymx/q5SBrgR8X24W9nSq4/ArVvURvZWkCk0yqZeWs/g/oKMHEBRznUg1J76
55RQPqpYjKotMFwFuTGokayH+aneVxm6wL487n6Px9Mk2QcU7Su4IdLwJSmMbRyZ
LMai48o374mFeG3MZMw62rg1h9gmKlt7HNwTwk/MOoab5OpJOxkhHCidOwPlFtH1
HlwRqdyeWkM1kMbdM+rsHetPeX5/4wDyXVkHziNurxfB6T6IdIeudmpQdJOzgMlN
JyOivgwEiA0N1ZhKzpGgkZY7BUx1CvTl7H7t8YFkqJ2k4OlK00eQ5QlwJST/RUI1
LkIOTnUjo536ae8sSJ4Gw/MI2v3lo1fTIb3rpNif25RJw6/sCGrUCklzCt7CwgM5
89BrSs5ctD43e9miLBqxxUmBt6f6rrXRI03OUeAL8y1kEZ+q0etos4P/gOr3KutY
o3OiMTgxoE8Xb33WKZQ+f2FxBh4aBw2DK5SVMTJLFoLp0VJIRoo9ZyLGg5WmnHdn
fI2pFZPQx9sYOKHDhGCmymp5Ou6ERoyaBcrgcjNqxPFRkM0gaQnNujuCrO119aik
tCq8PV27IoEgB+I7hTijzRQkK1cWxSlLkFVbR0N1P2PaGGjL2NWp27DGQrrBtmc+
byRqbq8g51vqnoyNvtvfUT4tw8sR2petugjSRWcejFJcaH1YSmqVuevB7s5F9g3L
gSKdyoVbMT2EhE4iCotzxvQUjNTzRP0J9Qw1ZbIa2tm9KS3oaTrBnUkWe512C5Sl
9Row2/b4I+q1/Lm8BsXZTbuQJUYnXhKDuhAfkvSbi1oQQr6J+JE7gAn8ekuvmwg9
I76FN52wAEjx85WxvYevP/KGg9pNXKaWX7zAC+ISyuoxl7PPD5uvWcotQt3CxiH9
SpsX8ffDzhIYPB91NfkijSavRVLRkK8CJ7qBAkJnhz3PMSg7L2Eg1YcnJYbYNh4j
ASQGE8IEdGWsx1u521NwuBiP8U/Za3EXlDV+yQb3FrEgRnkPfkb8BmKncan9SAEk
WYWYLWegpsO5xSxBhAFEEBbPrnnFh0ZutLgSMVDaCS4KX31EveqvPEsTeqfiryIR
nY6ZbCsXGB5tWa0p4b+uLQmli9EaJl/LoSSG93/7IOhq02AN2/DOtQIzAk/0AM45
7jTl3vK62XGGWdhIr5HuNCN3J+BDPzm7s+jNCVIEKI5VuRe/2+UtdJN/4o/YZqM7
QORtQIo0pqKrK+PUKx9/6Ly9wpt37rU76KPJC1TmSk2MStcJOMlWT6jT0VBWI/sh
6E0ugNMLT69bu8rTRkh6uuFSFsTyyiZQevZ+HTnfMStHqSoSocKOHpyEmvpkKXgr
oyNZWHRXLLvZ4e7+mjTkr795908duwmfbSl/IsqQVaigd3rsh+D5enoAOVfYxVvy
h5hxyoB4D6xLTvEa9Xn6Tz2csfSCn2frRFIv0YoyRTaWWdzsxXUdF1CAjrTdHuBA
bgD3/1j4MVjS7HrD+XwnWQxG680wbwvJarB++A29WRHD4Kg5pYDpuWR0fiQW3Psv
y/1v3q7Miz6RLW2wQkipR+udMMPvXKsiZ54y+7OiLfuFwsGt7b8onsNqQnjwXPZI
8Fa7XtIyFmJ/VC7jBTxHvkm0fYBQXzc8foM/NKXF+WYWQQrhxrE+AxlFJhGHY1KB
xoS9ZXCQI/aTCRY56ekb1F7rJ23JJ88RmwmnUqiRaEsOt5Mi32+xj3DFqqOF6oeA
tHxMceQhAeoZDxZoRqeK2++So2VFG5AQBfwjpWn8ZBZ+rf5x+yHIT7T80in9aiW9
zd8XO6Zl7jZQgQX8619hEt1qx6b06B0UK0StKC5zAJq3H7BnfPrAankwKC8I4OQH
d2Sa52/z1w6ov11y9kR8nH0luXVnpPfX4I5DowGW9m1JG+tfSajEY9rh9B6bv3HI
F49+4QQE7IMgGLtKZ9xeX6YjkSIAoEMI4wUb2WO4DPp5aaq0KBG/HT21UwqAjbR/
PK+FNOrXWsWoo9nBQCfn5soh4xwDmoCxtwfLBRsFWFNS2J0UtemprQzUkRS8pqSn
tyK4UlPdJ2wRLEh9V0ZvpqeDU0FjTuOdxHm/uGZ38F68dZkoaClPWdgGPInOug60
kSZh9S0gIaew/NmkhbpnAiCWDGoSnRd57ArC92jVvPl/gWAwqWq1yV5Gy7MstAuj
D5C2vblYU1pkDV812BVWzRLbQwr9NJTRkzLNzboTVFSVehs84GIeRbn/oSADJHOu
4xtkLJl7rKvkAP+1VSauP/t12iDsTAzCYr580Of6+2fj/ZYkBXxn8pB40OgQHOHR
MNUeCHwA+heF0nWZfS9YPwNhFUEG+q+J5nInScKv3qyfSRVKIKdBHbPehVwsUtU1
G9xUwiUfFj9zhnBFuOE8sNW43xI7zV2vLy+e5mu+S316GD3AFfSTz3Wjn4X1NId2
WypivuSSdHWsRNHwBTgmZrIdafglfXdXKZtzvFFnjf3AnfO2K+FpjstCMO78IYNV
fx7jB2+qFBmBhclvlxtODFjYpIIZ26XerG2u3RcOB4egMRnKbACvmaLeeIEl4u+A
xRzIYQD6wwWvec+W0J3BVbPUK7vsPIGcq1Cowd7jA7DqepfukdN0x7uSdNHrjsCo
DOcu46HTUwpnpXZQMxYGW5F2d4H2n17bIyU5T+rYZZveBXUMgHB9pVKTfDNwQUu7
kruGD4G3R15tye06rKpeSPWJkP1wd4mtHda4IvkIW+FI69uBTx0GTy2MCPed6QvI
7HZIVlM+cBYFv51VRFkRI2P8PINDbGuLLEXjWypJySH9dCe08uNej47W33nzNON+
PD6V+N2hdenbvnf/jwK5bZ2t8H53IpFSPlGxESWnKMoUX+jREZM5X2xK2cEAFbdV
h4uInfPaE9cy1IboxGO8uHD+lcjqES7SxnJKGOGWREMM9iH9aknTSV5ebRWAj+hB
BXX76ZNeR+zps5YhkffTyl1JEfWGuLu0AZevP+ytJ6xZ7yQyWP8MXDMHHXznE6If
u1rp4BaRvD1nKB1gbARvDAFd1GbqUhlhfjLrV2/LRCcUuF5INDHKQk7Ig6tl+moP
bqc+Lk+YmPNDSdIyetK9nkwm7qmirgqkJfvJxz72T/sPuTEsN8ZPyVinmLcLZjxx
3+SgVy+D1TINjtFAQeGj5ozXv9zegfde8nPHPTQxslwTQrr3Xoz4x4KUFCgcEqZq
kBF6aqznj9+iZRx46OsAKda0TDws+kmxiuI2NrLhmkiVTT1UUJNszg81t/m67PX7
mIa6Qt8A93KUiaTbvuIxkVpqbKlsKXbwk7REvmNF22ZKY9DtzyESQSIpjKv42Qcq
ws+TvaYwsYqV+1/8RYIt2G3wVG8GItVUyMw8fXCXuOBIjmxdUO5PflHelolqFQmV
+gPEFA+UnmDjuY7zaHxuBgDpszee5uRdUi4Kn1cJm44BzLKTifadISTcNLhbE/90
0k60+dS8hn9dhHOMGJU1u5yOvIapqsma1L0+23OJHo7wL3yxgVUfTSYLzcfuErJr
8dPHNZBUTA31tSihgnbRN9tVOSR+kFO85IETrdhjsihCTKj3P7cHAh5WYo9CQyxs
UrgCPcpYFCRPF3w04rLHvJ3hPJU7pM14ll/x5wfESoyqKt+3mdGcNzTPqDRWvsOF
Q7lnJJZXx+V9OkspY1BDhtM7kKtR5oECSuqeXpPhTHOF0WCafhnb+TWKavk/xfhV
bAeIn6I3KayaRsDkaoN9Qb8w4aK+VRotVyC8viFX1XHm533ATNkvxPyMkDwG+pZW
QBkktD4wPCvxdIKPAPxoZKic2Sk3tOn8aY8YMuNfYLFoarOqcbaA/lVyN7GnmTmx
KErEza0OX4KXXKm4VaC49nJUBJeltenUMho59m5SZ3KSVdlH4OuNKIVc7+1tEUGJ
tlC+/iXjRpbGtMepcV7QV2DPeONzMT3MOJRYJ9yT8Gnt5xXwe4E/OWRDQQMNZavZ
6Ct8VrJL2Po/NAGWbtePYtEHLol/vO1KdHIWT1E5EJmF3/52Q/ggoqVxI6pVQb0N
aQeXJEKHoiXpfJgE6GKL2AL9yFk2yNNfJNcgEnPmB2nejzRPjpTT6BE6Gx+gay9u
hCQ5w8/h0KofwEwmeUZID9ADaDa2Rxq6DdD63JYskBMJwjNLhvWmmxkV6y4hv7c1
CFipzBuIJggMSacfoa4He2x81Sbu856SyoRANQ+vje/kWKDRtpCk0/6pBlFNrBet
H/LzsK6KhozNFhe79hGDpxwugPITA4U/8PH0hjV1ZEpcKv4eHbSZVDnP1GKSvwgK
gCqnYvPikeRZ70PefDlSF5BW+KwQ1H2IkwShqtNwPE9TLz1Umdd+vdZWHcBtnTiq
OB0PA7Zf6vpacqYR3ShTd01oGl4KS7QFjnUoL3eXpNTxsZCmdoVHg0t1ZIUmrIEE
luv10RUONVPZmmbCa6ezS7lDprV/JgaNV8EIILrabWojX0fxV0wzlInJ4YzuEuXg
u9GJBW9HQMlFyKQHS6HiAB7ibpz6fI+NE4shzZWtg4KHMjXtvcik9bdRpcQ1vK3R
1U9yHbharIATTDMjy47Cbrq66G5gXZAEIn5MSpsH5dJt+6qjyONy692SKCX3u6uq
z11Hp7Dlg8uLbpbsXe7Xjtm9VKr2Iss3RawdxeaLzTMopq3IUoLDEveuYKBUac1k
a/rO62CXoE+afIQ5roULTZDEAZmde7OPVsoQrMHz7gjQ791JWIur3sJQkO9Zlqbj
UCFMPJ3AatCAcphBQwHTIPRQi3GCahZPMjS06Pg80pan3oN8BnrY2Ru4W9NdxSo9
LJXyXZEUVlOaTuC5opzYjKqbMgxPmw7WfC1D28eHGeS0wtuqEXqWIJcDleQ6R7S+
7qpJ2AY10Ge75eZIgQ0HrwyfROevjdYi/2U3PyqgLoI3in2y19qrnK8BRBFskFZT
G8NR+hS+5PHvoC2TbaQsUt9ZFK3d+xqeXrV0dyVlHiY9S2T6pkOsO9jPF0jDCTqA
ySW4Ji3n+snVDrYsm+YvoUOUrtIMenFi7q0NjBVE4qLwWZtg4sp1EPYU/N8Y3RQG
bSxuT9VkNfHUO71XAOQDv5K31x2JNBuJnI7aOY/JHGwKvYh31RG/T+MbibeqPGzo
Bjzlm3U1LmJCymrCp7Ef8n2IC65GiA2Ga4see5WnARuGMpVtX8DrdMWmInckKLRk
ma5NBZ0sxlgDMP2ksg3eLxY7DYp73Te0CqxWv5SKo1GTS/wMq6jyfyO5sPeFS6YS
J8cW1WgL03EKzmc1mLOhyKTHNjAw8yz4xrkN1QvozPDxlNI/T4s6MmYwE/Koo/Y9
PeHX8s7XaMiFZtkaZJw9na8mFjmxS4wRuYOV00dPwzw/xcVooFs58V63JvHaOQpd
IlfLnmfU7t++Dd5wYhOHBqFW0n9HZutY8AMb3uFT6mGUe/oukK6l2KJPnwczkogc
lMBi71wZr4ziMkL41ITBu435Qsj+mITveWNNo9xRF919PaIaGvxtvuiKZaI0guQF
aVte3JC6bIrwD/FK6v2jDWSqyn9TEsG8Akih4l8Tq1W66IAERftOnO2eQcgrY0XL
mtrHYBTkH8kDJaoSw52Jcz11rC0T8VaYoGQH8jeX/pxjIep+xkr+tPuAluIWWwAs
gsdHgOLhwmkWjOeNQz4GMLUrPtwSpdSiYSRoFl/l9uuisu7BC3BFMDFmTJPjxgpN
z2zoAqbRrqglgctaJZg93uJjGbDQL9lMxM7boOBfqEeID7xuRppwFJKWuvHlKpFx
U+4L+fjU57OCF9qc6zN8bQ1VtiNedjB4hTJuXexiHmZN6HomAKMevQ1C0eVOLDXQ
JC9d7QZfsZp0ezxLWYFGDwvv9T9BhCQ8EnAzQibK0xIWknd/EwanFHj6IO8WsjBA
nFf5xIpAuhQWQO93Ochw+p5lhXj03efH0VHZo3AvEg1JGgYnttFDAg9OXt1I0T1m
QGA3Dxfniuxh2kuJYyxQt9yICpuHtTvJez8lH60MQJtT1v3CU5MxoAOUqyR2tGR4
JffaW2FHGmh/H1Vo9nyUtpE8sLCh1rBCiQJwfa0DSwe4jDV5iBaqSRjkd7P1OMnx
knf7o6dgPJxYcjD5DGg9kK8xuR9wLs8PUKr5bQtI2pX5AZrpmwHoSBsqsqKh4Xmf
5qXMwiHk9qRNFJf98BI8+qYdoAt67sWbJ6X36Z1WjHJ3S3e9yEPULrlEKD3l0+KV
OGBFlkVUttK3b2SylCZYgMWjVWSmAwLEaJmqjJx0VxSPrzn6sDRoLWC+7f2qA7J3
QH6uC/KajRqK+fqxlsfPG+TDJBUOeM3fgC1Cimk/tF7q8IJpSsXDI6hjZdWQBRmE
aUjMpFDdJmYP4yzflS2VxUBgnNj/OYHUT1rAFYyjb4P/ummrlBMq4zklMkuoJTWX
tptCHcaaF2zNuFT2Bg9FbG0wJkq8U2/u+gzJS1fHFmZuRnG/BKJO3oJHOe1VEHU6
YnUOlvpoopGf3MHKxf5aPeOWmXKhtmLjWBi30KlL8heck3s4qP4lOSW8EHcUtThQ
ipqAZhaeV/TYajmuYP6lia24UzP2hlyOLLDAczAhAefiUk3owraL5gYy+hZZRUSE
gVCtT/ed8kzYz+DT0MBgOFDDBKn0GQyYyyKT2R+GzEr9iyv6stQrbxE4tAs8gbgP
SO3SCgj3lXN80PglS/HjNIf3nVY41jIJwnNg/I6qO0r36HTOICp0c61sp2c4HURS
OdKPuB9fy0/Rq4BltU3RZOuQIOksPASzPD4ka/9gPBciWwzHFGe/qdyr9R8fbJF4
Dr9uFA0AicoHjncM25xe6/IGnid3bW/9hMhMHRZeeBbSx/Nsd3ESZDA1lJKJYynK
MzMm+tnAGjhaeQBtlUUHY+bd4ywUv28rR6i6ItpclZx0WPmOSGxcFwuZ8r56YYgt
BHTWzfkp8pPkUkogOSj33nuIt9qB0vUfG1ck/Bgz2xvdUiS8SC+n6SGjl4hrdKdO
pI5Daz2lBNz4r+rlfAw+hAi8nxD5n6ZROVgTc58s6alHENPIDGHMs2qWFyVfDPZT
knNK3Y52AUHbPRD3jVLiDL2ux9qddMHXWCblvDdPKOCpAki8EgGgAhkKqciufCnw
DRxZz7mozersEuesgAlrsrcEZTmQCsdE4RopUGv8sOCIuc0G7p63uFErKhIuslUY
mvsTDkQIBNmRg7B4IoPov+TTiyLVSoNL8rrKt+w7osztxurgiKIdTszbcyuc4SfC
faSSSY8+EKUevod5/hV4jeyzShva5i3o4t5DhX7Re45fihpNJVnhBC3N5iFrFmTx
2+6KXHC+s3fGPI/TNgQscwL5nYd3HMyEK1bowEVsBjobZxEozb5chdvdDeW/6Y8d
W8vqTl2H403DMA/3QI4shJXompIcZOC5FrDNoWxIfzsBogCwsdDmyqC07iKgD4iD
6+NDu7ScZ4yctfjhldunjdpDry1CutOisnqfYNSllkxaAbUNXaj2scPZijTrWHIL
ecw+U3TEvVAktAPOrAAGiRonKjzuFKk28ugAzmYAWESQYRBSFCIawVrMCruQ/46b
69qrhvhVEH2dyWTP/CqoyWnpla795non/LQRGJweD5H+5robnNK3GNh02quQAEzQ
eJChglRlkq68WPhsPR2Krh0oEcvlj5anve9xG/1+YTj607iPXUoSgjcBPRMOfyEG
uEWL8kle2SqwYofDFa1Dvfz25QmQqvxblW+l6NojeWQUIWBwsv6LAholvv/BBs7a
VssMgi0uqNgm9gFiogMzSiH/S+EzCuzlsXuQ7yzVWTkon6BmXez+cZbcmTWdfVpQ
W23SXPc3AnZaFJ8YbXAMuuAm5+rBazywBfFof4I8SUklThOnA0T4WmUM8odTard3
MWFaY10gTXnSDVle9mJhY+wurLTYYIP0ypwy7Gd7XBiX6844o+Rse1TI9ij3Ocnx
5gnGo2uA7lvV2KI2ogzjOKVIfWV8xGS8E4XIDPXR7q5ql+fKsDstQVzbqHVusQzR
CBTXHyAgyFsrDaZJi6JjFr3SDDfeU8wWRUMn6qtfMuEdtuWPy78DjhpMZEpgRsWj
eN/LGz1VbMqep8VMyY2b2KWeUDYnnn9IEwTH/3SlwUadTqamE1eUuw2BeH/CSiFh
iCQH+S4flQVQ/8Pj0yp1Jved2yTik5XvIrhjkCDQlqNSHhjD9OWjfoSQed1qA6LZ
h3CG1BQ0o22dgG3nb/5vN/KptDypEy3HcQdVCiWXfDtxAzOb5T1RCcS1jGpCKw5b
MsKGHbmW54DEnL9RdUdCl4VrhtdSLeNboLWchGCSVlOrKSe5VS8Mg0rkQUKz+Ct2
JpOK4ZhbaCant0kJ0jFY7VKUyBGlLG/x7IhPvgV1pEDFWLry8pc4cSby8ujxWRlI
KDB1tDZBwmdGnNqQixfpC8OWGeTLPHmryDnoc2odsBe7CX4X1yC7Xsnezt+I9aXg
O6032Cja4VAOgBCLAkzAL5EpnSYcsNggN9pkoVlDWIImxuAtaMUPZ5FYReCS0xPz
vFiVj85zeVni47YUZYyy5jEgRdXgSSdxpnn252Exjm+EFMz7X+80F9D60OdI782u
UfZiCObY0GyKoJFXy6lu/vAIxv+RlmZT42mSJH5FyNq7JSBdb0+tEVof2FzS0LR5
RMNwltpiAMFm8XQSkCAChXYWkaip9hgUutmfULyElGJzb7bIRG2Zlle63T1ZRRB/
1smbXgQyKqWw9PDZGzhO4+ONHx9pqJBf/0GePeYzWS0TCQAEudHyp2voHDVdD4l+
QiSgyMlnVhJJrImFi1XJoJ2bxKeY2RAKgNaM/iyW6v6Djffux/zOUVvuZMDHitep
+6xk/KYIq6XcuKMNycSFFpdPSqxY5UBuJ5zXoZFbY4R5wRIN/hHmKr4zD5f/4jY3
dmtCifFiEkD5piJ/B9krfzddQysq8lPF8zhcjpOUbCDiYS7C74x+9vyDbDin4ThY
gcBGaUxU6LJ+r8OzF8YC858f3Gt/8o2apJNWF47xFnneVpAApKpHhjeEREYFSA0A
0JemXEmurPES0gLILL53G14ZOf/hBrHn23+JPHnN0faUGgOQq+BzYemDz/DRyeqi
Df1fqqUy6m7vkPRyfvp/mQdAKRW8cGwyt1Nlomu8Wuofy5DJHEpjW6ascu+pnssP
nQGSGSy2Un1tmUPJcql19vJjtjoHk0wkjT87C13eYIMLMDalF8mG1XDfLvB5mtk1
GQ/gttlYtvWC3xibXxHLaafIHSFYi0jpgmyp/q9TzEvmBr3DRusyMhP320Rr4842
SL4/A3IrDpVGu73ZRqQWjyiOOt5ztaZVw5gGdnivlj9nF92uQ+iMFAwxboCZffv1
wY6gWtj9VOtEUv9OR+jaQhLJpGcCOQrFuaN0Yk8WgBNLI+skIyNWFaZQ6CHJAKK7
N86aW+CqHOtfODLmWEuf9L6oHXfS8BGlXKSicbXP1WK7EXKmQKhd6q2ExCZnjJRG
n3wfeihepjzSNoBaOcMi2os3mWonh4wfBK1dm5ZFZWpS8wb2VWWkt5hY0oYoTlPe
/KldVCglEyybY6cPT6sIXUUDIqTpsStLnKm0HMUU2QHaDqY/SsdUziLi/jze+gHs
oSTaJjLg0LEqW6U3FngtpXGjCzX+jxH1+tPNxdAoT3SL0S2RRCmzE/N7sz6EPlwZ
pc6LVD5n1f6dbhyDMgLKQgDAZr/shlI5tagOyqgedopjJE+fXqtf9TXQbOU4eb4N
ICtq4cmy1LGnTBo2ZtD4QDLe8/+trFEedVwiWyIkiQxOLfcgXr6A0diU/4x10+QP
vJoEyFF+ZeBT4OHPQF5+2CsaPd7FrCyeKOid4GAszt2UJ964p/H4L5d0W/YzE6wI
4Ut5divmU4vZq4hQVoHXOepdp86FpYXb4CP+VxtsgX3cLSqsIyVl/OKPWW4stkLS
Jn8UvY335gM++TzUhL7AnodbRIoqv2rOtjNMLyJoSN8ELDyKlYJDvgbXla6u8llI
MVOQzrvWlBWl5TaGtSAXpQCjQPC6EHamJyiUDhpGroUKLLHeMMO0MjXNcm6zrEy7
AGcSamgkpWImkHfds5O9RUt7u7MiyrjeKxnaRVzETNFUXw9yaI2dexSQU9wanU1M
tB8uIrX84u8qoDqXHKguxCdAdWTetAzZhFxI/n0bYFn0809ztYqwOjijgWcU0TXV
3fGV/LxoSVMg158ONDPZ5a9s0rIIuI6gjxwPi3NPcZmXihbBrhg+3ivwr2P2HFoe
8KVU/Kv+FaII+lpPK8Gk1vAb3DH1jHtmy0Fsjc6yKohX8he8HAyk0B16ZXjeDT6U
z25ZErXatBgfDNc1+RYxComwNt+vSowKQBJ10LNuqHYXuNJ3dEOoAGhA3mwq4s8Z
C4HuntRzOQ9HQ+6vnS8hTPkUjWRTeM25akciqwyh16vMBfTEYfb2oR4F04jdFoB7
i6fxq8Lfl7u3CNhk4kOOKf51TiwNzxrhTKvg+4vyPzLRVdo8hwjpSWPfk8yyBF4R
tVEudEsNmd2VmO0nmOtFzqwIRCtWJ0A0KcBLYQEHRNs99yOzYLxvYz4MFHcgex/P
kK2TMqz4+hRn68r9pf/PaK9EJh/ZwHU9RAtW/6Fmrpz0SWnZDNPVjMRTeGdoMl/k
1JR1BpSQ1oQlpY0WVlHNHOdT3e1oltVEx4uv4w6S8wZFID3XjAi9qNX7Yxw63pzw
upaNLrxih3VQoaXDld+yER0eTjMUqW7jEmLZ+9rI9+QTH5dIvbWdfCG4DJJsvQSR
xKOaZG+tO+iDaIyh0QZVobtSZGxJ9Y3hHn59xnWRTxL0tx8wJAFu2fO/k+kwgDuA
PJggs8oAbIPeAy9O250ivaaaKfnZ8Yzp/9mq5Gc/c3hUNWLo18H+DYkwPO0XMfB8
jlnfsqe9GxsAXlYgXH6CtckaXh6oyK4N5a91A7YGyU43QFbV7ZSLa7Fx1uDKPF2Y
EkUepF3YaVGwv3I72yEwnRsHFXWpLPVso7KcxSnz4oNWWiT3GJLZVmJVZUIc/5Va
LLjX+XU7EzzzF0+GN/Ni4yaIdjy2Xx5Mtk68BYRgufZFxGziWo9cOiM/0NXGyLKd
RZZjLaKRyh6LC4t+6r3AYDPm8eiuetw9uiWEEJsRgYMm4K5ON1TjOph/9cnYHCA+
Sm44Wd842iSjKcgCGE5JkUvZI5uXpAgVQCBAFJFT45H9RHigBm1IPhjp6r9OdK08
fq2r/t02MsNXobxP0QDDbK901NbrvQiI18aGIgsSKT7pCSoXUIUg/Qcluc7K1Rr6
xAEQEyIoCdDI9AVwwzO7GDmYm+htBAkK4vPt5GYy1rBU1SY8iqI9vrm99xWRH8qj
V2PDAskNxxWww1Srf+4x6JC6bBck9TCDj5jhiDFHTmVe+e/sSjOUHqY63RKFTJRF
XpxyTrRpyj26nk6wOoomO983r8MwCuAeXbq9WZ4J0WmLELgr7OsnRG5WJcdtdxvW
nzeSfe/9A0+PlnFpRBePPBMY10c/v/BBLYCJsFscQL+hms5q/LABAZpL2BlW4lFD
EwgSNvA7ZY+BBRXzlVTdQ4gwXXx9bA9V4hLDrfLyD3qE996iOc9n5TZ0iD7QIaSk
gpKVfDJDAHK0FDWxGhuHnRYCShrFuuR6VKu5IkhMaYpgj3HzWnB5NPpNIl86VMQs
hlD4skcbKaJaMYmfVXUW6rlCd5T6SWEaHUR+IYduL+NDoYlpbnkpliiDWNy+JY+t
mgahfe8n7Psfrqf6L3baD/LpraEulJzEC297MXFKn2+GNoQBIEyLYAiGF+jyU0cr
ZzT88ejtPIS2yxbcOZLH/6t4/nG38z8GhxMvHG3URIgb7GDizcWJKLpEJ/1BArBZ
jHGeox1g61JmW8WkDnOtHFOTbU4c3zippynS3LShEnJIdf5f00y8mhNS2EmjQbKt
J0rR+mX+CVgW8kPDA/WDMWk1GfKFKuAV81sdaFtTNo7Df6gMTypDKpa8ALDf4de2
y8KeD06MrpGgWYbTm2Xy3NIBgAUa05M7eTnquMFeLCcdampDpcNG82gjrYRFUMp6
SqCTEi8GgLCEZBY1eh61X4TvuVb/PdPi1ykFiNgk9snbAcIYY6ixpwGRNxb6AKyT
UwCFOzwfkABEcehEkvbuDRq39e7+/aJBDV6+PEL9rSc4OvTShzVhH1IXf1q9gJWV
zuXzLxsd2Ln0ULrQIa6fkddqFQlk97T/ZZJPLVedFpaySDAI6pjf234uQn+UJg0c
sltOmggFcXYNNdd7ONj90fEPw17jHSKQNTppltUojrgaptmvoYlZF8H+Gx2gCL5z
col2xBCz2BHjJNbaKm54HH+iwj8KxNren1830c4B6ddpF5T9myKtPgKFmwiLDw52
bj3yb/R5x+xZ4WQi4YjNGobjjDfgDPV1gVnv4Df++qf2CF0uMTb8WnmbKPT5PYkw
D8BuCyVB0w2/IhYyaGWcxheNUBkYapvdCdC1ruHE5Cc0HCaOu/zitZ4Rxm0TWicz
08nhmO+dVBXIETv/91HkyeTPh8fpGXRGRoSBhWDhvhen95KSV7hY8CUhd5LKj7Ns
st0USL/eTVxj7PX9CbzAkrA8H3Hn3ul8uqm5taAn3rrCjlC2cIEqStWbD3Uh6RgA
zaPSI3RxS2FPqQJMVpc5Eqyu1GRMIMk4kucfzfZuVjEpizDnzyULt5pwpkgB+F9m
fOjAclwi8Dsu0nZv1fjHdjpwbecVkxKum14LN3365qOl6/jfAto47oLRcOtZrCmx
3m1Aky0e0JiYEfg1hakhnkf8mT38fXLAz8cDO+0hhCjK4nTgO4FmgiNFzeyH48ME
g31ic4R2yIk7ufrtfX/s8VNqCmf5znpMkMebPt6AZzXl8tBUcS9cDy8cIj0bx4W4
81kprJdvJgfLPeeDIFk9X/WgwVtmYxgtQE9GR2kyS+4F5n7fz+qMwkZ1iGPPFHyi
s8pcNHhS99XqwFGh9qD3fAM+3M7GxSeDQ2F1gzh+zqlbKZ7YblkqqQqAYZSRoQtD
atWo3HpMpPtgAUTa4V2TmNSlxHWAT3b6SZC+Ctjiu5yevWHrkkUTWdmQK+awUhRP
OYZOneXgunGgkHUh9jETwkNvMlEkOVfVXzXqA7FX6/1xMQgNOFjZjkCRm7qDZsHc
MtW9eVCS1sVBQKhPSSp4B9BxXvaBqc367Hxe/Wzb80ogMUjt50li9ubpYnTdHudO
EftYqRWISREob8czFbJGtM5I/yAxlMkTDhj5siAUyCqxx7ESIfs94MeyXEzZdwoq
XEZ3Y7+Pu4+1LwWc2gEALjNOjvQqBwktnGTl8gTZV8S9g/iZ1pwWnr0M2A+JnV3L
6A1hh85wribYmm1tXrNUFpw6jtvCrsqnT2qkGIgbyyUAlir7091ATbAaXRyz2iIO
iuSxniR3SN5BEHbAfJQUHKtK3dXiC2ifLJpw29VL5nizNYO3ubbVNYeZRVZg4wfh
DxnYcVWKaKFD2RbbEKyhUbAQcHEb675/z+4MFU7dB4U6V1VFfNnwnZNixSj9wJo0
EuGvufVAQHuLcmx5G917/vSg3duUPzOwb0uO0exWt3QqCWlBSGvZl/Nsd0R0YW4E
FHq2V3Gq8HjIU3eMN+EfNyfK99i5w8rkZeasOhM4dQlBgDKeJvxuvmUnpjZ98XRa
7xp7CTrJWmfbKcyEwXQuuHlSgO4eGfTsb2VsQ85/ZEd8w7VZFE8EVay5alUzMGH5
XkgmzjE2kr/ySTichFDbSxxP6JmgRdaUhdN9SAN8k2Alg/nUkMAnpReHZygjOA4G
4kUbxkqH33Vhde47io/CpFF8MMLMsQ6XGPtAgeby4wtx5IzpM+fl7Xftknxgn0TM
0M0EDHdSnV8BrK48Nj5cgbVzWggW80+NqRrOoByNQWI308zBG9Zd+hYmgHH3duBM
2RmXO6pJlDThHYo3GI+zjfPMfLqCSckTnfIn5PuJfsxTNDfdHz4tnLHgvFOn2tiS
cYlWBCldimupHnxIAPQ3g6RJtOhyYFyb7jymjXqBQSQZ1li/yg/3PSk+5MGnYB7F
FFH0raU3wuHMCRE2yv6Jo8iI6lC8iqgIKmVCThStrcK53ADMC/zUrOM7sSRbB92p
P1mc2rwWum3okD6mHOZxU0EHc5P0UzROKIXYSr6bQ5Pr1ilqv7v0lkxRYft1E/kH
+pgpm5T+1np2Vzw23xp9OTMuFz3QUXzC5It+7tpdE3aem738XLXSdA5+PHC+F+99
HDWAJMXiX/yh3JQ5fP7kNZDy7ww/s7rrktp6VC22yffQH4hP4zUgyxepLn38Oqy4
pkl7oaVXL52DlZqFRszZLJXkUEXkNDxsS6RPd53ZBNhBwgdSLn+lKznrGS200ZbL
uIqNUFIJLo0PFl+IEQyMG5d5V96i9TXsc2TkDtKV9EcyOv+enELC77TFCzPW1NRY
ks2PC4Fm5RIdiLFjv2Cacexx6sok5+aMEznPR9fLVWr6KQuHHhdco72idW4Fj4vl
RmaZTLH2bwNM7QJogSjrSdeH6RXe/Q3EGm5t/Z8ly4sZ5H0dIG9EepOJ5Nm/LvwH
uXL85OzEOTsbie21uIaIK1SDUgVk7k5r1D8HI6Lv1lpt9NjFSmQ1WTCTvSstJ56f
++Zb6uJLQbq+lxygeUWzIOHH9LeWVuBWxFF7gBwHspuOjXnwPVBKOAZ6IBh6XEIZ
HUkNFuu9P6VXcuQLW6Hs5Lpgm848UruInMOT3OjVLiPebTM0/xJQgxh7ryvdjYlQ
4h9Zd0yzRoJz3mEPTlNVcJsupB7hAgnsyDjn0VthS2rjfmEDR5yXmzFnPu1IFeTx
XgimzDPi/DLefQZ+n6b90riTu+kaJQCHrxup1qfZrCsnPPIPwSPlVPzCM2u9Uepg
l9UnvDAQY6PcgPx+NdfPECCVJA0ArQpAIjV1G9RILijun23B5p6wBCgzKGd2zMzI
ChjsUscliTrp0F7f6OGtYJypZ19wTzP3D6rJkTEY7DsJk3u7Xq344EPOJ4p1GMDV
C3Z4/W4cpMyUbU7X7qgpRZ6f9hNAuujdoGc/9VjQr83I4wspcOzYz+jZlVmJ5Jv6
bMUfMIdh3fjVULQOCAoAJp6G7Z6LKVyEF8uDdidf6icWPTS4nfRkOeF+EGG1UPvy
W87ADc9UAqpPX4Q2+o4fu8iXqjkuKpZp9PaPQFG7McFSP6Gec+kDdvjWu/VfCLNZ
/SGxeOsPkqM+kaR6uGoc9yFt1PxXt5d+aQKQRC1FVCaBfYUqIKN0xid9WDwmzdNS
8sZjUZqC9x7ms2Wsf1/2imxzG3fUwliZffHRVb3FNFSdcmfYqawBzd1SQeBDX3ZH
94RpXW0Pw+Q6Rc0BUb9sA0yrQRY5GI4lPuNPTzLvdL1QO0NWsQdQdpMSJAMnVPcI
WklDSUo7DZm3ejKqPB9gSF40R01dTzrNZnQx5kxnP4666PlYQ99DIW2MQGRMPXhG
ZWXFjrhu/fsO5wa01O26tSfaZiE704P8HAZyyGCf+Uv4I+16E9hlftp7kWsXkEt9
IzE9smPqkh3eJ7duTmQEtbPWTj6JLBE7TWeLAlOu9PZUrb3LKY2utgWAvoFfnCBm
PxISzuTwlrgx6RyVouRXK5VcVluzfuzIP2fAI86F7oSxjXfT1il6V2XoIU2CWb4T
JOo7/SLWa8R6KA9WvX+eaCjLCtLHS0L1La1cCBzgC0CG1DoUBzD0veG6DIZwypp/
dZ/YZc7IFQMy5ra9/a7/+x0gxhYVW8Cfopnz7a4mShQ8m9dxLB8znt1LubujRW2S
s+T1TZ9K5cVAbLhdRK1xd/pqDahmOOneHcTAbILavPdW1gUnlqg1euFYVnzY8IkL
oXBLnbtGwDsd5P1jbxOHI4MYqbpum6WF7yKkKb6ks86ZEufKmEYXEorG9iG0s9gM
p+wbrICFpYAkSxwI2m/ZX/HJFFN25Ob5DydRivVMBx6qyWh2TnXJ/UmmBNKLrK6M
JjnZoOuQNDMBMqwGCpr4SWffrDpG9YS9ZCbg4sF8dsrFW4+js7YnzHSKYUDfpLQi
Pr9XG7t6D34RjWUsYccwsq8s6P7ZGMWbgfrf54niTXfyT5JAC9FJgGu5LqE0kuJQ
CSJoSzRozNJ8QFLy955FKIpfd/Z9KmXm3o1nOkPniD6pchYg1q3wkh55gvr0WWWZ
LJkMa7Mg9laM9OjdXhjY2un1CEc1uZBsvlc5dgnp8UMf1qksubuiRPIt/yxYVLDi
KRjk/DmKVcYcypBR0XAoQHcVTpBKQpI7Ky+vdkxObbx9Rq+3StBJS9zxLXrE5VPu
Q+sHV57gOJiKbqK9qNSmWeDDY4wFLJ5K18ybA0ClZjrJ9KEx1+60VGCgdhJLTkb7
vM0rcUFxZx2FAco6OlyHs/nhWL2lDIqmDN17ioReT4UDUJM8E0EA9/WPyr2zqWDt
IsAS4cRIeNyPeoWiVDAyVnzHYhXkLs6Z1OPrqhCwmN8pZ7RRPcgIQOCAUoF6hhd4
8PGJ7s6X4qPDO4yg3VOVkl1+xmLMeuSD6POLjCB3nROGHVlRiMtEHtnOXSZzzLpo
teIGGE7CQJwV4lHBNBiDxPpv8wAZ9SkfWvGIHN7i1Z3KdQOJj3eFv8XOido0TNZ9
IDdM1K1Z5ZtR10i9ezCvv/bASRmRpP1C9M9Zsi56xK0Ru0an4FSmU+ksYtjrZV2J
/YDUMyR78RgNpjALXIw8mJ2T24omBDEEOtSISNPfcDmJpWo1UxNluqqdQvYNJrSo
lXPiUQApc8lldDPdxTHvTx/Pngv0Er2YvC5ZSNUgRzSl4qRZIyVLr2lT5oYkPZDF
h7PUt4hyi1gHoSaUyQHfVr/tUwocxOnt7aj5xXMbKCC8mChkVEI6qxdIINRvaxAg
3yUMJ3Ym/rZAgwnG2q282EPb95JK24Sx4a/Q4zU6S1D7e2PKLiwYG8SLomIpTTYF
iYO1HMUNmli1KrwB1QzYYPmzC8P6/9z6PMcyp5H/2YKuiGiT9C/CwM/R2kY+RYKI
mG9Uh+LWCjgXb595MPo3Ib7rFvLKRDhOZiGpWJ1H0qvgfiQ2A4NQn3uLW4Sr3gfQ
XV5ILmeCrf9/FiE05XoulobHYaZr1s82B1c8lHchEpZoJKIo1fZL7e1v34r6ekL/
7f9soHDXt0RrG67TNqT264RcO71XbUpIEK0UZryPuMMQVR7t+nZ9AqIgyOv6CAtk
m/SQkosvsL+ocqIcMD+XpTk1K0hHIdGQaOJZOhX5q0dnZeIAuo4wcZnYXXFC6300
wNtp6M/fhOArBM3DooRlYQBMujNn1BkI3jiHL6RwfZheJTLrRlurzb0+lETlSJWq
/M9ZgKKe9Ikwul4TpFedOd3aHjK8P2muu25dXt2oqPiKyaOUwTfQWgEI6KnOLCTb
1vWX26iKFVnqw4nF6PYHovjCCnvEU7i++LEH1We/FfddUjmVuHuntZamxsby8TN+
dSR951pdjRZjcG+V9b2/l7bloc+gAqLg7duQ3dvDzFm66jjXBKovLVSo5vFo87xF
RVxd4cqJgPLdmNuHJMRvw9Aw3uWCf0rzAeYvXM7GGUW7juEp0F+jw8bTLcjhMaXS
q65AV7j3d/R9p45HiaG1uCa0swBjm5eHSILRklfBqhSEXutvrU6ggsOr0q31W+ZV
uzmQZnmL5LuTYSMtpvKNJFqd/xDo4aamzzPsFADQywrHtbKmyBnbvJGNplBWgtFI
LU+HWUYUUL0uCrSJ4k075f95b5VFhTWi2IszF5rr1Le8ca46PCJsvNkdQGBg6Zp4
gzzVlbRskF9Xdq7QCLYevZVWAjEMdTLLRFI+K7zONau7UancyYTTKwpGFrYWfrbw
awSsdCcAHO5SjqoC7JIIEHlWG/VdjUpFl3JX9xTjjSogZXrArvm68BBV6jtoc9Ez
AmVwU2TBuvuEL4BL7ymht3hxR8KX/in0mj3I07kDZOqmkF662kCI2AcGevPcDe5q
DVKwTngF+jwrMjCNqQbIfTkp+K3pAPUmo0pxsBf6+ewHLZHqhq4NNbeMA3HrYmv/
dJ66JLCfxTDwzV/O0kgdT+K2lMsjvQFS6gDOw87h79TF7lsVozcJ8vQu083czRmw
hhH0iBfQ/ekPP2Pm6v6cEAG2Km8yA9rg8QDCLp5rshO0qTRj58y3zVAgUvOV1aA5
FjgMTzR9YxglQxXGAA4H8/62cs7/xywsAmeAnsKI3XEw/BpGZmomfX/QvVu7lu6n
iAoNiI4wTAf9AF4D5RUYw94TPCuQvLiwEf9C+cSTAadSWtluZYBmikf4+/BC54li
nsGg99dhSgvZ3//xUoCbfsBvZR2jJeoqh4l3HOwUMSD+xON9VjZ1+2KoqGU+6HKU
YwwiZsqXB9qMtD8bVri1rAkEMOjghb40NPXfZfJVIT6bg2QhOhWIPzRQPEu2tZro
fiQyEVpqw/AzWEeEs7lbFrPpKA46z4GwDaGEHUUQ5eFIt7WaUbbjI52p5KOUnZFs
vPCdAo3yfmzIJ+nluOrycMtERAZ5iIO4Iu+2F72Ol70t1MJDWN0aZwb7zatNCZVG
u6Ukt+K0gl3v85tAuBE1dE7d1cddsVFxqFbVRGxfYtWazCGwzXQVQr/83vfKHYun
CZ08ArLCxt3NJvQQlj81EzjRzxmyYphbfkSRlX3qraA8tchS62I1ThSLMbpvtPPT
dL37tXvj0Cuz4skj4pyPMmXGSx47T7Dl3229ixuZENlvC/4+DnoC123hb5VaOHQK
l/ALX+ffuVu0BHmzZCe9MteOSmFmKEzgas7VFoQHFiULyrJn2JTkTBFveL2MPuU+
IYsrtZOYkKYhqFvLWBGmJKaLcpQOa8IRho6JJ038xdsDDyabXvNZqZnPCIRkVHVG
wDZwGHgEx1TwXOD9Netfn2xCMiWjVYJ/6wular4jK0+8qr5V106UVLf/tA186x0F
75OQul8pA47HJoXO6ztWKq8/QazQuft3Pe7cohnQPGlzUz5IH9Fj62Rdzza0OcpT
r+C9LUjcqASXgbmMvTLgjFKHINlZ9R7SzfkSpAYiVhssQw25jNciB03OHz0akymO
Okf4drnCX7xPwkmq8/DtRJMxwuZDogJXn/vaVYl2TXjfQYlv4JIbSJRS9kBt5RJf
YXCFqc+JFtnnVNr0v9AWL8lckiyaYMMyGLwHYfIx5RVXGzDKRTf84ffj8GskmgpT
7S4626vwbVHOJMwGmPUebPSIpB3m+w3M+/FVmzI3GnGTbTWmqyC6Mssmhcueqk86
L4Qr/lDdYhygTpEdEmxIcINfLR2JgPL7nvQ+uj3npMpmQdYd8Zpgo2lRv0VBVF0z
RTVcTa+WFl5E2v+eUvzpJtoQMAwFAqymRmql436TVcTvl3GdTo74ewyBeMMD7juF
GwQo85RJ83KS7AY1t2oa99c1p/qFhXW8Ed2ZVzafGG4oDR5ZW3AiCyEo9qBccJ65
Xse90/S7wD62soLznHcBH1hp+Ck9QhvLiK/kU+msTaqeB9shpSuV+u4HkBLBaMJX
/d7bZpS5LmQHBVTA/HidLO/E8XSuW4RoWUawX+J2Nnh4Erl5tV0hlcjW0VPfSR8Z
fy7prBQlg4rRb7XYKgDaxXolpwbM6HcbrRSZ7xT49zRznv6R4ivCi1I+etcZpokk
KEBCykhrk1/3IJgvDncFHEUVKF/Fo3TnY0Uvnh5grZv1/yshUeib1L/zkUc8IHdd
4+RxMsNeYPg/o86/R9duKnFF3Vx6sS3moiAapadvSQYwdodrnvRgejnjgqGmP49h
QDcfuoGAOWWDsBARlX/s1+CkKA1Ni1UBFfyjf0iCtfU5a/iw0zRVzVdQhUduMRAv
tnRwUB+NljGd2UvjcE9e1aptEPC7wn9Fdj+HFSAjL2fLSyEr6NtzWvVu9tnqJu0c
gYcPsQe9pUFKOIMiIKT/ivei0JCx1sfuziSvzsTXI9CZfUcm1jw49xyeRqpmLr1n
8ovNMtSWe1xn5nMohdlIDki0vMA0NaFBm35F3WCUJR4nYwhqtSP1dfajEKXmjuUH
2AbfivPJrHLqwZbHeraaaBrkrRMg6GuvSLTPet2pxZWUAdT5ynFUaC/fHzdH32eU
4WXQz5Wqcqkj+RYi/uKl7CJKqiG0iPrEEDtkO92pvoxfXpTo+vfqw8/GOjpLX+EY
T/A0FTBYomnbFwcHwYXGsGS1jcjPDpOGDGk4KG9ilZOQzPW+TG/kMF8MxXC2oJrV
o8r0FhcQwg/OPsCkry29nQpTB1ZF+PAnVK/FGggmcZ67wvkebAPLbsyykLWnD8E5
65a6ur0hD6hOVZ641D+JAdJTF5A+GKSMs8Ahozb0L7LTm6AQpvQ0z71c6usgCKWM
ciWT9D06IhaJgcTRoABF8Q/fK3KDAoSgYMql/HtLXenLrtApMsvSab2CCN+jmyh1
fpZqkqpq0SOJpe77R6gZg/MiKxc/azcsJHAeTEw1EAov6lfFQdyUJTDhE5IeDF9H
wGDQhDfuW9FuWzXlbppIJLvKPBTd8YD9o1IWieiI3IoZjIAzzTV1Bs+HvXOJt48q
WRKJNOgecFg7KrHaXsJnqVdHyg4snwUWaSe1k1zcRbQN4F9bWBVveP7PoSLlJNUo
5KIMLiIT074mA4bZak1Rgj/VcSNQi0IupqRF2l1OTgV0Jl7RouN6+MOsH/MfzZsk
CMNhAIlyr5Z3ZI/gKZRk0akjTC0aKUa8PtHRcSzI3bKwl1Z3eV5EiMomnBQWuumd
E+iiyYk0Zw6deQd5eFMNJPxOar0lVcu3NjL9Xmc9yMCIqtUmbBrfhZG/op2/zJ8G
cH6f4VhQ9Bb/J7wqGycZKhCxPpev0c4qWNxV/s/lslUCCCbe/6qbO6Ku6Px9LYwu
rri6NH71z6MZSc9Ln8S+JbrC3Jea0PWN29NgvRJJPtKvpZ9XVlQiMgHQPThNcNkG
w/PUdX/94O1J3RyZ3uhNarBdwvzWGjoVRn6DGzWBPep/gbvTPLwOjDaobaP6/2mO
63rum6wkE6HTJNEawoOV4LcKU5o9lsA6GLZtTpkRjp0Zxr+aIOwGzmtX+kJvUWpJ
h4bTsdeux/jVK++9/Ub6DFi+I5JsUAmVg151YsVK00mhde4ing/Q3tivlpDCwItH
UjrBJ8GjuUuaAibHdDnL7GSaQuQlOctOMDjuMF03SzXmIl79LT26NvWwO43sSLuQ
D6ceK+o0t2CRZJ8t6pmCl58buJ0rv+DEIqaX/eOucGK5uPOM2ihcseqQUHDARjcM
+lzBQqvGCXRYpw3bSbDcfqtmSZsMEw62v1aXARLhZt2Oy1Hzru5ISZKx4qLqkEn/
Ly1ER4vwIh+qVET3Jc8vjuNWfsEKOHYNV9ZtT1P1fi1DtEMLXHTE0K9YssZds7C6
uudQQnjYHo6APd1B5aKXT07/S8jNwHgTD89S9i4q6mqginaHtftJTyHEfvrE3ahS
ZdJxgTBb4xhhF8mXf9U/JvcB2KK91ONAXvB3BBqKKtf25Mm3yFF2ZjtQB35wh9CQ
Z1mGQ8dRYrV8oBwpFetGmGWonRP6NeOOY9XxFcdyNw4yJvGZoKklDM9elpUevNhv
nwa679oLA7jHMKDk9s2Z9Vwcx/cRwlTnfiUrQqWpZUd2JFG8Pec+AUveA9xibDxE
gewz1xvV3k950KCyOpm0l/0ny3AX8sl7qevNt1smCKcDOdZSylPs62hIdWmdNsx6
lmWnCS0ukCx+G+4WwSixXFqYxWg5O+moWrD5G9HMRh+wEez2CdJRVct8p+3oA4bx
SaEEoIDbmjZivE7HUehLDmGYyOYSk6XUKXes/KdgI1DnWWygaHJnYj66PDu+bbca
ZH5TyZrXROGzOBGGOgiaU1n47s/RCMapLqdvSRH326aXlirGRe9YE7sPGIGdrHVk
pgvc1dRrovXSpazz7PiCOB1cdJX2frKI0qB08OlrpjSs4akGb5dtjf/ZrtPZCZQO
1mJtDVtCojCdoWUIvdGceV0A+pR8/KI3X7pCISu3Y36XwQvbQQqqkTOv5FvtPu6W
OKvsdnLXx77X7lEFC+d96lNXVExTfHzREc32/AqYBvbns1ZmmgEPYNUGOimLY+hL
QHiUOYGG+ms1w13rTfd+6JTR+jmFfni/RHncoaRXoF5MxIYBNJDkiCmCpmbKu/AC
X44VHhkiP9j1v1dITWWhRxRQT6Rb7iET5aBvVSG3pHOP96DWJEYoc6TmgEOYcWIL
mOOvM4riCQWAWinT2CEd4Dz3pA4KlyNJZFTCZsmVT1pKizmKfshUgReq99IVZptx
Jel5n6pljKWTKIWvuZ7ZzfQMPVgjSxa5wgxrdQl4GoQmqwxL9I++lLOgui1q1U6v
7vsrbI08SjDX69tVIJsd0P+MTgddWs1dSNnl+Af57//fRN+aKCqM2ni0YfB0/c7t
ComCWK5iVYZKgl52QUVlIV8QOEPbHSrWjYkRAR1glIneAM80AZxwIzr/a2+uLxkB
3NFbYKTDqPZk/NBAH31d7EkT2FGPL15uFBNvRYOZMOdT9l2ML9Ehel/U30xvyxJD
Smw96JBZZXsfDzjK5CX9s0LFh8M52KZZS7MsTWfsOb3o30ZCnEmjU9bxkFh2Ymzu
2OKIqds6GOLiqmBTFgzypOryyc5xltPIzsOKoYIsnEnaLZoZhnVAdvNPWOFMGXzZ
PoKIjAIkskn2DK1Qjm75pt+0hU9ro1CTor5AVcU8nwCALMO976y8P4APbtluq9Q/
kdEdM9u5K+SW+aVO6Dp2EcQV8z0IP2Jz9pT00upAHdA951O0ABSN2SNG/TyTN11M
5U02NwIhUQuEyh0NoM6vHZsHmv4bQ6xFGLXPyIM/UGqtG48fndH81RzGEEgRNSYj
rU1k6mL7kS6WxOEW29jlpWFoqmARbSCiiTOyYGhngD5/MLXeK4KOmSCN3o+OllFy
auKfghoR1+daS7zPQS5pxB597+LhwGf9GdCvfkypiq3coZFJ4KWoviJk689mZ/ms
3fVCeNj3iB0kHleFbgDyjQBrDowhWF9EESXNba2jsDpIC5zQ1/3qyZo2gQxuzSZE
k/mjXpP1PL+XwdpBobxI0J0Soe4qxG4QOQ9NDkMe+k3SPGNioMSN3Y08hFOBZSC9
xm/VW6WGFN+oNoObXmxwXjOqnrtlVsmLDFyngRI/sg4EnozKLZ2LGit/1LTPdukg
MgUEC38ue4zTPfjQdtKjAl3jgCfT8zszJPYLulLc+5mewX0zHV89mchUuhgliu7Y
2iCRnDDCfcB5w1bLgIreS0qvNxdK/knqG19oqCPc9hKbzgL2K+9IyJ4RhjLhnKmj
IpuIxFiSopLJ7zqC4AAqXJvpoil7EM/nwbZUmqzDXPT0p6zdYtCEg8MApqFItUzU
YNsi+WGYcNe+wdIX9ScrgkQIr3GtVOKRr79xl441jDoTm3Ww9iAN/TTku1NfDMHP
gYyvpB7onZBm7Q9ihgKr8rqXvKzgQwgU08QX/sJW+c53GNlBkkPQBazB+WBt2oCA
zhiYURijkjWo+rQJo+k+BfyrMi146bKZbVgngM7zJQCRuSvpgoX357pHJSzb9z2M
+NpP9MRUCn+y4dvdNSSaXWTvmitthGZRiJKg5ArUQvgB7mbRc2vbF0eV4oJmwo6c
WpG1fQ7Ixo60/qNqAKpsmXj9vmB72ZigYCjZPnxy9xqqNKNTazxYp2ip+ymKyvx4
bcbWZBDfq/q7gwQhR2p8o9i5eiDodUA5lxhNVcx7m2TZA3Or/LYzpHjJHWQ2rh2B
l1A4+pqeEu4Ui40YiEzCTEvYlorip54EdqIYeRyFkN+idh0HlARG75GLNLoItMmC
BLi4UDPyZzjc3WBhh213nh+WXDatweL1QcymBWnNdWXtVLyCZb5NwnWbPJM7LbVc
wa0YZFY6g2Cd2xuolzmnl65+8L5F/3p1KflRyCN1bSGC8lCjpGmRhEkwDzDuqvJh
SVArqfo/cI2XD/Y+xcFPa6/a5ZPa4Is57QY4AF5bzxZ03WP0KFcwb18uIF/XgRRi
3zQQHIge58HHYGf4Xiqt5hXsPhv8B2wDqhTmkzr8h+FEwWtf7ouV2dbto2K81O33
mcK4+nUy8ZAvjBIJoSKFLPYiOCBiGsIdYusO9I49Yh2jFU2PyQBNzPU2sp9+aafR
mOF9SPy41Rll20sZa7bDhkOqcXT62no2yZTbh4HC+JVOEgrEfzQEMrfvGczR5HvI
72OwtqEHr2HxeLvv5zATbTJWl3w+KBGvV8BPP/Z5nNXxFOIwcepwvHhkXgMxM71P
F4EIVmkv4Sxbz3hRdPFYOTy21nVlCsEmgpBirtu/uzSSM7qEOQm2jhq3zwh84SSp
qFwaLjNAZSPgSSECbqopZcNPiqwykT+caqYQlKiR7Kbp4G9nQC33E+X7YJhn/p/+
MxM6nmrU5IfOi4ywLb7RwdOHHFJ3Bj6u4+OlgtQA6FdgbDfgB1GL+Uft8AvxcA/r
I8VYtdNX4OWjD+gOsfo/lzJ87xh6taU6825dwE08YL5G5kmps3S3ZxmMSk/15FZO
rT0jn4u4LwqyMe+zQsm3gXu6bJfvD4l1lXlE5iIEU3G+CnLRyIg4IcbKRkQ6/Xyb
MeP1C3Uxd3qtEQIDHbjWmndaA2dSZ8WrLA62dDR3+8bH0nlRhGdUe8CZdLQTJr2A
ukshZaN3QckTr4Cw/1BpyEi6w4rjg3SxlAdBzwLFAL9h64g6D3/tUjl6C52Pum5V
lJaebqNYCt2vpr3VNVB3ZXNwdBurM1QHKgkbkfkRb/9UTm58f81RJn6IF5fHHCPD
+2hwMNLtRQcZhrS1T9/xOj8ejBwMEsgnqJKiURihRLS5qHBkC0mMvIVhjWoRcceA
S2jKh7+JNfZ8lblWnFLCAAvB9dKu7TZIJdcrElLkvAiqgf1JOZ1J8IuV0RCK3sYp
HEzb6g1Kbvm/S2vhwW6xEYlgEVo2VU+zekJVjXQm3M6IEZVmqksxAHFX5OjShQ9K
35apc+Nqd+lwNAmO0qJr/vFN8Ndm+a+vlw4k8LhzKzpmwI/O+iDJ/Rrb9g2rbe4f
DcQwqy6taUtE+feokvKQPQvx9cDLWVicWYFu/nA5g92Fvlnw7A1EEI/CX01LXhPz
v6d317svLaEaMvpc0CSQJM4JHq10vp+vyItEe7oMTmCcmxPP+hpu39X5a9oY7gHS
jMk0uUvuG675Nogloa/4wC8VjBjivnmwBbQ7Ior76gSQ2ngcCE1Wr3Vb31i9OCUm
u5K1YWSX2vDbj3JTzG3B34ULwMHyZV/QnKWLTKqwV2GZUWAQTA9Gvlvguq74WwiJ
1sxJIEOfgN6ugv/4Mi/bbAqH//t9xQrf8reWr1WGJrTGqeHSSYGNBheyYCvPRz0g
zg2OiTdJxnFGvWDxnIJtP87Fj8lYNGOMf4sVKI2h4yhwtpSQdJ3NToKWpeP9KVUL
qaV69EHLSM8Rs+maZYw31yFc5g9yQ9BL1YMHLVU9jUNjbjPdPXgD5QpjyyaOEHup
wwkuTGzMJSjx0nCOlfzphufp83lxxCs5uaxH52VvoDAK5DY60kYa4ffaE0ebnw7r
qVX4hglTp6ztbTig0FFpTUi6w/vkswChQEvkCJD0uj0ALh9jf3eaDnoyylRIAEYC
Ft0mJTf1XopOpaPb/2etBWp06LYGY7gWn7+MjbbpQ41pk6v000FM/4ECqglS5ilR
nYjCNrpCO7Er6wh9o2ikOkJ/tFoSCI+D63Gv8c5pr2qHXAS/+zzzLBY4jdTWNGzf
vV3P8vLCxUeo9TrRtf6IXt5Cyph9/KxbdlibFovtp3ty2oeCHliBVOCrsIL0cgb1
xHMDJfOytZNIqYZtTZuLS7/vTAHFlOuZiWUBSRx2IPLTzY1SBWm0IgyKKet+plti
jcw5NLrDKp3ZDj5TlOe76xpqGxessZmJHyI2c6zr1cl3IbQF9xaNDXAZSwc5g8Kg
PhNaug+IAxYTlmpOayLK830TGjEHqf9f15TM5aHcq0+bDN/BW8hTN3nqdlhkdRhr
RUS8946slnB+InHCTSfwE28Bh+Hpoto2zdyCInOssDLkWOlqBPSPF3UO1w8WVR8k
Yk5OWOBm1yIwxdXKDZtS5p5EzORQEDlmySlKbopInqkVOGNloN/kkjveG67b3me9
P8i+3G+mbH7pqXgAFvStBBzN9J7r4V8eD4TwjFEe8visohfGzZ6GBJF9AUpWiy66
htGbEQHa/4dr65S9BEnzruin9HCW3Tx0LNqy5G4ufwNkxSvx+lDIu8GY9ngEzF8B
u2dKFghHy9efeDcyz7o39R8g6/NCgQ9+ibm/ED53GLJThUliNss/KlBir6SkC6BO
C+cWHrBvvOfA0OhlCOchquJhhzR0Mauob1gQxnxLjfLwgnK5Go4Zvy0XhLMo+1Cu
T1qQMoNjQh/aqe8GkV4qmiYlTpyoGvJMrcH/LmbShOe4ljROiBB4Cf9B36ihkep7
Sld/SuVhGl7+43pWPobUO8wu/u5IgQRUtOiL/TUpR0gOzyjkAffqy1otaGEtb+xR
GFu4ktQqlHracXJEmieW7TskTKY85UCt9kWwrVdsJZQDH0wnTJOci/1XLsN6rzbI
NGstuUDo8t5qIu5ZaucZp2Te2yG/RwvO6pJFIWm//FKBknt/wkB1Rs4vAUjY1nJc
ZaT6kPTzxHToZObSICTdhJyVpoiJK0KFOzBvJsnBCHvdihe/q5Y4D92gWC6Rxc0K
a2XHyyC6w0AHHf0QN05LOSQV5lkZupaa4VdQT0A2Fmaq+RhMnMNTyeNZCe3AhUOq
nT9WpiG7c2g1BhtkRsuAkqc71EMbtiBcyVoMfluWnD6Daedool2YEkRZy09bQxSh
Db5IdxXJZmZt9xocbV0/y9YcGJgpH4kGZBnI308jJNrHVfAdFsCS+eQpadKAjTmN
tABl7Xnfv9rZ1C4m1cJE1DVT1qczyl4fKEjY5Zl9sctrbX8UA+qak5s5MWZZXXAz
STz4U/OqFCvy9aX+45D1AJC4x3hhejwBRpDpDMdXmFpG58lQmRH24KX9A+2J3e3D
o0pWf0E11NaHfXvzJZOxpAf/2NYLbq6xUTfLcb3X/vC5miKYJUWU9f5+8q839Y7P
po4usduGJZGDdoCwq+ogBFTO0U1Gtni5aj88duiSBEXyoXg4eK5TXdCYPNB1Mwrk
2ePn/5Dd5Q9xloG3ALU/ezCPdU3ufhdqK+xq9w5HQMb0DRy+YM6r0VSWN7gWjX24
m/tA5DDT7K3egGfVkfL/rpQQUYBvFF8wXVkkz0EqjeL60ZhBqLC5uMsSXsN6jtN5
E8fPh5ajo4RWZQ8nPDjWrJ2/du/Xt5gncH7SGV0yh+uQUPO0y4KpjbPKf8q3LfDt
xLd3RhbmTE4R1SILtvvJfdahkIZueMWcl+ZwMS0kbKwzCY+MsXWuQc+vOYifJ1r1
fIxizoLf1nlqPr19n3kRj+1VoFMaAo0IqA8AyRkavrW3Fi+VnI/lEwtfNZjQvyaJ
j6sfU4HPI2JYLaWSwCHICrrl1SMYaf1AhBwHaPDCExeBBlGAXC0EWWb7UN53MPMS
3wzUerDjvRYf8Q2QMW9/Exv/uWZfaDe1TdqQ2tH1bTDZYUVDlkitVps6/csMqTug
Anqmkuco8mKdCG0nlx5C8+GCYnVpAzcQX14R2ywW015rMupYe2QxMV5Zd4NNXRx4
iUnY/ogzh9PcFSZPv2hwHOpT098z1pNry9tTYeg5NAgbPLCNiV3xgrjUfeR9u6/i
I/Yt55Z9ynd9gTWX3waMmB+HPt7SBY/d3iorcbJA/wac8nm+QtUZmQgL5g0j9Sc3
QJaVA2sBGE89VQidN1/wjunyPDw+aL/i1DLwWgOYrnAQLxLJtl1b2pVUxsvOyhhj
yNTp7o4ZJibvlPFMBvwNNt2HefAb/s5QFokYeOoFaeK9UF8NTKuy1ikq2s8s5Cwn
hHTd3evwJa4umzZCYZWnlGE2oBH4gOLYLDq7e4PDALeGtEbxjFRl6vY6ybL+Gnx7
wfu5AGYpH2TRIDX19k6LRRjfTfM4wCsPclWfoJN3NDOVjMRdcsUOnLZ8iijN3BxE
WVpvYH+4/3CZZHKaL6LgZSsr3s1HXxIAHsJtHFu9BdXmIrC7HQOnHG21CjD5GkmA
YvIpHI3CMF2Cf5z6WOID4fpmPcfwjK0xgDSbKY+tNGQEq3lFxEhHMPX0OUH5PGCz
mETm2CGlc4e4I+zc/0rFAYNuWLB+ELNUL8EB1PkCO3I7iXSZTdYuR1fysAKLeRbV
6edFVTSXoIERaqwTM9HLSocuiL605ult4ppT3rSpUXurbbrAvi2vgTOGOXE2NuLw
1pk2yMRQUvVMIgT5YAoMV+88UdsllpwmS1zOAWfHM+n78qPp22gxTGJXdL+VzQLy
IdrCVYQWM3V0rlH0MXECSSptPVHxUPYVH5H7KuRY2UrSyX6MlMDwaI3iTGIF9JOg
+2pt8MfRLkhEVCduaZ0loNlLUZemFSPctLM5WIJT+K/N/9fIjxrsR23ei0QfcRNc
oJX4nlAkGIHqsgUe+xn+CAjiHC+TArDbMzpXrpyKv3/JwwqAqsL46GCN979/TtBR
5a6D+X2g81m5sghmvXG0Kqg1Y83bPfOrovkHNMLdGT19Ty+Lw5bSdEQ+H2oAprVf
Syy5HbwM8Hh9VtO2517OpxtphYZjr+okmH38DtMr6xFso7Yt0AnllQRFkHwATjfc
qun4VNk0KIlXhIwt+7eE7xAGSrtrQzoXzzU+ZIKkbk52BNCuyAJMy+7JmWGGqfL4
bWVIH62ZraQLAW03Zf0XSoXQXXXlqF/OX+3dcFyzBXsNde67BEbd5baxCtPwQLcT
8HTTZqq22hxTAYNI9ojtibILX0WjzNrihx91W35H05zPSM3mtwuagevqdz4265IA
ju1rRWkj/TddgPyqPXV4ljBTnIqtukax5YGvJpD/p5sUHgLb41+lSLDT90XHXB3S
Icmk1wvXYnWIkBITCBK4cFdWJ7mSVfc4p3xnMxu+/2gHidY85qJnZ7b2WEKpquec
h+hmgA8mzcf2LtjT8WDC4xukydh+RetGLTzVCbkaUu/iul0GVrwYlY1C044t7pjN
Wm7en1hn4Xz5l0qJznOWYogSj/jaQhySfgYJEOSSoho2q95tREy7FpdJQbYCCtKa
I0VcfCBXl6WPnJEELBkOU2oPOb6unIRE25+PDhUsLKOl5WwtleFcqvvS30BnS7zu
7TM38JgA9OO/HR5q2N5dxA21SCDPD3WLKbQ+MUa8+6aXgAddD2k1BBzi37iRqRPW
FmMvnG0zvTBIGvfMSRxEnzAo5ie8wgsb7Vhj5PbVCSbPcIRDde+X0d4GsmFb+T0p
6SkF47jTVX2wWfThHohnXWJ7hNEW/Fix7fURseWE/ZU+Uy/5ebmoPe2OjlrGMtLI
X/mpaa38XDp/bO5AAFMjhthkGiVLnFLSOVeJZHc9K3F83n5OmXs/aqWMjwnC2riQ
hqtPETTCKYXUqTWPdCVac2lcidcvQuPMg5j5fkDcgjQ7DoZrRg6tcx+uJDvh6vxF
JQjZHeUgZzB1YT2CGmkAo/tsiFW8PyXy7xubRExx80DgC9TlAVgVARSVDEDVuCD/
vM9JXy50q0Y9YiLm5kR7K4fosTNqN/ei/xlS9P9VLCpIsFaixNuThFIjBKht+0t5
s2rRu1SQFwvhyAYfxhMfVZIOGbSco4mIAtXDZKVmwhx+iV0t+241KHN0e7hUfXI8
Eb0jexKzSk+FYP6ZTrStt+qAedrHA9FWcrrvNSCyfyumkZrhV/DQr7BBaHhTkAHR
lLoN3BdaxESxSi+5gMOdn7NE9CR61mW2Ys2foJjNo2vr2TV9Mr1w/VfqEn48uamZ
9fYRrsMSCP83hJ/8Kg13zXgJ6jgccpulIMWhisDBDDjjKNQaFjV07ZyYolTF5y/o
XGfoZHp4gtxx0BvXaFjJCfH7Y5S0EyoKPaXUy4GhPuYX4T7ebg9cilnJpJCG2dnw
DCvAf+H4aLMMzQl9CToPD/YgTyVz5q1uKH7CD28cIuqX1OHBU0BsbAYODCsLqitH
zDkXVOisa/kjiVKtidR07va06PfbzQUaRg2qVJWRbNORJBbn79kq3/Vc/nmcOHJx
WLeQx6e9xw5yNr+iaRq6GGhsi+HPRfSUyFOV8H6YmBZhmjm9YpzIGKRrxTnQx2dY
wM1LOQqNyGblWEICAguFBU4I2s2mDLk4GjwFLoLapE75TS4nkVFGaDojsayM407u
Pn9OXvsQCmzvCg7Kyu20dwtSzoeMXfB5Gi6g815325sM6LtlOVD/+h5RsP0J6dMs
zoEARVXhWeysaSKH/1UHu98cUnFLYQPYMwLvtTkL3fCHP19hb4mo+o8uSTbzCgku
TyOe5hVJ1uE2QaEExlVEkbFH8Kc6MNm7rGb9vZDjJACck79TQR3PHcGUlVo2tN6c
EkpwR49RDsx2NcWyc9/SkXsi0dUIRVcLYgriKNoU7zFSRc8MwYnzzUy6fRSjyjuB
iRAUkUQsGe/qWPMQmcWg6CPRmHmM9v/BsB72KZu0IlLHbJX5M+55o5jyQ+ksgq2P
yPsoF++1G9SqG+peTbPjLFmbia/3YZplIGFdIzjhf5jsRnJL7zRXWwHSg3jAf/Na
PhPZ+GLJmAb59+jywfHYQNmjHiiTY4GnrDmyi0zwUp26DezqPVotOIkb+rg7T1tH
zsfQpI0MqaaqbrojwjnqCbBWDvr4ZNGTofuZPi7FeWKW3U4EP2Cl+dVQawUOVEN9
YS7nyUPah1gVosS/1dgrgXyitkGVwlrNKhNrNxwq6JFbZ4eXrlCdEc+S07LVxjPb
Hpqx6u59GP4iCh7np2YnkcQ3oGqc6FE1yz3wjWdFL7D6/8oR/YhICWIdGS9hFSEe
qOd5930zIf2trgIobOHuGEsm4fAgs1pi1SzFRKGq5VB6sdqJWFtI298DRo+ziTg8
RRRLjzHYbZ+S34ySiBlOnAb5LMuGUmyzL3CKQFplNLPKn3ktDow633+KJ61jvRWP
lQTOfLbFYK0T55KSPdL72ny0/SrN21o2Lo6cfrRbwH1fQ+F0pZ5ScxE9ccZOpHYe
kI/+Jddlu8QCLJLKl1p5O0qFKRxIWw3+E6NasKF/8IKNU5XMocobi61+UNt1SRZr
ocPJl/yunCQPOV8jLv29GVwLkcVp72ezxJVSmS6uyw0UMsPKMIIrkne1MtC5IL8/
oeICci7A7pFAUZd+Q90pxkHADLVo+FnR+wAOX62XMlGc3iVXh8VL7rjC/gVlY7og
1Fh0MFwiiKDpjmSjYxwyoahPVQIrN0/rSzBikjWfYbxAfFF9hm/xfwf9dXDx9YDT
rCH5Fko/qz6O+DKrUnzMGWy7jvjm1MNv01okBzt6ljgsoZFZDmCr2bSYen4FzK8a
asycpxhQh9NvlTrKBcjL5J1m+D6Y477dssIuf/sCvpZL304v3Qfy7elgg7L+dpjX
/OWds0KdSXJ8/dGOlvxT9hakDgCvrdDc5Y185P0z8jbfvEfU532CGWyjIRGI2tMF
4ITE4wgFOxdT2njoEdH3J0XQ9S2FAsaLPvkc2CMGJ8HQ7qtDhR5KkEsq88Idy/RO
sL3VH3Jk6EzqUkIQQ6Vdn28mRNgPdwZLlHzlqZNvSZUFhWMeZzT4oWO38m4+elHa
lESGKJS7fvY9AhH4K4bCMm4S+jZRm6rhSsByviUuCEVwjLyVckN+zW7LUmtu5jIR
UrqpuMdAaQGWLQsqIsUoiD54vxqK58cE9Mu3lkVBwIHOxBORg+tUa+7zSkfRTIJw
bjNFdH4kyFsj44oEfFNcUHCH0snuY7HxpMxQrBLLmzw+t4mzW6BVRtX3kCliucfd
/SRQl+X6TYRTSdgoTKVliU01uZOl7i4bkDg+/8LtwXqUhBQgKMyLgyRpUGtm7vOs
fj6EHPqmQCG6VTE9bGOv2MG5q861OHQMpWQkvwENtTlynZBUXWdnhYURHj9KOiU/
VYmyBqdsIWy8eSIpSkWpdHkR5Ux7ADaf6gv3oiP1UvtS9aRAK2hEUozri0aQlvKd
DeYUNw1Z1zovDBJnjPmeRyjM1uq4B0Jmr/f8A174Go9M103YtzaVgtye9Dj6BLmr
gqKwFfhKxF4ivWiapColx6lzpdWaYEbP0rzXKH7sPPkecKzA7GoRlNJvIu0p6Gih
Av9p2331sFHwFa9XNVOy/1rFsw2HflkOiQ7paW6eAJBJpuYNRgqMHxceWU3vmWeR
IB5iciPJ4qdATbzHOGlMyrV/RAQVNUhB2xtFyr9wbKl8RijJDc+OHZLI5wYFQHYv
SOqNbSGCJ6ar+1ANama0lN2REzNC7/6nJz4sN60AQJKzmkGKYjeW+Zmuh1etgfyZ
IsLaN17odtlyAbmKlcTRBaIYgWjACdztmAAUjsY7OX26WNXjcEnx3pS1xb0VBjOv
2A4kqe28fvZclr7bKdcAq/HZUFbBNWmRcSYFUl1uZDQG1YTTvuLHt+tbaxkWRG4X
Sow7o1Ce1lcyUTfn/zgheNTYX4Cg01OJjjrFlKYsYj+/Ka0Sd/o3ehBaiVy4dtQm
U+UPBSZbXMhfcWWo7vz/4wCZFp1QDGJtgfH9b6m9xoakXyu0y0q4uHnUJ5olnxL4
3xP8gHSVKOFdKe8c8nYxqPw3nKCwc4hX+Amf7ZHxCD21++We25kCEyKyy8toMXa/
2an+ltC11odJ2grqIKAXtFKRMitQobFasU6a0/t84cDY2skPJCooXr8z1nYXXOOW
g4klQBtnJnyDviQLI2SGBrf7LBRF8vM+ssOzRQvG5Cl4ZdoM1+9uMJHnuAG4brzY
xC8pYJp2AzQ3cBIgFnnUfF9RYki9rY8JLTYuAxi2aDlOFxgQEqHK1/+ix0X7AWmr
LiU3618PE4ICNsQ2eMa/SUiY8wQSwCujMBm4MTyPT6706hBVGVf08vCD2PZNXsLd
gzcoQgysjrqCkYRmOkbi6CgC9r9tmy3l8dqSYPe/rL8/8ONdiAcd+D35jzY+21EB
Xhu2dEsd9nVR5y8eS+JEVPSHagHF19P/nPoev6U6q7N3on3t+qv7EpljYYF9Lvev
B7f4YUHQNJyfx9H+qY90tRRQDZtF+4VuJtxByIobCn8pKDtvcX/lUZToCv3UsDRP
w9DIC626RGuw+T75sDcOaxFTdelt86sv3iDqLQ/1g3eYtY7S5+K0WtoKAuhPlfcL
WeW9zfs2G90Png3MtGQOUXFfZJ8euqgjdL7LQApkeqd5Q6Drn6JHna9iHFMBmf+R
k9LdsKeJNetcdsKSnEacEQ0dzQx0z7lQLaCeuqGZSfRn758xSnuy7o1e2LR052nf
aYLqsrPN/IpsY6rA/a9eZwH8PLNK3WnaAw/3dNLHb8oNf5JfM0xQM9UgJgjmmCrY
MsEdo+0RZxCpZzGvn5sDWUpvQXSVbBrChG416oT4p9t3maFRq6oRzTWokW5tPgPH
ge130ac7baNoyQno94O+7p2vhjZBLthW+pqCuzz0aw4K3Rof3h00GD50fiWoAOKU
SSv4R3pyZzGSjQiILihuO6CaRNy8ZaxiPGfXi0Qda1YBNakXfMWWi0clN9eCe8pQ
h59sXsCxY7jtZfQ5e8V65yZd/lRTfvKtKePeyBWt4IXSRF3epTSHkY+dZ5xCDCr8
zsLHbtm64hqaouej3pPdCKVGnq0TMdrjKPH0+nvH8T1c6ObkVsujA5wrXTz+kF3+
o6PviKeKV+VvAT9rRHtm722Ky6XfFVWSfxB5Ps+KrC6wyJI9v8d1dXZ3lbkas8PW
x0oYTnMtrLhVCXXzDlVp9bYZMUbeYlVHWT6PT6mB5b8m5C2aumudl+K8Zr4zfRI6
lTnHcTteBrCTIkUDpr91BLXurE+zsk/GpTTmYNf22ghPtKAARNFFvsUChFfW2dKk
IQMW9Evr4uhMKRTwmKq7SUkf+qlNgzCEoPwd8Lo10xlZUAQlgxd2KBD6beTQ+UWH
zZ7Hrfprbm3hQJ5oKRRh+/RDhpCVwhwacEXzeIAzUi7FEN4O3XPXdSirk4VXVEm0
2nFGvJkk1VkvumA3f/thd7Zcm56HZJ/zN3gOAbnegTYLup0xYEWEJGBZzY75C7gn
1sRj0KQcGajxzMrMzzWa7jTXixLmrHjNNXuz5Y0z6FG3/IUeO+AEThHD/5e14ETh
qNI1DtCvUbdgNUNC7f/qgS1vJSlyuf2q0pnYQBShZ2gKnMZh9GwI/aFe3oazH2iY
m2woVa2f/J36z50BKqf3Wal7cZ98FNfhIZVdPUwQ4edz+rdmekO0xzZYwNJk9Fq/
w5OqDRSe6XjsjMwk+afEVfFvOnxX2ApT8DRDprDNrujwltBRCoITwfwFwQgdHdTB
dq582tYFj2Gs0+Dc4insL55EqvM5qC8dEZK2eK+IajDpQb/xQKOfPbzXZKh8Fs0F
3Ytr3qxUBlRdeG5OWrFfSx2SnbMMVq0vGSY4dNx8g+pCkOXSUoitbHw7ysKYUchf
FERLOyH2/YzcJYuiTQweNqgKDnvadqf7uU+gMOR0RI3/UmR/5QKK4lwCx/huieaQ
xq0dybTzX7k4EAknSYU3KqMH5DSMUErpwdQVdY5gPqol6NagkzgtjjigX3yq55lG
Fp2qQsXas8NyzfLgOqvzUJ4+6eaUCDKlb3hSjFEleaN/qDnHt5NySSc5QGrwgGtC
BvNPNIMwiJHmAvk41n02A36HzD3P3i16cYUcv4RAI/FC5EzGjQPHt/svw+/wCDlR
E1++fVvVuiIPamig2zOndlaoPPBTgeNiyy60X/13VLNHbq+8UA9C+1FTQtKn5nrD
o7TMAWk8EDojAMmafVaYFzE1nD6oSMbxxM+w10Hhb7SGPDfwvfN6JPjEqRCr4pTr
eVYyOIk3hyef0h+oi2sifBABeZMnZ9cVQGwbkIUygemHbBYmpdJVGBROFDOLC54y
zEcCWBryDbSRQvYqf+/yaoHwZVpahvMpCqa2aoojocmIl9GjlXLKwz/K/Di4RAWs
29AJyAJ+NxZdEGPuBzLdq3nzR8CDJEvfTzGWP8duzpoVWvKHbMWxdbkVE6S4JmXR
PFLSM3aY6TrndPPa8CoC7PWvQsEZAmepa6hnEj/wrm1V9Bwo4Lt/su1kRqjbhEq0
V+0IBvEURG1JFiNoKQ2uPDhrY5dAz6n/uQtgJcGm3srI01AjfaY0jRt8Sub3pZ9a
Rlztl2mBphQB/BuGVXY28klN53/7kg/E4aL8wafpxj9IIxKYvPFak0uY4nVnyRZr
kOpggvf6XiROrT7XrtOdv/HJGgn75G3xC3X0b1AYemSZFSyG0VkzbsQDZh5Ipd2B
4e/GK/IpAmSB53HGxSXg/r1Y7/Fi1ELBXmNFPupD5YU96yKzWFkYtWYo5d76s+ZH
/92bQWYVRD4vQn32nNXqcQw+U76jeT7uNjQyHAJ67mJJMzh+PS7mZzjp92JJMzWs
+Zt0T7wN3D8IP1mYZkzFMzV2ZzUDJOROAgZcMwBuR87lngXj73qVoKHq9ZKB0C22
mclmmzoXEa+tjDYuaB2Z5F5kYFMOKqyTyQGgwWrXNj+g5Ydl01YBW4ulH3O6Pvfg
9bjH7hhzWcUuGSqNTd5//GUQZU9eOvztkuMEWSP/KhA92EesUGHHgMyOPd2ysL/T
x1JFI05ySgvI4axGZFrVNh/ll61gU3M8ydRHl/XgNRS4EFu0uURJb+KQd8jof3sZ
0vRYqzmn9vCNY10IrQz8qnEiZqZP1dXrTAQULOqlWWCxqCT8lBz7ZjfbedjZLPZ4
+OZhMY1f/4WoiaRBikxWSynJ47gSOFVAtCYcwhua0WSHQFK09wama6iZPCpGkDOl
ya48Sc5BwSWwoJt14O+6Ufgzcy/ICqs8WjCjCESCmlaSCG+JopSkyIFCw8HuUYRq
p+9fA7K6Qv/ycmL9PTHk8C6QDHEQKDEfHnYmIRCagkj+gZ0JoTVHNnGCK0F+u2SB
SNFPc9XNUIOPHg1mNrvHr2hMgVnlFKr3PqqGVfnHS795CJ8HEx5n21QH2Ll6c0F4
z57vBuC2Z8YoEPRoj5sXh/AY/B8rss/kl3tMg/GolM5TUkrU1+qOmSZUGDgwIZNf
Eg/BCw/TwlNLjJtl+Hx2Jo/i+UcHrlitTqOUdpCbLVzuUAKT/4+/quD27X2FDcpd
Zu66CD4OfSJ9g9GvMeNTaAkMWmFuqisHMPaMUytNSqJPe35HsTa/JuMkQ/BQ/TEa
Yj2EJ5Ny0KxuQuaRJvNA2QBIzZg5MJCBX+5MkpVYAWd/B90OTRlODbV+1QO2fuVB
H7BcPwNwWisQ5vdvFovOQnJRM4gDqRKcfSoZLstRQzsSoVSrHe0v6bWZ/dNYnOEp
2u64HdE+HAhiNcoXU2N4/Mmd91FJHK8VEmiGwrhwEhE30kF6ruYoL6CLDTRAsK1O
a8V/vxDwAg3ab4kKb3TLT9XHiSShwGiSEMcaRJr1HjVA4vy9+pFiT1eul8hrEjrR
lFulewqpVhK+vuBWrL7rixpGuJCk4WbS5LmlQEU7WMkclLdFjbBR4rfZHfh/6NRk
GDGWBmGvFWcWijLhByqyYG7xrzEt0orVILqBskc1lXepU74ctJqYn9IlyjUD1B8Z
ryKUml39xTRwkzt0x0EomAK/1CkwesFj+Vki8qfng7leoUvkW0w52KoBp7sHPMI8
NeLLevmBLroqD++JBBq27IPpGbKzJ2CpIT1OlL1T/XUi+6NsSEISwM3aYz4R/P5W
I8bw6f6ttit00/YgC7LoWU3Ndzi/QirzclNo1r3jI9h2c+loQyN1gGEJk6mXg9lI
mSJu96R+bdpVYm0Dxe7ywwI3c5DooSYyKCwM35dE1Bu3SS19ezvRNT+G8Xhw1V2E
+RB+JCZxfLowUw1YDSP3qTQYGflhj8ifemzkIVqnMDeuyTUksNW/zSu76DIUlCCr
aDevS9neRL3P9e8WqVQgX9EB/1IYnC75KMCbWfvLWeJSHeSFoVQVINlzNYalp8E5
V5TvZ5fO7R/Zovcm3CgvdPydFMsyEmNexebQMjmJE6O6J6dphVxBOqXjBkVxIe+5
R38mz6+XB/sbBaKp3Yy4+cy9IvUashkIhi/E/5t/feR/MlzA8/y5Iu3G13s2LQrq
VuVSe6fVTrDTAcRMC3JMv/Tt6z65MwUii8+c/jpsjVCcoCZ1c2kX8al/i9YUw/63
7rq9lJDjb9e2mygJNS/UIoBZv/ZaquM1UHXGIZMkieM4+AWvZ1PlkjdlyFZn7ytx
kG4VsigZVkSuoHrmjk7fdmpZHQKOCiRHIaqQIg6JUygZp4IvlK88NW3idInpN+PU
4hadMZVWmm+/Gs8/V7H2xl37gSWYj6jdGRlFLVcxiOwVk5zrf3pR23DKmppYbJjI
OG04CPLWqPxisb6E9BjehBaMD4cw80PWu0NQ90pM/BDVLZNBrh4jqsG9avtbYbWk
QtsHaAQZGpr7Gv+Tqq8BGaJiYJpYvyaxqAYqVlsE+EitwXxV2Vg0laS9XnQFd7N8
QMA3yAsQjTb9M61sqv0YH8mZm9N+ZO9rxej/M8MA/XwcQtRJmdTHj1v7oNzISSBB
imOvtUztVq6z5gce6r/KEyl5wVUzwQ8gtMNaGtbIh8YW7XGd12HDVTWZAuPOHl5S
B36gd5DGWWyayRaZpHuRyil0uootRFieTRIrQt3RW3VrKhPQHo49oD4aSiTTy1Ss
p1LGGdf+CrJgEDHNaRAnGLS154btgujQn9mfCUof7xaFCcqr/RUmvQHldF+06IXA
rECWT5I1brcw30S9/kRzgjLsrUQGI6NMt6NyN/9usTNcL4UjFbLqItNd9yBmsvcy
qv/mKknSKNV7FOgY57BhTxtR3FBCasZXU/FGbjSqdh1ny1AhG4y9wawjpxBjQ93X
80yppQHpFtFaxnzHYQfY/NoytyQVvd0h116YUbo4Ek8TNamfk0htEQH0OxUNpecg
C43C++Ojot07pgLrFfIPdf2838M0CpPucBVw43bufi4qQX4rNqBlZKuhUKlpEEjT
WqocGGxI3xZhMG+Ua5zTs2irYM1RBOtYv8qiGtgwzucH1MVRbpfGLzGcG0OFM6rS
fdmBxMA1nD7rFxe0DuK1Acap//QK0M8s/5tMtL8m1Qi6/3TobyairlvzyKlnOrXZ
bGFRWr4CIVHrAh5Jfvd7KUFDGad4ww9fyVe1YnZsPP11itLNP3ByRpSezD1l48NX
C5VLiUyCvTZixQslVms9U0XIh7u46Y2GNg1mfN6xcNOyW53MS7aXn/7sr2AYOofo
IK6AgMXDUsEb9+XKgaqX5+r+J+NJVFdO1T54upZpObK4zjkuozXdZhROdIeYirNE
hLsLa32quJnC4Kp8Hd3RdcuFYA2tCzG6NhDDDTJIyQg+p+U9pUdWQbEUvapiVDue
c4P/u2k+sK0OKYC74td2q7DYaTZwYs0OMw04IyYQ99gRqFpsSUEmEqCVu3LyXXOY
pMFFdM5xLq+RZlvkN3KQwC+cDQeoptVdCj+J5B+AbEXuTcAU5OUu62j27QIM2Hcf
fDrCwA1Xpqf8AMflSu61A9NQmgy/9GzHhMIVO7/NfzuNywfDZl7XjpfaoUYGdt5F
7lOfhoJU0kZ12XFBRTtsoG5UvOixyKa+J7B9p0lJoFgaLkA/XRhU7ckZuV0fan17
bFNPM1T0loM4yR08I12U11OcfchjNLjlIQStXND9ywH2xyzy/uPWeVh8Kjbsj5Zn
CVftTcu0Vhwbg1aLMexD3zNk/9N0U+zP0Tdz15y5yY7WYTmfBcR/JscIhVwxI09Z
WtTuarpZax41opwZs+mc0Rm0CZYkB+A4hzD9VckCxzzMXJVYyTX2QY5fZ0Z0GLrD
zPCT5HGAFzlNk4YoqFQFcC/xqzFvBDT4iyUL9pVvfETDpMZmPkISocK+7LGo13mQ
xzRszMeMwr4yjThSu+v1aiJNTp7RxyZbaKQWckSqafbfoSPJI87YTQZm+6tih3BJ
+1SyeIKADGw9g6i3zRkx/kEVYZPo7dHEDYAaMedcUVP2PWVh0AAm34fctTU73YGu
i2Y+C/7K/hDoJC9viknbRmRQ7uoSHDq9mybw/HMJ6ParGt7+MS8aDMbcepZUleqf
H+6GZDU5Yrcl2Q0wWijp83a2pLDCTpOYHl8sbHHqJ0sf2jIOLO7RDGjGFM4/CaSQ
YVzneXILvgOuxXPX1W5RVIms0wyw9MKRQPY1XN4lsjRd/6FE2zJvWiluglJRTEhE
6RXOU30Hn8ei4yD5F1g3OQfkrIaIGjzTNSn5z3UWjSO+1/XHC8O33rbXOjNsDls6
NszOjJaYEAygh9gkGB6jIYb+1IgqsFUVR/ayfkKAvJThgy1AmOPR8l3EvjeNEN0J
0bzqeIAz7wRERhVCPwo4v+7pM9JZILvxqbKBhtgd6MBh0MQvaHrgV+1vXrBP+zJT
BTuTthnG6mtu4ihx7CQq2OIPRyaF2PE3IIX611AW70KyzPLzZ3VCr/KzIs5luTCS
Yv8AY0pzYQZBp0gxfY+zpR/yGtS6u0vct6XeFIZ4P/IqzirX6kQx22XgHi6XuHG5
oZoRk0ZMK3wpIGHim3dWwNSOva5aRZ+ItdBvUgwPwiSkFlN0Xf9uQmT7rLmj0XrC
UHh4UyTc0ZhKM6bq0glG8b3siX/gMq+TXUomYNW/eT3qet/cIDTOZWU7xYMhYtIR
pKhhFrpLmCQXp7+6gRBRkCqNapixZAEuwL5Q42zixtwA6+7WWqSXjxIzgD3kKciI
aOlUA9gEZ5HVDRc7SbWTshqmfSq+HJneN29h/lTiFt+Ntu0ZFIr8MdSOccS5uGcY
Hmm2ztBx46t41flKpBU8E7MHwPtec8PKUPYNBKdZ7i4jGva5xU4eHt8QItcI5MWh
AUHK924ZQJ3Nx8LjJcvXEnuGuKvmFMQZ7p8mklPmH/3c5f2DGrgvOm6BGXxlyaes
3G7okGWTQ0n/uxOVsXM6Kfpdrpco6tejMvZMnS0sr1GAVSn25LZPUD/XOcIpeW+D
NeQVAofz46zJxnmbwW8mYqVevpCO2H67K7/3ulZCPF5gzLp8Lj0CLl2C0ugOOvJs
I6tDxKIcPOLlN/74SAH7GNc86qN1Izr1irTeIebrDAny/0jms7HczgO7F2Qj+WYA
sqRTbWxQUxmMo82ADkgo6yqW0wUSwyvvCh2biw/par54zwXBZNjV3jW57j5dDxem
ouSH4Bb8uWjlbOTTrfLn7THwZP75kOesCXzt4erdBGVkJQcW5SnMchf1OIfc26CT
7exE0l3S2ArN5mRtbT2ITPwlFSjSobg3aqsnQLsoh8Icmc6b2p5K1ztobOqcJF+G
HRAtv++hoA5NlQwtUvjmoEUmUo/yZQO2eq6o9GzMPAabOkfpATkmj5Pd3ym+K5wM
4QV5WzllEGzWOOWs66WxA9wNtozsKyHoxBx9qmbIZ4DTcMqb2OHpFTnvWy/+DT17
5J4aoYMvbCiLVVX0Ed0UM405yrzCJWnhfg8apfn3EQyCLslx0zqFMjZmPoNvOLoo
NCvmmITK88p4vkKUhDvwdnBhT98R6yfH5rOorOgRFrC7ZLhUBjCGpM01c97y/n+g
6Jo1ikoJQY0hG5CZZtdmhA99vp/d17FiaQiAZqz0SP6mYb/gMdztaXoqwolJ4rzb
RKtzeMhcxvTG94LIgFRXcqhE7YYWf+0iq1aimfG7n7vsHbkk6hrQyMLwcBaaRLHU
uf70kalflkqLqEpPGevE/su15MymwQYc2aURTP1tbOYfoAd6ivWqFL2gncW6sGNT
WzWJLf8Yw+lHMK+A2CwwSEXiTYui6eM5biq4Ymsf18IzQYYtFgaVYhW7x76jPpeJ
vVBIQPe/o6AE5hBpXISJnzFvg/5OgQqanrcPCeR38QCmycJPESRhZYFhZ4FE7w2d
K4bnz/2TYqEvg6MNZTzCQR3f2mPX9+GdEB4KhWxVYrbyQu7duMUsKWJXe3mcUg/S
jDz6yiNAHjPrZPy88BaVAiy5beh8sh+8ojpPIX2O2l4w5M77lCkQuZooZHEK0kP7
fnUQKYRRFnCafezXk4EVBf9XEuVSSwCbys/N7tPP6baJ8GkaVsZfZlaMVKuoTbr4
C2aKXU1L27D+mQk1AZ7JgWBbJU+bCZs1CCKXfzJM5we09q1vDH5zKffQ6A6WIc6O
CeWXs1J/mC+mHm6HGS3Nzqode3yg2LOg+edi6qdWYpYiLkfdRkAzLYm3Y76YKEkc
B+q/4C+aeF1aMvIMPPb+Gn1gFdGW7VGFmDCD4DEuEPpGifsqlZGZBDwvQtn7CLOD
zTIoEMMyvAScq+kiqQwbi9nHNRZKi0slT142QCFD+hs9S3UFtukUBfzhvyiCX8sc
UnEddXRnfTgKld6ya+LiE+PWtTwOvI3OJetyuR6W7Y9P5X6oRpbl+q//OHnAWgQH
PWvwB2jJPqLrL33wAhaCmHE3zVyptOw3JhE+9vOkXzTOgSgiVS+vTM/my03QZuog
s8BrDyk9k1jZq6zIYEufLG3CA3ob2FmMzddN4uW+SLRZ5Loq+Z/br4Is6KOhrZd1
UuRkM+q0i/vaLd/uwQzkkMG2YBODT0dyzzBeHdxmcEEDOmBPhSRSVhDQew/GiZsE
i0BrD7T4vnnpDAH0qDTXUgBweDK15JEfBCzptgi+nT0Cr+GTJNKdVVBlAQvBWLU0
bDU4G5hTczKa5yWdl5BeOIntKYzdqxOmZqPM8eqlu9JaXW6jSkiBZyD60WT3beiz
cFqbXRkKCuRaO3mnwxf0pbseUg1jNCFhZjlUbUm7geBvUGj2gzIkmahFSxjNu/re
W6gduTHieWnqDVfQmDkJSSEk2c80f0KHJ0oyI2NsQlMA1s7s/BOrZt6Clbjai++L
d3//4aKDIttnmbGNjrKT9PMAZYMvTGiBoxaF+Bb/1hs0jRmf8IYkQCzWdtZG1ms0
xDVqlmJswlKsxfucF1b7iKwBfSaulA7cn+eenJBCCSF/bpvmepNc5LN3THUlFnqX
UsSW+e4Lnbhf9fmrk7vBOLdmzTRM/BPade7JADS6GJlAzdy+ek+9AqkDayqs5hey
YIuN+wZsMgRbrAzfQ4CI/oSgZa/ax1y0wtoAVKwArRIhQJ6BuYL64+pia3L06KMf
YgNsexSof/wyqIcpQ/W2eIExitr7wCpY77JCqGutLs21DQUEv2v2LGkYNXUQeqSA
kkEA4u7ZT4TwO1Ox3/286AUTZDa0yncct3uEQCcfsjapI9m/9BAjzwI9+BaHLkpT
00+BdnZb4vWa/z07zyAYxzJIbLh9BLhF1h5b9Vh2s2z87e9qw0rT0KSGCnj5Vu7a
5OcmOTMtGLfrHb4b24Ils3Io9+YIXKbNJ+t/4P73vVmSQjcrWJxAAdExnBHoB6WU
2ZxoGp4lzbLT+BsqQdqIy4IGpi151eUgboGgloptXBzWitwXonOD7kWFZerQZmBH
XJS9xCyUTn87SyvMee6SjbYTebN300/Bod4cD2HNtTLbyaHTXaQfb/lhfzxKVhmw
yVeP+/NmyOZGUnT2SM+qQ0HfE/5N/T1u1LuGq5elfmlq6i0ArFzZlCjj9Q4eqJFX
ErvuFlvbhBMnlBUokbQVcUSGlhN4RkuZni4WRfVFlsjdwls0cMaLDwgwOUHoEHRt
Jv8Q8n6e3qX+KgGB0CJFtX+cp/mTetjMLQVj4QlUJ/Ad96kk+qc/WHeDEdlUq4db
tMP4jN4eSb2TQqwTWkKrF8IrwvLqktO4ejo7ai5s5XkZJgxHZwnaQcjvu1C4Gcoc
vngj3GgkNccTEB9T1d8i5wf/hZfphpw8itQ0Ziku30R3f6vs/a/TBhKlcBnkQNvQ
aXcz977jIrKT8iH3SXOQf4a8JBrWjMfAZJ0dFB5EZ8ULegIeMXyvhdwoaTsBwDzV
JKz8RF9m+OrdZ1ivFfWl5LErexU9y4dzwyLqJrtAFKGjvafHErJHpCxq4mCoG+y4
RsamolXsquIOutnNSstyRUhMKop43SL3tVpS2HNya8SCAXbuKNLJ8whLwPmnlCpR
vvLO8FxYimgpWwwH27IorYoBiuVTAtdw/ZOLnlAcVQoMPVNVqnK9sz44LqR6VHiy
Q9HLzzAO/UQ/x2OCCijeNhwpABd+dSeFbZFXNdmE2AKHh+Pv+dbGTXjtdoMdqemS
EywnnhlyMiI8zgTbm5XaMU+XRTnN/70nucd2k1Ova8Qe6oReuzZvihnfzfd+dm+4
Od8P5Th1FFg5fmCfvwD9ZZoqkJyFeYUrVzVtP6EZo3Rlf6QwoZQShUfPQ5LM/9Vc
cUmQRTekA2EqJuETqcqb2C/sq/VPBh135r0Shkl4qPFesKvXLBzIVrA8GfUBRl0A
L68RXGYXANXJ0uAVJtHXExPWueSlRh+GnUqNRp1MZNNDDJC2rdumk0sqnG6+jXNC
DpTjcIea4HL51X1Q/keB6/eJmznlPLErOegUjBLLfRueYYZ1M572q+rCQnv5RuzR
7fTazVjbbKJFX1h28Ytk/bAWdmcWIrfYWvw2W1i7dHwJ03UkxKzrYZ4gbR8XlgT+
saoUF95SWI33KGuvV4Lge9tlSXc+kgQuPUquPkfGMCDQW/mFdKCNAbiF+n4K2Kjg
ejubS/jU0a0IK0MTRWkBi80iQe6eQGYBOk/L1XYfysur+8MlADxlsOccansAYTqa
rFGNPC7jQAsS20AUghUd3b7Nw63QICAzYOrSYLu8XQmhniNGfKJG0dp9yj4GKG7F
zB749TDGXVc4p+x4KDDQADEDvVTKM3JkTnXKtq6LLslx1k5MjcO0rghb+UQHgLwv
BTcJ1F8rqeXFTaFRfO3NHrq1oK4yb/dXYH8jHtzBwiAgwjDVHz76C6Vw3HRxjy/d
Q4E9hshbZ+NOocvfFIuOdpGPWEf6RcZ/wBlmS8//MD8Bf6SsB5SK9BDSZA3Wn8lC
DF/gCxwE2Tws6j6icZEvlG4QPe4SGq66SdseWBWwnNYHTOhWgFxIGcecK6ZU7VCa
thwUZnqgqLtVuzvBLChOwMHuqA6gdwREx6biIrkj28ZSkLJCHtkQrq+FjLRXbE7x
ThaMfWe4ZZ1SKMpvZHxbhNPSbYQaB4Z8I08KyvLknrSMD/+3LI5OpsNYSZlLYftQ
7ofMAFM4MzHJwfR0vIumHn1g6sjmIDJU0+K84n5T/VKvWeqqVZzj4uX/p/hqkNs5
HW4UZa4fPZIryk5SkK4eHL9ZqVZFjEIRkf2lqTYrdbBIf7JYzYUpTWPSBUvRJULh
7Ti9ppv5BfenKVOFSPqPoVEgoJisSBuVaq20CMYvQ84D0LizNJX5kmBuUwlTuO5K
6w8zhpkIkBnWV4WoulkTvHdGOffLQFA3TZcSGENd9dovHNlS2ytG8JMbl7e5PDBH
e81YptOaF6mWBqDq9Zrh5DdUvR4SKNvMH5NdR0Sh37tfoTc+uxfIfNHtX385pcG2
WejWZWoAGTAzd7tPEO4IvKZnZqMbKuYCzU6N1YR1iCHhNb0ZWrGoCc6XhgFQBboi
TOoaoX/PKSECl0JA5fhlLC5On12WpBmtrFMX+n3yPbo9VbsWihtMzfKTlA/Az6ct
RcWyOmLIEQqeOlJTOhRbiATFqS6TEEo3Xoz7ZreQDPjpaQ+8PsfNYffVBQpigHtF
IUK+l7w0746YYDA8U9Ux2PQzMKgmY/nHXVTvRGXZxDPPnFaJWnL/s1rzgeTDFYHf
htEkniiCfL9OHXXvaO6xbdt0jS1vQlYXnjQWA7Cr9C7q8PBOu1dqez/2PLB7qlfb
LVjm2C+C2uO+ukBT6DBkEEOJs4qtAD39DKXiVdSKGg/nE2ryXXOGXpvBJbXnx+Nt
IAnDTAItFo/sDLr3mN1GhuZ4elSkINXdByBn7Q9s1nXgXgLbUVarwvuYXv3MFFmU
CaHt5t7jWgsnpyRCrvMeoiEboifvLLps4wiE2Xulf+d8oo6bng9Uyx3PdqOKuxz/
52TxUOzv7Mnt5bg1jd/fm1TdtzmjF9cOORZKH3s7+BwtQzaSUCBJlR36k/6K17tp
6+OF7YA8t/lgmKsieJUKGxzzQbtAjhhSdZ6OtrTG6PE7EizreweRujj+R3b3dQVH
uHBYaU8AMpA8BoQCCqtTp+2Zk/YlpD44l7DaIPk4+9aRvVLY7nnp3h64c9nJ81Dx
Ok/QJdb8y6bobk5FxzvZbcbNm7XJEZdwxNci7LLe0+KFnYMgjeGvP1TrxH9uuqL6
e8MQQw7bEErbJbUSg9YSR+6kSX1Fbh9+40RoQUsxAapYQs4LpryvHfNNYzGhISBt
mxfuydavBR9Y+llUVWGnUNoeNf5+ESC0WucwvuGENZz7CpzIN28Ba3sKjTzLey0x
fkwMWZgu+syTllNzqWnyd3RzD+JPGLXL6PVzjg6mRtgqdBEkxRjyXkd5AnY2bQNX
sMDnPrS8/VRMYrbLCgsuofsg6gs/RmQEYnIhWCQXkU6bld5xcS5oHf0rMLQD7hrP
NqAVrH+A0/PZbS7wqANKrbWZRErjJiWy6AAf6ADnY8bHr3K6rlMUOU8aJooRKR+7
zPI52qxdQNV5Aq1/aQNYvsgz4emjoi9WDQbfCy34G1bJ0Hmr5wgHFllGj8M/66bu
WXL14fS2fC0Lo6AQqMngBrQ4tFrcHMbxaCz2X9lTovZaLtESqdooyk/VS1Awj0es
fVbaHt3VrPsmi+nUuiGYMAyndXlr/DHXhRPYcNYMpOLAMeN4GmFfUl7bgaWhpeia
HJb1x3DTjHXNhr+x7FGF+Lewbr1UlXiGDv+PRwzMwB1GB40SJabDE11TE5RhbAeV
JNeC/wZgMr4rbZ/g3dBc75yJ5UTvW0P/dtkHnIzqU12v9AHD7fr7++WGF0HokKY8
hglm2zoJBP381WqqDSeeql+sLqMbbtESSxr7lmgShEXQbrWfVuu8f7aDqj1RzovS
wiuac3XmNoXRZcYw4HRHIUfxYut9NUvRMur4/2GopgfRWqwYJeQHBxJiI87ALW2U
bg45JcgBt1RXzFMLDKpEGhybJ6yM4Slrb+weS7YlEPju3GYYLKUX0HvLOc3Ls6nu
oyMp1N0cebQb/ZanN8O/s76v23Yq35UBR1B9w6+fpbm3wFxymiOnOZgQEquRqLi/
L/xG/zdhz4afTrKByktUUo8dq4+UhAAT/olRRbOCJf6LQibe3q3jAd55fxZcYEFg
OZHBZS6IDeEYJ6/IpxafkO/uvEMgobbAhCYRWju5tN998vOl0++C5JCEY0a8wzpl
/aWCdyTe/He16Y0A1CVH/K8sJENKrhwIvG8TPn5fzUOrP5U6t3lifcUxU2jrdw5J
tADs66q0p9yJsg7CbkBsH2V4jp6dwuvyhU34BSCaKd6RsDTkK4Et7lbNrAilsxSZ
6wQY6joCnlZMMxo8czivEE+Bx0xJSszZLvSTHQnqbjTPQ/LCWxY5o1P69w3tW5bi
VTA08B7i1SZAkcEZpp87cWZbkSIYqusMkVfz04gC1D1ifqeW73jRPljPAruqdXtw
PT4Kd/wVNHCpa0mKJKRG35wJ4CoqO42vgGe4owG1OyRPHcF+9vC5RHkK2DLxrtpE
Vgg1CD865PgMSbSs9uSiLaBtbP5sumFdhWsAGwXUKt78RrcONnMmJPvaWkw0aAh/
AFStFafCMkojTRB5IymEAMlUKqEl06dlJt2VTM2GS0wVTk9XFIeTRpN1ksFkK5uE
gp2uWKSEZ8qlk5f3Cu1TBmVO62bS0np1JuX92wmC5VG90Coiwb4cYaRjyWn6TFXw
QV2X+0mhMLA13+ouaCEFE8yOqK2WgakfRFbkBuKpwu6tj2e+79XMZC5cCO85ybO0
yIJMCKiyThK5MeQEpzYsdBmN1fmkz+Ys/fJxN67CqK6QWI/8YLGNXnmFucFYA7NN
Fb0frTifZWEi+d5F4783U3LZ5L+DYLr7X1fskc8iguOkezX7tiM4F9E5BnGiiUcW
k9KLgzwZ+eJ7yuNd/UsBeTd2D4h1CuZuC7m1K8k+pJHMt7jRffMSobM3bSREloaL
FR7Se13zouMwZ7V5uppgIpI3XPFclF9Hhoyh/DqC/Rw3udRP3q5CaDXJWBsB+5fd
4NQMOmNJUmIIxryep80rI0ZfaVyQn7jBj5HCcIQBwH1ObL2RrakulG2neTjZzZ1e
tCBmtxNkh8X8g9YyctnCLrQ2dat4siMihEDh8DJ2CYTDBWDAEG32Yz+LGyPRtZjR
XeH2wlh0CUFGXNqqPfSluGqFlwZzzAl0r4w0mNVJagFJ3Jts6hpVqz4HPxWYsboF
zLaK4xT78jHhSl/b7z7gCAPMEfowfAmgj6hbY2GwUeh2s2d9uZJBPbXWLbM/0vqT
gLkt1asl/G1A3kAZ+TE60jIxzm2ABHjWW1AnfG4x3e7NIu0gwBL3mnItc6aY5R6D
kpgqskrdYSFajJaN94LbNgrmwE8QVUKXYXyMPwYubZIBEGSzEFM5WRa0BENpvUwe
DUEsVyj6M0uskbcldyDREmdi/LnfM38gD06RMSI0DzBrk0AAsj4Dcw4AVN7YXiyo
WHbewtM4fv+77HvcjY6M2RdU65JgMe6FA3teNMkxFCuw0J47j0dPaOchktU4a7zq
xlQ5mLe6eQwVA7gyDBY+yp72PR1j6FDJP0rlKJ6Zp+8sRCEs+i3PTKroFpyW4GCV
DERnHoigNQAGBWMuw9GhtKM+xWKklBpeymDAp/jh5k3TQxeZaEZpZlAtGJDbYImP
rYDLC5wlUGdl5fG8HBoSEt14S+jqSwkw9Rj51enuBfZzjKlhyCiFdq4RGFL6czO5
KmDSAeuYErpIkW1OEtcjiyO3qdMbbIPqJQ5bfiLjja6udPq3FjZPpx2aJCdccBsh
E8Ah+Q+FMgc6jV2uR+56tebvqCGySdN8CZ9CiNHJyFs0qqXIfOTQYZZi5ACouArS
d3rBqjMYG9iVTIR+jBdASi+1yWctFPKIi0yDH2AOL0K9YV3oAghrufZAm+Hj0/dY
M11XdRsCYGkDYUNS1WrEmNHiEFjxA8Xe6KhxychRJAlNXpo8mFhakD5JOEGKJf2N
3OUR/YwRsGxN58d8C54Xyzhb94EjaGaKhO35MbuMh6Oo+WDwMgVHeoDvhX1zl6bf
xh3hMD46jw41KbV0qAplatNorGoHw0JVXKoyQBRWTHBcXYJF3CKQKvgB5sfPzrXL
RHQjkBjy48YQgzc3t3+fk0lC26ZgFrkpnQ3kln2OU03lBDEtKfZidXOjh+LcXEZi
HVP9XK5fX2ocBRdzpwMR+lNAp+uP180fP3EFcmY/sc+7sxJR6NOvoJ2k53iUCpBY
0YsBPwaprNe5sH81krLHukj6rQqGVMl4Tm7SdYaKUnQIGx7NFDfhe0QPi1kjajmL
cOhpcQYWF2iMaJ+Kv6zM61gnz/xyYa0mn+trxu4ipT4sIhHOg8Yum8zpwuEpc8qo
C+f7iOav7NYyeSjFOBnXGGCyE6OOuK0rvWsLInzR04Y2B7LY9n+wvXfvWFHFPCw0
y8eQVoWwZPEKDp52aQDUwnlzN8dKNyaoNFmgcBJV2YaS9RBEpnW8R0G3LKxwlTnb
lMdliRRrkQ7nq0tipBLE1/meF3us/41JTJKMOUHKoi913qAhhzQ82Gg+iO/ywDbE
j2WCzYctcV2tebX05/QwY5+OtbN8Z1FbomovqLSFkh7SbhJ+jlgJ91spwPvoqloN
VnfHga9Z2oxKch5BSXmMQCeeT8NXZYaDH4Uj7EhHzIgNAs9XXquHutrz96pi07sH
zWyaCpsKgGDWAQAzwxeM6xtvc8a4fKvepwUsDDr2bFOoduSbuSIjAOCYAov53bfr
6HvA6EDRcQy5ElBXxdryCIxKPbzIVJ/lTuBS/fcNR8hkjtgN/GKh/hjBFJveKpAV
ZCWgCkDOcPcJPIOA44GvbqRks5Tj0DhxzridNFCF4RCMdzJyUX9VyHp5c7PdsWVe
BflIiaZPjxnRDuhdrQE8nDqUfIqheUwSt7s1yLfp2JJcLfvqrMdNo4dnjo6DSg55
OgBYjFtbTvomZtNptw0TM8u2Qv8r2mieq8MLDBrpNT3Y6pUhs+/8TMpR93QPNldG
7mrvHsEygpjdV8JkXhm/TQaJ4MokYFSYLq9Wcn/6exJIFbYJgtWO8SRz2y4KDegQ
bDS7Zb01OM1t2+o9YKAPk8qguMZ4YlHCjtCBnxcp3X6aronyXS44eNaemDXihvAj
5VELlvOOIQzcsoQ4Jw76K76CSbJwS/Ehr5+CV9OH/eto1ELqv9PLxsLjIVy2j1bG
9r/4sNd+OIFCoFaX4Ur/r9UW6lEsi2NH6Cu/vCIu/mZBq1JYkUhNLj7OwbsGXjx3
IHw6Nhc40fModJj7iukpNV/6LBRYD4gy38nHS4Hd3Vey7yfWC607n53y6z+Ovv2T
f2rXum33Bi0Q7ZYuz4m2BkaoB599g+UWQibU1diNAqXjwdL5NuDye6Padj9Opp/C
qb/6vn0hD+Sc8pjQtY4lYktrDE0g4wBIlUql7sJD3OBnbCf3bk0HROYIXNfA4GiU
yITCrPG/NkkPOqsxQTQafteMMEMguCz5SHErNk1WsaN3I4FS0VIPj1ruFhbToETo
lEmPjhA6VkRELlo3clBkkTtI16zxmE5JT9EG18Rw1QJ0gesycUpLC/7Nqk41yL+r
b18N/qKniTE5LJFhrLWP2Qgk7aFY6V7F2Kjwbu/RwF7TiI2I7NiCmwEBTspqElD9
3Cgl4Pwq+GfXzij10fKdHnqNR1ZHgLTY988rHH5RVtxTd8E+zYME4s9hONNWJZ39
QxJvS53VYBYaFWrahoSyAPtHOLJqNgGmlDppeCuT7CF9WEfs9EJfMApP0S6foca5
sHR6Z1bOX1RKyWBGbhUBuJYf0lVGSudlsQzi6sjQV4lekieK9h54fQCFm0BbQ8Xs
4145i3tkFWQugEhNM8CcDS4o2q4ENZclExbTbOUaL1IIAjlD7IrcO4TPePGjFDNj
iyJO4NJFjlbrRvc/3dawAD5A/tc4UnwRdm/256B+tTqXk64W7ovV6hwg1HdzxvVt
xsMKzazQEAEfA6UNlM2LBWpVCkRXEd7tMbr8AB8La9o35HfbGnPV1nCwC5OXcfQz
zjNW9dlDbsrIifTwJ8kHYuUa00WeKWcOV1smwHMIpHpDLqYRESmCgAwakoGXsJ+1
+wBmu/1qWLqe31D1iYuf2RBKEQYNtWmb1jNS8Gs2R+UK9Fo9z2WBb3tMx36Vr7Ed
OiJKyVHK29sPiQRs77bGyVtjTnL3yMay0tU3MDMjr73ywyV/ymdblGogOQrTlsln
OOanP5mO7sfBnbiXfbhd/Qg0uHxavmxR4qaJU8ZcDJEw2PU65dR3D9qD2ZXv/Dfj
/c0qvhkfeZCQdBppM19KFnc+TuVTPE9sElJ+/H7No0vPi4l1oFOyZbL4hFnXUlqN
pgJIptvKyZ59WCXfUUFLVhYvlxfDZbMZJqdNC+0wh3grzXr7bQikg8g592TZLWdc
c/ej8bCyB3M7yg/8wpQbJYkKODp3KZRFQE1n1h2dFtKFDyHpX35OtR3BEo8Quqom
iOk8wSrHf8/dMaC1zBT3/Sa8lzo2OWM8Q+SH1a3FzQQvow3hHTbDLLPWNkSMWejE
+dPJ99NM0xF2WmxAvn3MTZj8VyxesRQpiSD54QmIiyUhkQd+KPuNP8VHNsnAGYHP
9+qQsbgIDhhGBsHPHYslAz7bL/Ms/JZ2t9GIzrok1IRieugTcTAsj+4Yilt6VGqw
CTvJ0h69Ro1+KDz4VClNcWvlZroVjX6TqpsQa1MxeplVtXZq4XIVMp/+q4Q7X+Lc
Zpxxf+dlsStw0/lOSRQtdBWHhMPVmaXkM7o8mUiFQ81mrzjRldmhDr3/icZEnm7J
KmAl7KF5ZhF3lRxe7xu6W80zfslEFFveDGsY4Xu7N9JlfCzlmhfouSJIJMwCIbDb
N2NREs4S6wGdNpDXwA4xgjaU/+HUkwbWVDzlpX3IJWZhQOvDRLLEGLyWns+6TdE6
3RYX6NovbUMSUwSQp047Tdpel54w/MPWs9pp/uwlbl77b1k8Wn1MRAqLbtXQ46GV
4TvsCjDRIgCEHupcKHWZxkK8EK/sb69GvCN0clzIJqQc7crClFoXWpGj43ZGMF0r
9zdKZkb/Gfo5Dz4IfP6A+nzgpC6VNZLnLfFx9heHBxPY28CNkyGEWT5bGbSanfzs
06RakRwEnYmK/B4BzReKROeyHcQ3mUT/SadHNEkc8BKHBwo93iwL+LspMLRr5/Fd
knmGSbSi3cCUC+eoABNwNW2LnlVT31KA8aVF127wHdTKgVIPCWOplaMHFWVKTFzl
+/syrPj3YOjCMkzlKfYbeFfMIeTBiB/hJ7x7zrYWqJD6PzrFOZuW4pHZWfiJS0Wl
0ZIT4qskUhZ8bdtwvp16ym58VMgPVNiPGbOWMjBQ4dF40ZtXHDhtxLtrc9udg7+p
oxdQEyfCeXZBdrehBw8/32jumsRjHg2zJ3IYAFLnFP5QJjzqa49G8o6EOu+VTGUk
3GiUL1wGoXaEp6e+pPUMsgQMO4kVin0dNSsMQpytvk42aiec/cFRAQhttv7+Qj4v
OZV1mYBsMukwH0l7xSPHxvdtILWiMHq/npb0jl6ZMIFgQY0dTDwP8KxoohzaEK77
RXipckrKBr/jvwkLBWqTf40sEt79B3nYLL0YYkKwlb+LMiBc3JUyFMrAArgLKlsM
EV0DRNMinLVLjiaEG+jlgQGfyoenoY4YV8d3O/273jgt+hhquclmUF+7BI4rNbYj
bfLtWrMv7vIZHUgUk+rb6fQFdjDwt6wD1BuNwV+UDEapj/PO845/c2xKCMM0+4jS
SSbH2sK+ltjeHzu62tB6G2JQ7NHeiVR1r8tdCU/oShGOwacgBLAfvTGmWSNwhL/h
9tHBSTYLxG5H1lEI0fEMgmBdQ/1LHX/qOAhU0sOzrQGfxfcMxpacNpN/frBBINjT
41u4QaYRjwPTxWINbAWMJfclrc24YhpSAWFz1ErRToARoPK7JPqKjGsICp2YvcGe
FXgWIIKQmIhNT3uxtuldbfzzVpy6RmYU17SR+8KehfHgVhflB82oNgIumk4GkiqF
F4Bcx3Lo2AF+t5eoYTLuOfntLSuSiCLjAR7NsLAtt3d7YdZAHwfRKlevZP3YqsuS
DM12Mw8O2fLmiLkAmfEJvq+rYgSbn8feRvAreNTEYgfUlB275JNriqV/OqPCjluA
QnJwtr/2CPn0X5Ng5I2p9kta1vNQ6yeaLCDHX5cET/7wrZF9yVD3ww/K1qBq0VNw
neYs8pzwPHpankU4L2KySVUIHRi0mEtK/LUD85K4nlKnHRUyp+FJGvdk1q49Hw0m
oXR5wbFj1ElVIrlKrTvlxmjmcK1zn0UZHbCS/dUrT2Xbd0hoC/6jS74Re+Y6K/FF
B76UMkXVeGrlC2menhMkfCZeWL+NhB3VotgEEtLDDRpaVsTWPKr0yDsvf9CzE9KQ
A83XhlciClizg+uJUQd0WDVA1xYWMxfn14PRyxIGw9v6OrLRZOmdulChGsyVehYR
b8g8Cb89Z8WWrJBeKDKH3GHAwgK+JBnJgR0/GDUyqq7wsLmzan5t+3HgKVCxN4GB
Nr/bi9lPhMP33NIdMaPL+uC/0OKo3XkTdleUuyzh3Yw1lL2SxJWdhe9ezovFoqGr
VCp6BfM/U/vICZQU+NbqhdL7hh7UH7xh6RDSrg7xOH2NvlXGq5eLFrPKzUbjOapf
jjUhepKCQZnDjMKD1sX6MSAsJWzwP8D/tnuzr9t8WKZpOMVMDB1SomIR36KTF4Sq
7elbwjXSJSY3z8hrJZhKpru7TkER8Am7L4ut76TXsCAiQLOCifyATpE983ZqrXxj
RqMTPxsmc0OrezFv8GMDg9i1Tf59OHIFWyr4wc9Pned+S7qA445L9HLAStxQ+wGf
gFSuu53EbzXLu+TybuYzICMFwx+zoAcI/87V8dQ2uIFqxoYkx40HiqBGcTpggg7p
OWfUM7cD6iujJX/uFD9VQljNpf2cUi/lh1N7SsgEqf3wOLNxQYDKmFA2LgBDcm5u
2rRUREl++Z7Tp4C6b5IoGPOEDVVszBZxNjGiRwXCE/gdA04vqQ7AD2G28W5eQlNx
ztfjwf4l1LwCvHXPTC6Syfij6/t4NhocexwhiXCKo/iYFCwLjClALHkAxkELvUpQ
2sLwksI5VimhcPopp66xxHIw1b6df1ZAtt2opvEt7HwvPbcY5gP7MS6hkGFbdEGf
jwbYab26lztgluKOQShzWjbzL34KTuj0DImmZQI+pJfbIRFHvvrT0FZyyTuCXZlC
Tqk/WnC6ykSl3oQfKanyOvGfqjguuLGtP0T/ebJC4D+opTezYx2j9/l7DYv5rQpD
A9J2IXLX4rd+WDITINgOD2icu+HhbnDcO9dRUXkbq4yMEHncSEpSKAKJe9xKS7F4
wLHjmGrdTkH/VM/4koblFSt9G48DwThYWMZhvcy1OtV9n7eBpqwCGNFN3Tz/8+ir
e3seAGQ609tGX4Cg4yYKVYEx1JSJT1QuqpEMVahgTpL8BtwERM3OZGiy63zmWA/7
SnYgDaZmLITCUyk4DluM1ySvKLQaAgvt/PLfiljMnoaDdxX+pop1vgMV4ytOZ3hi
FpLDihNBWZadbs1cRPbm18sK9GjavHfgio+YapK8+uNfPNM3WyvltA4K8Qf/y4io
zy/ucTrgLLfsp+pSSIurxlOYLLUtwRYz1sxLb1fJUsiGS9BilmvoB+n3+MxWLfNN
ImaaB/FFUV2KCYApPQwdWxnepgu+c/obOAtuLJKjyPh4EtaTxnO0w0xSHaI6C71J
uXbzyMbZJOdTLxJYa4udTx/M2bOB5/gSV+V9JPL90PEKZIgcfIPMz5pdd/COsbWT
0wTrdensKrkwhWw6MNRX3Z+zRSy7wZFq8XdpZ0JThI330aF1o6v+Zs86M4lKb+94
UlUTCyi53dKEdUwPAnSpGhtYfBtEEi7DRXKjRSwAbDJOGcGUHniN50MMUQyVm0/j
QxX0Wv/dBmNEKl19lBhliB6OvX7bVqlAoSaXhGttRKqri4VbJRpjRZNB15rxz+xb
wSC6DLEOA1R8UEn8CbuyF6C8wd03lgGRI6RvqieJoBAYWEDGouy6duS9KNZokvVU
tdeq1Ory6lxQi7aFGjCEgdYhZOx68ju8UdCDgOg5ly2a6NKW4EZhdPmG6nu/IMvH
YDOSwHU3EEaaylEg/MHD9yqK44IkBv5Mhd107RGqAE12MP5j3kEyExEP+ZqP/Bzl
NI96LLU3lN0cKND6lWEeJmphVHDbOBPEeGBvBXr9iq/tQlz0kjDtdjOfCMHUnUHO
kVduc6VIlRQb0xhv64QKfbc12UDwB9ibV7Ttl5UFa2XbTmYItRa63DLw/cHaYFcH
FA55G3dapkZr9rLNW3uvMufeza7GyVYOvcwxbAKSrcKV1slQe5/riUToho/LBUnE
7saskZc3rZfH+wANiFAsPZF+hFU/oQpzIrxHBYT6AFlJw52NSih1sxkQK5GUbshn
3X2rqIPoG6c+eRQAlV8X39zOPPG0EnsAwla2qBQKGj98pEvPY1KnkJ3Gs+96QgKk
Ye7Ktrx/lCEOstqJcZ+vqCip0tjGSjs9c1NA+fJjZ10BMXfz9szjwgYiagflSWkf
F2bv65Nn/SYfFZTYDKO0esdC9KqZ99mllY0ROmM0Es7dukNFJSW1ejHUf49x1fK3
DEVboRnKF8FsGpgmruzMI4owIq3IYcblS8qSvm+NNKBdogwMZA02QRLU/O4++5TN
ql/G1v8PA9K2OFuV+dcaQKapulYMQp4ayk/N+ii/GttQx7ONHqUCPmhSMLJlZr2p
Fxfr6XkPkSwlZ6PjiYN00GVhK1OFRKo6HQucecwByFjJ1emL7Zc/JB1Vz7B7Qmjp
7FUuJZBOGZOUFXOh35yA/ZSq5gKjZlKEBBOLSUIWhHEbbG9TIvclh31S78AZwi3e
0NM2KjUcg7niDlVpdRTI0mXD2hNGimJHaB7EBGjVd1/kSuNiL0zUVv41DnkuHkYR
JAdUvjyHTkjVYz5svi85E/lQq52hZJHZrw1F8JTrp5RSlO9zMqUoMkSrglSTHly1
2AYTjtv4rQktomq9fQGOafZ4IzdGSQGFKZNc/OjHy4T+XLzBj1+soNlnAjpUy9E0
fVLpXGWveCuTnf+oH2rRFnVrLe0lvJL3HFxMXMieNN60P8ofK24F5W97E9lJ7OPP
H0gdvQt09EJ7+rQGpLUbAHsXhxS+Vb3yKw1Oz+LTDa+T1J+dWTcMXELdYSkDza1a
VFH5fJT5wdE/5NLCOSt7Raz/55AFYE5Fl+2GbHVo8dbRoe3u7hy+rs7eOatyVr/g
QOieLo18BarfgmZBVIFTXD4iE9/wMwvFJgALTXPaBHwtl2WgVzGKu0m1XqPCCWxn
jpB6/xBHySKlBt/Kvfx3CT8hQiHXJZVQBqR1+fuuEQnHxpo43rS1G4dzbdd+8brT
8LvDare36fpDnUoWALh5RT52KA/DtxJfGGhzKN4qLg2eyNhFVumOboQQKMaoudDA
MNCiwnF/e/8b9aAsRoWDzS3OrPCdFtOPHDo5SR3lEQaBtywgeoAKkN8JDG4gf+uW
7oTdYJXM92UPPknhIdAHu66OUN1kyNHpQm2OmR3t0vTVgpJXMTrVG2IVQgc4LaLc
xqtd7RBvERBpVsD5HBebUQBUK6uWHhZ9GQqJHF4oDZXdTXLl92Yu3pcrpyoowfDt
7I978Q9uQoFstypb6tIUVYdSzaZWKjQt1FYNTado36g6RnGi3NT1/x/Bratbnwzl
pEmc6IoMTSIs2OX6oods1W+RdmjC9iMTqFS2xTJVSTtoEpmVxADacdpNoz/qnOhe
FXxVUOJaYFIKcFN2WjqQZbQmBD/ks3EMaSifWAnIbtAhdT4puiCc1mdCqXvq1830
GgwV+l7o8hZKC9TYgNcgjU5WF7wXQ93EhpI4tzapgOnJUE6yXCLGNBRDG1R/PhMI
YK8xtx+iHXAOJunbbwKKGCe/F9LqU2NZXOElmmIKNKAPh97oXdxXeEeJZ9Oa+EUR
BeP7vR1jcY4Qu6yCw8hTYB+I+Hq9p6hnbk+sN9UdS4yGEm60IoMRouHK8rfh1sJW
Zg0winJYtzvUApwcUJr05G2nwbmS7uJ7svbFElst+e2ajFdGVtCeGA71bT1xcNN+
jK/DZGaMfiq5PxsW5vfMz8JjoGm5ALPXRnXTeBmS4VF6s6l7CyuEvku2vqzT6Ryo
KHfvV5zKzX3VdbYvsMNr+K8CBJp6bh2hvLdTm/JA4Yt6Vh3ndgwu3kG73C/EH3V1
mED9vEgKy89AAMKJOG9t7ccTAaBhoy1v772BsFng2quVo3RTFhphXOMuXHZ5P72x
c6lcCd6HEDoM2I4ablcLyYkeZ5NjYpgsk3VcM1hAQegfvetZnqx3NAvdsjkfryLO
AjY6LR6yYTAAUIqUirC0QXNq793oFnDMGku2Vv+tSC2Ng9YM//pQFLO3VI3JST1n
adZvSRyhbK3U5ts8MJ9zCbtZTQ2Nn3zJ0gCG5DZgt3xLZdvDDXIoiHuBOBcxe8qD
z+ISEyn4NHH1oauNxl0GB3C0oIMuGpadmKYm1I5cj4TAH5RKhxJeVVLdlgfvdxdl
cUXk9rN03KrNXB27B9fbeS13UoDRPbl81E+xorKoTb9Oo2yZ5DyPt/5onvKKeab0
86TaBoG3bhlCdJnJ9YQmhHHXxt+Lam/Dlm7Pin3WDCsnqj7kEzEIiLOIhqYhrhPv
8ixRG8n7eKgYjKH7x1DOvJiLHV8AhSxdn8ngM0oyHUaCBTVQBtrfjgEu8FSbj+RX
/JmDh5eqGhvmYotNh0x1av95Id7ztefRkrdUL0JJKhjFRUBeoAYVnxyX1i1ULEGg
0ZmcMdeSIUeuIo8iT35TzDu5zVfCnxymA9nCD3SKlN22PjMUV7nK3dpNo1/rrgxo
yNF1aZowB2JGMfgbtfoCb2KwzJ9fRkZsIMJxTMrpoYms0ZlEeeLkKjNuT1ACQ9yi
ENCvmuNxH7jaZQH2qmcf4qHfKMLdYq6JQ++8qioafSwiMQVLIHsndEN0+YkAfcVG
COYnDBEdzD1SBVN6KQBnO3jnXpU/HOi2CqE17Jdi4xy+HIteToJwq46ScaMyZ8KS
syEwku/DFHb8Ti0JurjZkpiyQtUGed8gYXralgSajIUwt16d31ltfkvWBZ5dzi7h
i+6/I774L4Iu5izKujxTPQP5rZC4KeHGUvxdIT3vh+MZq+D5qMjUenDZ+q4NvEnS
hyQz7I1oWsozq/aHFIa5FxtQqkW5pA3aKeU5r1GSrEXTmYJDbzu3C1rlE8HmHNcO
H8jCUFKsYFoUnFfyAzHC3pUnDsahs8kQPLIBwm3RIVI0Cs4q5s65zq6vRuJvrxnG
OlA/nqt5IxgPm09XF2+4zkgqj9aNtcTOLdsiRAWi5LA8HD18KD9nvd8/WunhHvar
Y9IIMVC4hhmWzQiv0bqopKRLnG+1uuvpZ49/T3oauTSjWzLW+LD5/wNARPPU0QaR
cg049MAZTliGFGKwzwOhYcMK42LRvL+Ih6L5WguUXQwdfPUOsK79OD1/XAePep81
b9rnkUF6EOqkA7V2Z++BEXH4C2M0qqPAmm8L82g+0oXQyrPlBInx5Sn59Kunsd+p
cFM4aaFGc5KEaOZn3nblmkLHr3/498XNJKEi1RSVMebxG8ZZWsGQy7FioVuPowNS
PglWpw8V0zszvLJf87UWrPVU0QZsrEIgaP84RNCM5u/TBunp+DdsEmBWuw2AjaYu
K1qwZmMY6kMK62kx7b7mHmCvBhuni62ieSSUS19fhg+b4HUeHlONBnenK99/KWdS
8oPBiw8oEKPsDzUGMRoSUm+XZEQk4+4aM3aCmz5y6tYG8MaDzf9u/APh00XyU8tn
yyp8Np6HsPbvPYhdsRFgRUIwqdIGqsP8zIYTEhvD1JwO59adQ2/dtetnjPZdmZPa
JHdBG0pacjD9GYjPLxn5MN+/CfMhXTT1fJrwwAu7QitN84HlxiGrIxJxH3enDJA3
VBXBv/c7Ogh6+nsxRss6MOAbDsmUruMznkmmYzhPQ5HKMb+wJB6YQ45Bovi6ou4I
3kBSf2es7z3drk46FwoglrRwkLYEwr+AIlzmDOv2A8TrIQd2bR8BvR4cZabNoo5v
eOb0eCkAov3hDcHoFt1kNDFalGvO72Z/NP+w+3EkkOaX/7eDnNLqgBNe5nFVPDf6
bLCQB6ICuYVkiUaVeU2wmuXJgwlQXrP7jDLm4zLXlflT2+x7BCLe+gFTkiuRapFO
B7Q1SUqP6tDSZGJcV+mHdoTWsSENE+SSUfmU5FfM8a9/Sgt2bHVudScl6eAnzC9f
QB2+bvppmgQjPR/CemulXNEXZr0hKDLbcV7iWdHJeDxitq7QyQclSvFplxMR1AJ/
4BGx59SEDDtNSx+hnS4ecfXNqa994LCS0sNJVLzNvxD/IjY94XKl6/oCo6r3l4A9
/kXLbWHLBx8GRMA3OpOxIe9drBNIMgcKZF7A7yUAbDNaB/0u+ChSJVjQSgS2FHj/
XG8PyRqz5QgBRQWVKChjMODSyeCmeENOnugtXFd5AnQG4hjwUYYHsAu2KwNawIUU
6LCrjvyTqvV2bp94Ww6dclIYNWzD4m2MAs7n07OymYeaX+YqSl0nq4VIxBy87YTp
IVbpdBW4rf8BlzeQXXY0zOvdjHyssEsPj5u69V9wKEbAwcvsYpkBYwOEOj8Nas5k
1nWK9te/zPv1BW55f7fChybeYnkvcK8lJbzmTNO8k9bHeVKRE+TJfHujLDuzKCHy
30Cb0UZDM5/hTWX4ehiNSez7nihjUdTsBEIxJnAombqK0RufhV9qaTU0+F3J2S7y
+JSzwYo3myrhrXb7o2r2T6fQgGn6j4HBLEE+I/Afi1BJbbaHKI/8NBwtmbErKCQO
GgCILaJKqcukN3F7G9D0VMycojSRrQ+adZw04gGq9MvJwApjlxiTXTRwVXkYZlBQ
TbwZkU7dvnjlkOxEkmju60ASKdDh8woduyISNg1fExVz6nWb07NKvkQlrhXq2ijs
MA13BD4uCB7tdigL5jA+tksPf57ujvU2TjoW5pO+reuaQh9jY44cDKhIy/HOlLG/
+bqjjSKq05IQJfNJHGZCUnrsguv8VJHG2zmpxtgtwV/5IQvab9yyXpx1ltEFiUZ6
3OhuZDmD39HMQJ/LXcDL/EyQCnpQ6iIfEatw0mwb5PBYqj7HuGqMyU2H26AcPXdr
o3ZbCT6AZO37zM032aUdG2mDxvYF48/buxOWmqe0ZW20C2tFYhNZXI0trxGv++Ib
dCYW8K0DcBKm9IQdiMu3jIiJ7YwmEMzetnjV6gKBzIEdd+bRQzY2QVXKoY/ehkJk
nWR9fRo4PW5VqQTMCr/unr+612mYXo8vbtOgCKQzVJzkJCnlLzmpt+qmjtM4CMWs
mPsN4HiLWKWPK5wW7ifccFt2qZdDPIdJ2Wpk4NIY7Et1WWX4TH0T9Kd2Yu6zNYE/
DWdV2IXYn11Qaa0hAbJ6aW2fd43cIuyh6kxEplxSrzJDfW3cRdqcwPg1GMVKVHxL
NO7bTnMOFKQ7PWr4GBgoeGuCnTbS48J5EBJOE5STo64yLRBhZ75E+gApNBwMCZWo
ZGrB/hA+ZznVMhsG410Ebiuye2P+PWZsZFvrDQeq8M13RORyHyoXAIUumae+3frc
KtkaIrAguX1sVFFToBUM+FRggy0c1k5EK9OASF9zNYpn44UzlSeZ45giqF7b7Bkv
teEX3qEqJceZ4UClD7eFkEs5vqrjOHOyU93K5zegWR/Cy4xA2L9RjT+Co79DxdRJ
nMcstpbbuog6erC0/7rf8xpguukcghGS49q8PA0WibXCG6TjABDpojP7mhfdccwP
zZfN0g7O3RAnjg0Qp7M1M3WOjmLsOpN2KS3kNffX+l+mdbdhtv+HvFtSpBxcQKYF
eAGFk6ughMAm6ERX15Eyb8cYkAjdlEgYsksrf0LgiJe8CW72cT0zvGI7xFVXZxAr
hnNrrOinmtKRX4Hv4uIwZenFanUl9EnT/XDLfvNc5y8GDov6mlbhtb7+ft73lzwW
ZO8/GP8YCZ22kkOCDWmn/TR3TUh26GIVykZwBBm7yra10/fK3yfqOfUTfs7QmTv6
K0dNl0UzT0f4TU2gOvbRHcePscyDHs0Td9VIRbYLGM3Gv+wegXDhDrTbeBgEtySe
G2AeWlPnbDyhgRSKyonFKhpFPTXuKV4v9+SElDogzqw5zWx5tB6kFoNG1VeGUk90
acenXwqLXNbUN72IW+2D3uADpxMSYTqmNDQWxXMzfZJbkY/fWq2ls7fLUSdHKsW3
/JEw1KcKEaDb5crszftVrpE+xE3t5PFS4ZKBJ/uHsocAvWTcewKGa6FR/LleeXoC
V7KR1X1CtkHt63CD/f1J7gA4mrjE5T2KqIgvOgcmtatod32fPIpzEk+1sCZGNRZJ
hw5V7d0Q7m996w4Si+IMU1Zs/o9W/CNh2bDjYwiPTNnFrjwHvup8wUvGQHjRpo+k
79cR2cpWaqO/H8+aCFsiMhCYrUfKhD/w3jGMHX1YQRavENWd6RQwddPyDxugV9qq
gFKlnCfEQwF+i8ZctfEPtqG1ZIbyzk4uRElmFsqwb49zk0H5KwLWPWnoH/7t2JjM
iGPiqGaPmOphfMB8PPfHXBY7CnAO6Lxl/LUGF9ig0Zb1jYIDuZg7S5s507qQKhTb
G1XrZgFHLPM7j9+c66znG3k9uC63y6/oG8GXolMiSR/1CYZgjsseUqmqHqzfXxH9
JyjqZ+o2Up4NEFDxEaCEjH3UmuordFwL6xNpYkz4SHmSh4bZwG1Tr/OFM5v7LAiO
CK+XiKPf2CWBQNm3xZ7xOB0Q286vuP767r84wuyeNJxvofy/U3M/oIqUesdNBnOy
JBXe+uTsoFdUqAgVW2mcHdhfokW9RIcKzX2YxjvzPZbU7GvRmbVyYA63B7XCU+q1
0jTYwXtX2fDJnMS185Dgi7VuZNItVNZSx+Xm6GrshcvZbRpBAEBHLUX4+iGBWab8
Y8r7Z+byq8zehsmUpUSB0q0pjspzWCZaEQ7oEy2idI6juVHL49McBH6XWNiYUn1q
k9SK5JKV9V7iI2Vd+20AMe0WyrBR73Lw+hKHoY0S3BT6leFr7DxzhQcXT8jIeEr/
ZNfiPWz6R26Xic62ko0Oy0yKvc51EgXEZvsY7H80LFnSM/ohgZvEvnl8HgCgV2KS
wyjjm7+mA7X6NYduGHwz0RyMhLwP7PJE88o4eHADDbBAhzI1znEROASl59tZ3Hwe
Yx/C2TpXtVUPOV+YEfX4Y7b1Froqv+YjJRBra1iIGhmlP2TswGsmJxT8Nr1qXefM
IqLpugpaRY3QgLljYmV4E/SfImeYTqQuIt/24hOWHzoMRsAf7wfNdm4N2d2jt0NF
x6IO14PxqbV0IeQnl/idjmiJkvat5bP99iCJ3naoF7SdqN/ndf6rG3vOGzzzawuE
NmK8h6Iaj+CQCfX96QpkFPwF/dIArlcGXXP+0JekLsoVR93aoio443xMAXww5nYJ
Q+EaAfqHo03TR6XRunDtDV938Aqro91n3w5bkPRMXOpNgwzUgl1YikBZvVW4n3eg
kbp6yzuI2GJpI26FTlhAq2jx/91USsmDGSaoauFl15I6gHQkVnEgwHX3X9CZqWf0
Gcbl6fnzUcWFMQ8UcaJVuUXRQaaFmLkOaLro1+q52pVboWtayVuiZDFlqNdNR3Ds
vQQP3IGPU8ePDYgD3l2Dsb8aWyCVf+ImY+Nh9Ck6D65ZbSlAJFbmmM7clyoLRf9e
VUUPLUEhY2C5wOzpFpFn10vnvtAO/Np4+2ZQptElLGRZfLyr+CVv+EJI99T09b4L
tMY7dXGfJ2AGaqHgjjl3d9IeCmqArFgz8qW3efUeQIanw/Vm+T5hRnlIVMa0ORwn
GU9F9lQ96j3G7BzmLngK34m8ZDdAHJi/Zxr1iAkxl0QC6nzpxMiF2O2eIockeYTL
BoqYzF4DdZWWVaww3W4yCM8PhqpctGbz0K/muYXVZVpuUWugpNhEIxGZk0epZoJL
/cxVlE5yFxM/GbBjBaAIfayS3F2KgpVmsP+m5v6/6GHb7XFLUjUDXg+ZSrMMhW3k
uCHkrzOT7uvEd+N4naAhtTMFS3HPuuR5z8aVlmJIXqwh4T1K0wYWXwqzaaDEXcpA
JSJgHsqwPw9S2QYxHVHBF3RiHdmKlSa/qcOj5WrXD99SdQgRZR/zYcbOIgqTkU+j
zsiTRs5FSl4KtQ2i2FDxv/ASO+C3hr23daU7ZK+463yJ2WWLrCw9UBuG9Uv53vJM
mROU4tIOPdZ0cDSR5fq9vpbipWxETKNdQcoFdXW3I/04dvDxavuuv7ts4Ovtofja
mluCSrZa6ZIqkh4PqeTO/Me1wSZNN0/2ZSXfA40RMnbr0HTJwuSERCCBHHC8XWWf
qsWOuBIlGwBlS17vIVL3/PE629zZwP1oaBAOBhSFvWhYo/gHdJGSAHZpfnvTRJ5a
fwc3IO53BwBP0mlj6jrBfRvNYvyUCh4jaOLikqHmyhDl7rj+DKff34oxn0di2Su2
UBPC+HUzCMX5taGs2jJE4TglZWcdHNOHs6dO25KsA1Wj32FU2tGatADRp98Oc6OY
yR+f4aHYLf0MAwE2tZhaMMsWqoSvW/B76PsKrs61cGDskvY+V8nWDoaiH7ixYpWI
M0lOuy6DfHMTESV6GwQ2ef5yPAyfY/TyNk9BNO7ggjsRVhXcIR5YHRymzyqqzn9n
ZNZ3bcbI5ZbSuhdZmLeeRKaxVoGCVF4Rxg/I2eMyQv1uZTIuRh9QKPfjJ5R2RCeF
CPpsidwv7L/+uWZLKM+Wa2v1DTPURbgjgS5m1lLQep1Lh8tx/AcE4qh1xQDXG+PN
4NEdVBh3O+OfaB5nYOntQU6jzzhUUt/FfrLbL2jhT168YLCNFIcD2pkiKy0gsc/L
n+3+idWQklDjx5d2OZlvPsX9EySyKoC3me3W1v7Cww83P02I7DGda9VBfXuYEEbj
uMkosrXwnJSpE4kXbnvzOgu0kZ9kc6cu2lkM+41/U4F5NfSWXDTXf/sFSvoExSNk
JBfaUHGNbhuK7cOvT35RShwWjFq+WEmAviDqP3mNjzLkqClX1fWXOvRJhn10FEuX
M4oOyMXMthFuUer90EPNSPDzB2PPWp9i8y0Ce7zhDFh7xwKjsmS6GoxVFZUO5F0m
qEc0DU5hiB//S0CeZ1TWFxep0ijskgkYGsQcMwpEuonik4gqqLj/4v0B/8yOKL6O
IjbTYS16I3PxRMpjA1MwlZdRTkDu1U1UtKW2upa94959SP3JF9qYgq3IlorHzA+Z
8ncgEAjI5rvsDnrxZvkZgNVKEJjDyEervLDdbcTPOMw2/U28nBsZZoKX1d4afURP
F47sMYnIHW1VQjwbtK9TDNfwphx7UzA8Ecpsz2ASjPs6coUQ7Qs5055HbQzvYrYi
XPP4OxOnpGuTBfKDoSMvY/GV8LqmA6bTnaYrbQuhD6CY0ZHR7/OkzSteX9tcJSmO
t8MyFPUEmjLdBexAU0FhLJxMly/ly5WyXQZFB92yBlpvIe+q2YAbCx4GTtaJAnSc
WPZLEgsAwfqhqiAQ6YzOfowpqMchPkcTEthFt9b+rKRvv8NrsIQOQog0r8GdK5xq
mZ0jChJPt2//MNIstm/ZzCBF1g0WFkQTqtr+MFQIXiZT5KsuDux7L3Dn0GUPpbS0
J42UWHwLovUgD02FixJIlow3VcF1AU+BQWelZxUQ+p7sYhfCHJ6SrvhvWt4DMwdS
9vgDxj9/ZaJpVU5Hvqg5SXLm8HhnjXvc7/k0D3Va8qgAphiaPDluW+PmTv6Areei
o23exSAFptu0r7K2dWe43r9ttq6s0fH5zmys/b9v8rggCZZkX9wwyDBPMEpS83mG
QHv1dN4KN7u+dV4y7MeBoBC6gHJOQV5TmmVGrjz+x6GGKy5vGPrA6P1OvpRXlSW3
grMKwCUxug+CFbBIIKk8K6LY6LIxnhYGHrOxdfFRDTMbgTXo+U99fPIrqN43GuHN
buPYDqoXsW+ALP0azIWoqsu81mN4HeSzpH80Ju9qEaNlgWXbwL0HDHsNxTgx28EI
ztVwR+qFQUklxs/k9V3wWBgBAQeus6LK65Cha9fWoaQTInw9YWve0ujC7Nknrv40
Yb+4yzje+w6SpI0BApkhTrXWkzKH/3sZoqggHAj6Ob5NYyYP+DC+EJruvOywESuP
Hg4Pb7o682yQx7MzKNPal6JmnTVJxqEfDL6TCxlVXjp9efs4sjcuO+EuFL7G6/9u
4M/J9RbwG9+GWtche211H3na74lBBZncdiZb6d07UhQms4LuW/HzOa32yRb34WNW
b4achShb1RGVsvnE9MrheHjduwH1GOlhLoNESVZsZmal/cxBIkaHxnD+Tg5qnSMh
UONXfqXuz+17sXr/GRJ9wa7Xb3LkJrfaq1V2CK95EBz1+Od+LKfjI71hRJ1faJr3
tqY7kqAtlCzdDA2BxXZ3G8KACAk11l4+EcTsXktV+PzncESFTm6ruwJ3P2KNG1yI
udULUXBF0Q68aCJ/eELqoUfGy/G6mrk2bkaf1q8jWnC/KValH/DtpPMxBS3MLINB
wo+IXxr+5/4z044DCcVfp8OLll4xLSbHaYSXPHfaZeTsmOC5SvPxbN96hWNY7hq+
a5LneM83ewhF/PApwxGqJRwaX7RR3LUok5opfPb89x8J6S6fFdKHNj6WLjSyzZYE
39LonxA14SFXDdfMd3PzOL5qctGPpHA3QjBwWUySBItmad+r7ZsddAkiH2Ngjqo6
h8BuSqEFZCyf+jbRtwKAVM9BNfKHfXuTa2EV7jW2DkP7gdnAvQTthmYZv7KRl5YX
JMkSh5JVEFztsyfz3bmrJj47oEj5t9DMnpRsPS7mW1XTYmzfWbbcammuRcTea9S1
sMUtH676UdAkHVr/Ymi46LYsNE9EKhDpELnv+sMddXoEdMZzWA2AfTyEm4n4YHW6
W1bEZf2yH2rmB2pL3bXWcQtEmfzDqhbZhmvfBzHEzxlyA5sSli8qdw4KPkIU7igG
/udeh+mbSLYjYf2KJLu4SF5Z+oxvJBeojenGSaS2LQKqRarBBXuBHN4HaSWUltAc
O7LTOMESWGr5M9HkX/tMjIAj85LOAQLacEk5f7spsVPoUydK78YbQNE7lN6rVl6J
Of1bD76Y5uONT24zFLtxmJrHuQttsm1MniWw1jXnL/zKQEPvyL3vcLUNBUrnQfEu
epHCBKV/slr9ydhLNN+dXRS9uyykIm+WodjI5ZmnNXm2+fYKMWkWr1M6yMlxRNUy
Q4TT1jdVuKLUDYWkE1lU4YlRlr9NkyCNyrdpkUku0fBUObYMbKs3AR9tJcyGbaCh
c3MOcyqKFPhPOouwvUMHZz7KcYixTFxpysnRFY9DonrE723OT52klr6txxVCRG0f
3aRdcPdd7gb8XB3wi/DdJzZT40qT9O0m3vSTad3nUlwj+XItjZp8pFYs4D/ArxMX
7SGQpntfMsuZ714bI2MbTPEekRTDgMoEoQdDvHNktIJ8lAo6MBdrvn6R2+comFHR
3+fBtNoNT5VFQqFS0eDfQTpa6/p/wHbihIIgMAWfUn3z89IDYjxi8ncZAaO0bRYS
KEIkNlP27HkQZFKWZL1ruTkpbsc7fkew80AIWB8X57GsnqLrl7dMxKGuJ/XHq1ZS
NZi9ga+i2pu2v1zd09Z3Ouwme5Cw9NP8P3ED2hJ7U+PkE/qJMxTlV3DRaKcla+y+
FGZ3hZHVof5y5Ii+PIHJtWRNhk9YIhttovvXbBWboGWOlSBKA+uYHpTFluih7eF0
YkZpi6AlnLvLDnqbDVXpGMnE29sk5PzfyKjXh1rIQtn1+b3/lf2aSuYcG2M/bAcf
/PhSb2anYnxUNo3c34imIFWR2FudBPNsAwyQ/y82ubsl3ixYNZKkgF1Gl1+WtmFl
rxMGs6bB4n6gnbvv7oyJfcPdh2Xm+S2+dDDXUndpTlN/07Rq1CL3kH2eHKep9n6l
QTY4GdccdHoloWeSqwJnmMDmmN2a28wXrInBBY9+spQzntNzYkkQpa53E56y2lLD
klg3tGvXzdeHC0kjDU9anHSuo1Aet/P655asYlOfadaicM1+h2y9o03VD0+1d1B/
oq79Vzro65nP3lFvQr2BNHNTBUYIQPdY7bRSnV4XJML63ba7TF/Z6p9J2HG2aDJU
NQiQcuGXtXipR1vW++pnmBQypcjinKbu/GA/GctQ26iXR+P5Mb5r1Qr810kODefa
OmgdZCmCkplxI6oGdbmzKwWlr9DiXPKTTI+S1Q2DJyBWn3vh9OoUKVsD8Hu8vxXA
I5wqpTHQwQXPagiXvf/FizzQhI0KAE4nGhb3ZmE/m2vxLHFWeugkCiMbylwHkHJk
N+PWGN0yS+5lGdOZAD2lzGkfsU+crCnN8RfVcdckfBsjWq0/QUA07m5lIxCBOn6n
LaBzrhJb4vBBOpzseM64cNM+3b/Nw4nEBDE8USnOoJjpuj4YSixAuVtAALPenha1
Ili0DG037bfHALD8gVWiBAqh+HRAgJS7JSbElnYjmtguolqK5b5d83isNIHXIUgp
x4DzxPZjVmeZ2zDBJDXsc5NJoai6QZ9HE8Hd/0kqutrbJPACPaUi4TENcGlWk88q
tqyOGHs8BAskHiatQui+57cbknGb1U1JM+ZPb8LNegC8+0ACCaEQBmPuKy9DJH2v
Y83vKSkuld+fbRyWOcgbOdla29gcV3kGIXbyDXHFDfdmPE0+Zfm3QKgr/qyVmyC9
1lqV4RAXmJDnkAK0Pb/shcmSS0J3ZYOToyBRM/yme7ypIsHgl0b7TvMqQljZVa8W
CC4LHQLisEnGn7Dwedy8iKlbdq+nWHvU/nsFk0t1EYO7u2nqiZzgROPutBNSSBuv
DYw+Uvy9ppzDRyzTAJVO3sUj7IxlwoonrzD9qamf4B5XZACKsHx2i5JR3+AVgnG3
S+KTtRr9/92XXOkWiZCVJO46xSNBS2j8TR0cK+abljaHA/ZE/lpFMehOmR2lOnTr
WeHJFhx6awOsTzaiaBK0KkKlbj1u6FabcgK9wVDgDH5G/V7mZNPlr1xnqN1SyxlF
+LlEFZp4iaR8ZSWcKFJR/auES31ltFpl7yE3mLoO2QoZIGfT3Dvn9EgnCa5ZUrvU
9Waine6E/dK2wLwCAipUeSDtSXyarqaCWgtNTD6xq81M3uzYBKnG0c9UKsxi/DaX
aZkp3o0dUaE4qQUM9owyTKr+YdXV/XT5i3de47CczUEYEWBosl1vALFKOOXsjVyR
X0sAFAwQoHQZU20z6HgwJS2R5yUn+yibVd257Ivp9vkxbi2B3UyZeV+eMQrqEoU0
Ojl9thH88TikcDcayUhSOcZqwx08NOrsNJNYA3FBE7Q6kLuW5zmK3EDyO763YE9T
cBGCqidolXIOug9fpB8JsjbdcO7Y4FlasuqyjbDb9BvlR2AaIZf/QdtCLEKAlkHv
MsDX3OJTmgdDzXFAFu7kPLRT90IDRV0TbK1D6d+eh4zX+5K/GSsrKPSVIwQDK2rq
nYO8d02WkpGB92fImdRwaKL1kVo6y1xwM2DHBhocGYtbocU7E+eYamdHHulWae6o
ZebuG6fUCFGqPseNPAODaDMS9sqMS3BzZiH1R052rAWgzj2ms8dw9vCC2M+7Dv3e
u86rAqZJGXiKQqov5N6b7EdhhSgZuQicllu1tMqs0imEfJBizFeVaanJaibvqdJc
5TsilTaWi+QapevgGhKwVq2GXzzYZxQ1mXnH8pcXYTHmlvslTDEn/XZhOnBRxMJ6
kgBpS4ImERKHqzskZKv4peDvrfk9zukQbQFtDrQvTrsQ1X66OVPLRCSijrPKVd1W
OoOAanEKHx5DmmGDcJCoHzaEU3MnnyCSvKmYGU1WLHAEAxDKvV0G9Jbov6RnbyN0
J+qaC6bBMSxc4pr3N1zCZxF4lrHpawll7xTNWMsib7IgC8lry3kg3zuJWLjCn9Hl
SyUJ6Z03N6BsvqDz8uwJU0A/7VpVkUG+3n0MeS0URQ9ynGfqfrZzGauoVR8+3sN2
AyR8qCizQzIjC+tkKOiEti49Fc33RJZPK8X7eJ31rEzRYCUlunbMZ5prbqY28ua8
aPNTw0+rHwqyDdh20BJhHhxKv1V26w4S5ZDTPS3VxBhUUTAos8BV36uK6WHCpL2I
HQnwIXiqBaAPbigileoKQhe25WY8fAkvmXgh/YiSQtgMfmuF82h6VJFIP8nj1FcS
c+A87Ny51BXvSqAw3ZPmePPTgNYdmDYoYmYBWq3QnKg+CEzDjZPTtWxdwjm6DukX
8Q5YN6wasTYOlkqguGl70y2rRLKa3ME/npUbZWgWagUndcC9grLt8K/o1ux3sKHy
7NFHfIALG86HS8Ab3r1CEF4FZ3Ei2A9ZVT9xC5k2lIi80OCpv8DKa5O7JjpYHIcL
xqhuYauvdvlJCSdtGjqvdfhN7mm7zI1uWrmJ03/dhGobfM5EfzaRWkgonQdJZoka
T/EjJDv9uzL858gADm3lnQVj2rx4gMZNyC5FRW47bwSyGTL+p9WQ+ahpyltv35c1
dGfyOH8uvh/f7e9H/rfc0ZxpDox5PjLgiKxwyFw6oEXN9RcgUeqFXZ4IzZpHbRTJ
eUX/9rR14XT7CmebNcsmW3Jmbb7XsGhQyfuITsl3ZOheAShVTZXgYbUMvoWwJAMD
4wWAUQ2R3LFAkbQFueIDjKsS0qqKmh+Q2ohfByXt0s8lUTmvPvW31oUBd1cueR7o
BvlbXU/527aH0n33bW2n5xQY3ck/MjG2lEaYau9f+eniAHRyXp9yDPVlxZP6Kqyo
OLzX8tRZ3HKdT1HLFw94wPXcA5LCTcGwnrKeW4Cri1Jo7j+Ao8gUqxsZDT0lQksF
6iDJjUYH4gfoOkxGqhgnFv1FZQqdX6G2H0Czk+ThMgyeLoI1JiPSdnlzldAqBmp2
2NzoJBqTFjlJ2HshLnd7KPe3W7Na/EHHNwcYM0sp0uhVy01GkMWdxCOK3xH/Xlev
ZJUDN52yPq7eznOmqhA+uIyksf5N4na+4HR1slSigC55an4D4zDokPBfbi9jDOlB
XZpWyjv4BYzCUQZRxyHhaOy26SaF0W4As0QS7hZ4MYSvBUTG5PZ4R0zH4awYEq5/
bhxZJLs8+wwaX2thVZSm8gZzr4tvuiEgDXf0WOlNBDoyYJ56RTcH/SGPs4ym2aY9
kVvU8NImHpffbN1VZpN6xPavU/NS7iHu6f0z7mx64IK8W8PnbcFOPjHt+DKwv4kW
FqupAaEOlx+Q6KToIpby30BOTOYlu+rdcVAvLqRo7GD3pBMKUiQW6gKdOOrxqUwX
z9d9/5nyryyro9YLPWsqBUxjBMGAKTBm4NVjUktbEFrk9Vt3k0qTk8cj8WYBEVRq
7MWaQSn5M7CSGFqun1p7Wf+IXi5NpQZzm/0z+deLyBQGYdU02+ZJC854+x7yrZvb
An8ry/5bApW/Kk+KyeMgbSPF+OrdsZJm5CqDBkm63m9Jv/WZkbyBgYjFtRCoOriy
55NXGEVqtB1C6Jm340Y/B1mNwI3pV9Sq3eG7PNQoeOKRzB+3bWc4ZJ1WPti0sP0w
7Twt8/JY+7e8neyxMaPzVpZ6oH59GN7m+MIY5pjgyauKG5KUhCu/iPZOgwpd7WAd
SviAHdxEQa58KKye5Z9EbtURN17HMC2Ju2A7ttIe6YmMi2KTiRz0k1hhC+aBDDuR
NBoA/+M82X6P3lCk70fe4mfrcs+DUu6d+7Asbli9LkV6ttSn6E2+gy3ckk73dF74
d3KYuzXU+DguebGFAb3bFkiwjOPSXskWaBR1qRLE9NLe5FfoVYxFCx1vj2EKWI9P
LHQg7J2KvuerzntSLdLUEC1mG5VLRRu+/Mo6rA5+KRmTGVLMbQNHZ4Cj30UIqhNt
UQFa/SehEV8R5fFFMNjs7wGwbe1G0L4caVjsx77HrPd+glV6HOk8Ty8EW39wl7Xf
UOjYZSitosYkZRFdrreRj8Y6q16LM6ol8g5ywRdsxDz5ONGjcnBcWuhCGICt5F48
VpTQceuYTd5JqEYqPvzv+4pgNpz/yUucbAr782NgDpaVLScIVviSMaIfdaJjFddb
opMwsoqO3xvL6Tys6vEOhxer/0VK/b1waNTiVBMVMFUB40E7KrMNxkQfomFJK/Bg
1WRQpJEKqDyMCrQo4ld96GSp1ESInfZbjmj0zzrfRTfo2BD7K6/5HNbm4QXqnY+T
vBmQ/2y6Y+ql/AtXcXPtM4tCbV+HbsqexglsECQOcnrj+SLjDDT/MfO8Oymo+JIs
eXrYAcWbiLK5sQ4V2/1EHwFgP6dXHnoREA36y8e2BIYffLraS6ewPf9zU7frQiIj
pvI+6+qWdKbO9ryZIIwG1Od1gMYrmldayZBAknbsPe9hdorb2luMJO/bRadMSTEu
Rbe7yMJTbPymQ2Bl1AAy66ksKxapvUbDo/29MNAefEvTRpTKnpBI9ZhMNDQmUUtf
O7x5HyvRQyvvfuncc46KWkOfDrLOiCPCBG1QpAA2PFlWOma9ZD5audKba0zyo/DU
VIpv0XExZ85QEVjC7BRJb7cII1c4W2rEHz8GZOrDelV0Rbqdb1bSxZdu4VUoMC/o
DFNzbc8PqIw8xoD74X6yUvSji/eansP0feZlNuxbYU+WsfdF1y44KK8F/oY5A3Xt
RVc61H9+oTNqhZyf1/hSH0rHTs8Fu5rFn1KL10ClR5eWUK8lRdir53RXwJfH6Uwy
/CoqucV6F8kQytrHa2vy2Sqy4Dahival31slERKqOYBMVmQY3DdBvXnTUSZMYUr/
KpU8JjPFmjL69bm/UxV0sg53r2bEJNvUg2hwSFl2oS0TyODgFB1JPaMNHSpfuIUR
KRXYWNX4oyMFY57YX8Qqt0LCQfLJlwtcjMpDv4UwmXzlzOgVowpQCgq1jxX1qQY/
+qoTDs4g4iBTYIkDFZ/Hjl5d9iCGnsYdMbM3RgkufRxukQLS70CFpiiQ3FtxrZjs
2+FDTwA52Z2+qBeVvV/tiewVuwe+gA4xIVquLdRAr8/JdsRYuzVLhQla0rEArmY5
qfl6FnumY9N2NmwpQkcrInLGpO3Nrgn8K5xmUAGyIxAOtpQXlb87tbSw3O9AF1ZI
RNdzvfxOOZiyCPohFt/uyjXK41Nm0jgQFSqFHOZi/CbpBgmiHY1ybgcowwC4LH29
u6pJsglPdPU+Pl7UnaSv+bfv1cz25H/XCWXt1Yy2dtaQRFsfYFl2aENwV4mlXRme
7C2CqAT0XhxCfEgV+h802P6W5GotbnDNU4pJgaB7QXBIXvqOug9W3Pra8CewrHf2
ecrxxmfT/eep8Nw2hb08rtgcCkO/LUnhQ4DX5Q2FOWsFNseMH9z8OmEIahG/g2OF
X3xzwPn/bIFBxWY/FTb4ZwmdxCmDqhP86y8BIF/z8wNHE11/hx8ZsDsrnlHPEaI2
JpnQMw5NINvHKEBKVqcTbVPBfhiGWs6sOsbGsAH5L/BSFUvDWuSAPSIcBSbe4fRo
x+ZuiJmSWHrduGKLgi9V1YRuSLT144KeCxo7R7GDbfhkygo/klnWcLEb5MEg6RpE
IBjsrjwd+9a/pH+M/BsPQ1y6KlwYCEkNeJCu6U2EAlY1LlcWFWw1+X5a7kYA3bOe
nGgWA0lNRD7JstpWK3NVcM4XcllnrbTytNSJkNLX58OwnXhde/xZEF8p8XTjBPlM
Ot0UaX7CYk7XjxXvAeAHEIQeAvi706ENNk8/MzjGW8nH85IDGvo82xCtLq0TSXxU
S+u55MRUrVF8+QdNZJUqsR1pyde4wyfhSnK4OB6AKvSSKLF0D6ksym2x5gBuV0gn
7o2gmc0cAoxg9LB0fTOkU4TgtrRkzqr1XrYtin2jSX/tzOZZ2baR2uPDc+839+X3
1uf9PLWGT1cBuhBxZg4J+Fh8boK98yl/9GxfSFJYqrUJxXsxeM7hnKnRERVVzhZ4
AuSThfauipRGhoZNFuUECYDLIXjstbjcezxqjYePrsF1GsunTdaZHEQPwp+tPDVo
It7pufNDSSbSkxfQDlHvJImjwP5LMtOQZTllSDYGXRgCjB420G4BVIJKLNV2sXMh
Q0NgwZSqRPaQpngHPY3u9KXjN/3g49w2tmOkgTyAhVkrxJqI1xddbBcVSHhiZL/y
dx7BBhpbBFkcx2GbeeJ0OCBrLLxRjlqMkm4hQTMoeUpIws9Zg7yirE58iuUjRYP1
1pYdCtD2dkQulqeA4YBFnbQGb3/GEXOAdVl5I9y3JlgI7qb0lOAO8FmQZa9ZmaWs
+fxk8W/jqF2qHWv5tGskfcarm+N5KVVSv4QsmQaVn/hfM1kQSxfoDOSQUOPfUlJ7
JIMw3JS/OQZDSE0klIoONgZnz9HmmCuW5u6nAqxwA+yML08YxDG2PAC43J/Kt3uw
ayipco7FXAiUmazX9Mcm2uy1ph0zKaU9fgy27lfThL5cAgRN4+nbV+aCc+qYWS88
WMVG79gWu2QZUQrf6s7reTZKblPum2gSIa1ZP/09OJU6vUW6VIqBxOM7y67Pnc1l
oxOerRF2u0CLhEKTFk55ZzUKP/DrXZ4p5nZt1w5PUWt2dVKWk0Mm0Otx9VjoD8z0
w2eHvS6rETLHweKHvWHGBVwzfpVd2Npek/wVcRYzM5a9RkbTNW8cYF37B3Z9QcTH
3hsz23hwg5q+caYaIBDwuuz6Fg5bPIKtBPV5jzXGTt+gPGrnrc3ijHJNCn9u6Qc6
wdUvBPCZejtagO0261Fp1UBnDv0Nk9m7Kb9JrwDUk5/m2uadIKBBqGgdKxUoYG6Y
E55b23SG/K5sk7YpvQB67XKOfPs5UWJkRIrghaZEzgdzQ85OTNco7aoUvXUpWKB8
sz9KaqGn+OYc/d4k0f5cUoe/SK5Crv6tzhkfuTEhsVPC6pZCYfTAtNIS6jMYBQtC
ag/Rtiil05KLE3UE700oYAoPgP5RQhmh/he1mhFq0LLjh1UKwG+FMjEqQpUSNblM
SkD2FkBr5GYt96y1FMkz20PQA7i/vSZH37ndvDXOC2MbRbXRzSunQK9fRu0B9FXJ
DAciwBaPGhNzMLy+rfsbjvj4kYzBZ7YIFBkSo85NDNrQsgebwHLk6IjmkPwLfsyj
a2E0uef0tQCGrbc8fpHpWkYX7BwRJ6Fi996jaebb1ehf9OA7DzNXYgqD6fsW+nd/
nLKUU7DxTvm4LHu1wXJSmUFktvyLf4OfAgza/xE9RbFMA1JLtc5Y1fe+Frddhjmp
CwWSkkygKUlmrXbSXKSWrBK7/PW3/M+yUB6ZkH56GpG5nnEY6T6Tzw/k6wY0o3d2
5IM99EpEp6PcO41ry1hMDfUeBlmQQLfz0zBEimXnUOzU6wb2RQrUoirYQmwSssEt
bO7/5gbBFEG8CpagsG5BgG7aDIg12tSGJR8FnP9tvCqF4UThRl2XwlfL9dA5cwJ6
WaKwiBkG4NJtEvM1N5xA+eZYu8pREIgQ/CoPaflArvNtoF058/tesTYWT/3VMkUU
si+DMayoxG3wPKBeeNxyi8W4cQAFIFwDNfnspLJvTQpsBHLvdClJAarloMjLmVki
/z5OAoeiPUwqclzks4jjRhGp9n4pwxY3f+SV0HyeOybWCw9llr33wORDgO1tDCRc
2L50Ohab94rEGU1rZDStL94pAPxUBAmYqyp8hjYk10Bl6W2MwtQfq8CKcjZ5yq9Y
VpbUJklMgMVKL0xKlTYN984x5T4wcODwClPLArzQXGd6q2qzANxcovw1ktPOXq9F
TC1D9kishOXiGKu9U2PvmmBZ0k7Ihh0hpJ08bucSH36cFO660DGW+a91+FCPtChg
eRTLwyghBhFn6AxSYEnvRje4Vo4uCXoNcax7ornVhUstSF/sOHUh6v7RUvgyfq7l
AXJeKS3W8UXa4Sw3NOCEQTdzBLIvVxQGAFaes7OHfWc/XIkiFRfrBM7rs/o05OZR
1jUQe43rMToCyXFrKDkVX2Kt8PV2zs4xQPLrnumMJyord9UXgx3MeyKTRVxU1N68
knZkUAeplBy4JAldyTt4IMtYGIM8zfzYR+lhPqvUwN6IMdSHzhJp0QM46ej/16T6
sQ3VS5u9HNaedi5hbdEgHL4hk9tH7nSEXH0o25wdwbXiS1Yhop2V1d9n5FdrRRbz
/OQzRNUsu+wkH0oZnEG/gI+mNApeXaS+lpFvgu/5wzSxY0lrU/F/ieKswip6MXZO
tM1QZU7jSPRrS/PeJ3hXLHZug5u78dVBTms3eeD+pDW4LbQeDQPMajVOImAFzIGc
JBpqks59FeC/Ox3EYAO6tQzKeziX9Dg+cEU5LjdNTMIapHxa1UAnWXXwrFDqggZi
r2QFGCgXflVcQ0p0fmnsiKfe89Yt/UEcL9uuP/+8jBO9fJTyMp7PfvR5PwY/sOKc
f89+R+KNed/1l/hyC7JbNdw9kDYXRXeBM/mDWVx5VuQ3TSDLLwyaa7cg8BkLVtHt
CG0puUzSbHbVrpyE7ooOCebr0ms4mZjOzg7CHpdjt5pkLccYRwDnVX+ixkAUHnx8
yPiGZ9UIyPZ9j7kCmoowqNAEcetVGVF7jAe/jExiPLryfMHf/cjafgOEBXzHrei9
KRHUCNE3JvJ/ocX1bJ8olwfJxe72fxQb3qzajwOO3bUyOrB0PyQUPo6kHaTnEsBJ
R24kIfjpLKScEcl4umoLrWl7/vYQNZxwMvGznwjBrBtomSw0fUY1Jxkx2E8ceSEm
kiZoBBAkCVk8nxvuvTqppbQzKCgdqPVh7gJR/XssAsqvUXKWaZgnSSl9i7JXxEIa
dfiS1KCJIdgjZ8IACEffIKLt48N1HUpJAN1pAeKMPti3NKzJxNAwYHzZ9S03fSrO
9cMOOh84t4EuCMyiewV8bDaORvI9UCztcTL2RwLOI3WyibkUpU2a2WkD6PpGt/Ol
ZVk1JdFBXtTa3laC0PM7b/EmFTcLbZpTJo2MK74h4hOjBmFrVKe4Gu5VTEO4iADc
YfI+2ESuonFwuZwRS68b5RFIEUgEgaPaYGlnbQpWXtTr7SN9kPJ2sPgocFAtNJAL
UJI4uvscf+75hDyDI7SFgVmN6apDxePfWpSZI2UFXZR/LyfQ0utJIY9ny+BoF+Vs
Hv6lahlWbhAOtZt/5rkEe5KoNJd1PcckwlJO6YgfgupEcSpZheYHKTiVDi3qz6YV
9dRVFDvjMC9jERAIivbJklxEvdHlS9HAyQvIUtZYlYtMaDpcCDeG3AYUKrlf/m1E
/GXt+vsqepft7MU/O0mgG393ZTXpd75ry0hIvu5GnpA00oJtwHGmgrLigdVH2MTy
DdFqf5Y8HdsNzA1D2skcs/2HTW6qRQi0qiSGp+C6AHiXzgEYx/b1AGTWqgIz4mot
506jjRMm8zORd16KXiRN3jmF2yVpiO6afnXADeFvTAVe5nfubZlJsSoI/fgy8TQy
2HY2/iknXn6nnpse2UoHu/tHzpNNgmlSZ0K3vgBXG094HMyCfG9h0ySXznETXVhj
NN+rap07+rWUQqOXtUGOcPZM7UlpEcUmVDmWt4YXPq0dUC7RUb5/2ApXTWsF1nqd
8EDUXg3fSs6fV+Y5y9xyXaku+Ga5bNBEmyMJHSgV74W/DtHSQuFQBdAPOozzdE8s
IjYNhoZwQxTmGAkRQWiWxzEK2vI7q4mdhaeU+R8s/aLME9idILSiP963dK/AY90N
zIjbJIXApsZ5oXauJa3bINFps+OhakBJeUx5Nc3AmjpHEcUgATnZTqmYUdm6mtWu
mLNS/Uuou0TPeqzZcdfZlUEZ0acEMsR/KLr8zg54up4KVG+zcig2RE67gHvqZEOp
gHfAHGjztYE2VNHhY9QyqOFWwk7e3/hf6kduZBgak2uh9MvK9QGqhWO+2hOAplQf
rfXZHJ/n+GUxdHFMOpusmOu+dJrAuikAxGBfsO49G6UewMXEmEDk4URu2IBzBtO9
W0zHAyzOR9yf8XTnWlIOG2MJlS2msyQR+PD1kLvtaa6S5DI6IbEOOqwLpIAuWFIj
3Tltfhgpw2xmwEYevY6S4lXLyVZ1mO0iOMjNxK7sEY8bOCrUppUgmKe2VSwTs7SG
Qbz+YFhJlgjV8H+jtM/4L60XbYZSiTrEV5TeVMhJzvg4zrghJNEEJpoMmTMGYBrq
GC/5bnWJBq6qF8gRa8iCm4Pv7HZ1cEbYAG2gG2/MHoWZjSB+MX8Sb47ig+dvDn54
xgttc3gn8xOB5c09rt4DN7wbmkexOzfiqTPNodQ4eRWMf6Wnn34Mh+KwM+aXNQ2d
Cb6LXh5fSWv5jI0HULLN/NPLQ76sHtJI8ZO7ubPwyoyre4w/2cqh2qi7RThr4bCT
wyTs7uOwMgBMaYftZihDmj0bZOMkPAnaciLDDxD7/T6cVVAAweLQH/9E6oW0wxgI
vN6+pYQVSwMAt+SNIOHGotdYyFRC+S+rtMz8d4GuE6yrwKZqsgd5OprqqxTljxin
zyti3LDKjJDIW6dhjGrM4Ceh++7+9T9q/0ygl4TP5kSf930JMGtgiNikQzoVzIum
Zz8sL1zlFhWW/N/kaiDIPspOM8s672dL66L96t47mvLU8YbazwFJ3YbWDjiKfQvT
fPKK769y1MfbdlEIhnLEX3DVxtiUR+SMXExLAV7B263H7v4htZ9ObtsXKKjFTXEF
NMZ3zbYJJ04hpdUXAAwM9iFOA4fbyBJO5u0bm6W8MZaqVfhH8pra4vsKL6l1IzqY
zzP/Q+umZqR2N4QFX2hU60GsnkrlX6m8t2N1UX+SFjsvOqXhP8YQwLbOTZ5VXEpI
Y8bxrIv+HxbWb/fVZpPDlZtPRWjpWi7r2iH1cgtqjuAYEsiKRuJpKurqPu8WpG7d
Ufca16kQrqARMnXdZOBjjij8grf93/EfDiHcUlOb4oLHSBItraCqGe2OR+osCU+k
sPsMU7OFgG/x4gbpMe20atB9chFCP2p2BFH/QbkMRZsqX0u4ec+/p1USsWVGxhjp
XJgfxvOA1vZXRSgOMTP5zpWiUvjKQCNbnmEQ6o4njhT0pwjh8LGbt90c033cBUwO
kAIlX8467eAoUukO5YsS04xILEPPjWsvZus6XAHQYlim/F4HVGqAXyBwS/6ADouD
T+Ygme65XwdbezKPq0GTQphbRb64FjqkWkpn4/hzJCUv7Uh40ZzYBCpAUvy3+p65
9hjwdYKyhZ3gaAOvD5hP0SA7nT5QhE6CQutTC9WHlbsnnNNlw6ntI4AKI6L2QHF9
PWIUYkax7ScD5sjTqp7Fkv3xoAefJa4MfTW7af1xWwSJMfgv1xkF/DszxjdYL+C9
SMzjMSwLLFhabrragGzBk/b1/0rmlFm2RsGXqdAIgwOs9ko6ITsUzeL0jnv2TQau
IHQRUZvgZAuKuzSKqvYeUt7MOYCM9qHP7ETh8TJ2QIQ3oM4WQBS6gjPPe5PjmDKK
7LkCshJA1fLy8iiNbrhqxvFVZdB6/VKbLiU7GcvDcnTV2ve8fKwrZzfINC1PNNa4
ykLWgUQ2rh/gdLmLzUEJdG5/hUppyrfQA2U/l4Ky2XD/LVshJybevt8HBJcr2Msb
GRUa8iaRR7Ej862ILXG67QhfDOrGnKT4Ev0ePyCY5/EAY8Cc5zPWD+4RCe+DqTRS
qJpuRT5La2/Pojjje2iq+YLSxPh9KOBgrFdA1Nlyk2sTdCqZh91pRajjA+H2jTSF
vPmRgcvVF6bUzgpSZzKBqtcY8TBowJHdADKUxY/MWgdAbe9nffvIDUvqKQUaMXou
MOAB3a5dHtz7nM7eDjyxCLSyPo2cFXO9OwqzcWGvN+R/+MRIm+MbokktQPBVys59
1Yc1/EvhHZ8IlH2AnB16rfYgFHaWEUQ+Geb8cAUpfD8NYmNYl+8UaulqFFwSKJQ5
bwQWVtzhp0oclrVsK8sZnXOcQrvw5CeISNJYNntTdC9vJt/I+vwGNwSg5CZsJ5q+
JpWvPt1h4O+x6npcsBysUF2GVQ7wj5VmnLxWJGyaZ8PTEQoEKyPTFarQFv2X9SoZ
h5icIiwWeiflq7wes9/hWjP03uLmlrwUTDu/rMcHPCjtf/aIKodKLRF1pFLBJczE
FIsezHZuy5TLv0Td+uSva0aHVIdtaWt/d6vsjqTDhGGmmz3NeEqhGxXzNqc8H44+
ase1O8tlJW7AkbvZh6qVvykEJCrMPdaXWTy+WYVmr4G7KomPIod/4ap09ABfB12L
+0AIJH+hQUF6Z5/zK2i3SUZvhsbYSEyGiWxMliLfc5SvGXF7dJiqW8Q/N6JTAOJk
uAvOGXrDWlz5JdH4RkoFxe0oQqXyrca5S8CiOSyA4t7F+caHrMz/U9L4d7Icp0C0
GeDbh0O91bQvoycrHhw2t524Q11J7mDe5dvRgNPVKcGwvzzXMv9EPOA8aie0jwOV
oO9DDC8C1Es8tRtY9M+xjuhc4QJ9R6RXXdOimHuZxHvhApCbz70k3gW0oZX8fE+r
2iFAAW63cszAgm+ZEeWuD3tkWhSWi8tyiKUJIr6D3S34M9f1SQqJOle7mtW3odiV
L9Dhele9JCYz8o3MFZr/mWiBGIzcQuySEF+ON6PIJwuCKOHXkq0ak4Cw2Wtkiegc
2MLbu9vneyGw0vM9ZyLiYImt7j32BhW+rcDbnk04AvlhRCsMyF2fwNfOMqzXsSp2
Lm3igUJ4tgGrnRa11Ju0USxrdw0hOQrZqf+lz3TZSngOSZVUR5vncAf88m9hTpEt
JGlYLsmcV32/+IIwoLYk/LN/VvvBthGwNh87oHuTrRL75VjG8kFn0Yi/28yncHo4
h4vSjQyEv+dQ28Ohkz27NuQ2P3ywKGVWbU2qoHkohYR18tqH3kKzYsvRbnBIl3Ns
Ru1ao1CF+FJnLB8/w6eOxqzMxkC33xJNbyRApzZ8eqOBOPkyrLpGh0/yBqwGmeS8
ucfVIpJeKZszuyHRMR9cIm9BPVO0BD6+zD58Cl2Gd+292pRKI8mfVwGLAZKpDz+x
pBBqyakIQdqA32n6JWxXYEtXPlV2IJGd484kmmVKGDjQvWf2qcE5BZbAj1xQqb/N
5WpXG/FQOqiibFZeQS1rhQ0erJBOnuHlhryInnTN/vqolHv+LGU948jaM9YXoC+A
n7IZ7tWg70pRjDpAXSBzSRMZoeZHs/j3YgRwKogCPOaUj4o46H75+l6ttp691uje
Hz22ysD/bz5Q/0PQdTtfwUt5uo4k3ZTCnvF3pZBySoqwmmWOlHd0BSRXHkUCGLTr
SsSdpuR72CDPIRRv5jbk2gLRemlpTvBUtPRL9vuXD43c30tircNYXgyGbAjzMHxm
TjIjU41w1i0jvJqxrgM+Ib96DsJ9YDelFQCetoV1dZNO+ROJKsFlYDj0+IYozNha
RllLISX1WOpA0Xl2nyXEqS7/ftyzBgI/8Z2cBr43ItWf6YyRvXoNMgce5mpoY9X3
OlGY/6VfDRFQS2W5G3fcFSIaHBKFphuKuCsvjEo489TXix0hfTr70iUSem04Y/X9
j0Q1Uwz+TD3FrsndwHSrvH7JsPVLNjqRU5/JgdfjrI/PcfnYwXrOwZPwsPJXZ3XH
Fkh4gZ+xjJPgV4MCFZoHJarj/tcGso1dFqHtxzDcQJYcV7iKIt+eQGY+SQuqv5fH
texWOUH7SliIBY3CnO5jTZWTDEIvUHYnb3jh4umLwf0yEoaCVvyjLU8PCYYtlY+Q
9/XhKUwzESukLHz4EPPyJC1w07hPT67iN20VgUlZKh91YDR21YaYMK/aiuAQACu4
Yo6K5n/0+gghjC8eh67W8H6ze4L4E9qKUF2LPc0avMvm5xebOR1cExAm3BQ+mSeC
rSGwyESvtkSNEiGPTTQfDPX4dDXS3ZRvJ8I2U5xgkAMtRqY7ohaTJlawjRQDxWXn
5KFMz49yqs8E9He7uRbmq6SUZrvkKNRn2Ie/dzf+aPLHlVtJOays2BpefqIuBLBH
/wPcXAPPPBJbsiOkO2Ew7k+kJDSMfjMRoZsPNFh6usDSIMu56IxO+l0on46FLcUh
tHxQ+nqWOW6MsWh5UzUSWT6vxsjYScFEGHQiZadDkDgkXEFAjTKY6LIJdIJWrJ1Y
HHA96RAVSYGeSLrSa0d4rM7ZJCQ1ErG7VdwW2UdHwwtcDU9E+u64GitIkxfmHVYy
OArqfDr+Uz6ZElkxG1SCXJXojRmKio2pvTl7UXaxaPnDpMZVGnZa1lXJckw4Z4Nq
TwphETP0pLZuVBLS9ZbhhwPsuL1P+ZTq6xtHpMAauuGmyVHtmedlqXTeoGWZMO0h
pYTM1m9URM2eTjs3PnyW573hMvq8XqBfhD6PwlmBK66IPs0AfQg1ll16n8vsr2o8
lMIn9ZGliv7tkwe6bF8vGjCrn/3s+bhnO3+Oj64pRkjcbwooaB6Rwf4nYycEigwy
D7Wv3yJGrtchshVgE/GeuBrndorodD2vNE2zNEVYaq4cIMNt0PjZXQ4HjVeprCZA
tJnRG6kVDUspUiZ83vm8MjiFQzSrbkVdHWmWG1nmY7MiVTIBXA+PmsQoG3WwUx0l
LCZJ7WAKh8zbpe5kHesMsQbah+2H7Bxk0saV96NevcxTSFC/OMgxKrdvsH6tSYTL
W4omTMzkVSfioiR9p1EQOlRwlvm9Q2dJGMwBk+ijSDT4ACdEds/F8rINNWM7/DgC
66MQLNIyyhT1VJXUVHiiwCRKU2VzT+KKuvPyK8Qkq3Ncn98VGLVnASPSkFmk5nGu
SDKLQEDW/V8lKOJXyDiu0wfudK1ebQf/ucK5Yj7aXounVK8+OSETzItoGwuWAoyF
aJQdj+VdlRCN0HnXnXU0m84LYTafAiAh9LjkczafFLfX4yMAIoqjsL1XM4XJwDW0
lFFmp7BlQva7+tbcChI5cp1r94H84ig78cFsIPGj0/abdbDg+xDY9WmiZ+OTZ4RF
YxoBCfeaLwG6rKktzA60/m+KDuLJDEjG0coM3e93EmB/D8a1wdq8WSDe9K9nxjkt
2WbcVKTKDhFurG5WlHYqDRhuFQW1byi20ExgXoXaZBHH6cCrjQkydS+SJK5Qm09E
ZnTMD6Vf2PaiiVVidaY6mLJePy4TYJBy5pIzFeWzO+VpCCffU8nwapoylExVNlGr
Oc6/cR1LbCfW1GOUtvvVgPMpOJ/yq4YeIq2Z/J0F1Xp600KPS/X3QGvRfwz/74pO
r25mpSk4ARV/hD6po3bZAc+mKRV+QYyi3EnEkTjVzLCKSCCjhxASmWE+z2GejvGt
MHNEfFOKiKQj3eryDlJ3psn38yTnyXqqZtTLZEr6/bzYKq0M6KS3oauAC02LFUet
xeN/YOQ1MbeNAixeaDo4TAkq7ftLlH597Ck/zOmMsUC9dGaNiDre/Nr59TRvicdu
ElcrqXpm8XpSv+vIWrH07CEScLME0zlCvmXeGFQ8opStiTcBeSKWBQiGedkqwxq/
Mbefeb6Nu5fzFFRI9lb9dsNu9nNh5DWRrTZ+ESSCJBP5O9t1UbIX+xDKebF85yKk
qmCo/GUNWnRa4PzZJtuX61dRk55oCsvv6V4FWoAo5o3DsHl//rst4p66l7uwwMnK
xu/8+6W48zGqQOTMhmP9RjXh+LCeamNh1ubdPpH8I/4SJBGxqzk8BQcZucboxbLh
8eRlkzYTJMCo5phbSi3FMRcS24aK+MXbue1wPxViqUN77r7Ezv3z9w0HYGAF9nPc
lgBExMTjIxcK92KwSHSnjLMf+gKApn/oYs3DizmKJ+NaFimpxnSJmXbD3TGY2Q8u
iTKnQA3jpcHINu5Fbq5dPDvwgBgtq6rydBEZDr+LcgX4NCdxMK1vU3DkR8xOVuKf
ZGb6OfbAbl1MA3AE4FZBDraGvU8mOyfikKLi00pPFpzPkWyfk21CYDbWREldXYij
+eMp8giBX+xnrhpaTffRNM4ZBn35HCOT/vGZv4NeQciPQLQ2sYyaEOcl5rTTjROQ
X8PAaK50mPKca8GovQPyMkJGW9LobuCMmDLoKXfsTjNQiyajRJLKptpKgAcRV5ha
VvjcEmLoeSajSkvvWGLvfqgmeSsb8SViHl3qyczR7p+dTXT+kLRODgIy8U/Zg/AY
4kU6D7TGBWYN7+HFcV39IxG1P4bVZxQW+HClDdWS4MMuGxRQppR5JCgGwTNystnj
IKOcXLPSB65Z5m2RSqw/QwNSuTXboxK8iLwiTMimfh444eyXf90Qqkv2MCyWRQdS
2WExsiWpnaqWDETgk1ZytQFfxL+VczFKCeZGledlOVL1maTl0VQVr2TfRHZo8thB
we2IjgbofdYhup5fF1FoiU2oc8+Rzy4rq2qP1+FiBahXQHN1UJTo97SCoicUUzTO
+WOJ3c/jnzqEwXmAlC9E+I/+iH0PTMGawUcxtdxco0MPk7xe+FImWbY82dFNQFTe
NKdBkvY9jiM3f4aSwMj14WQjVVi/T3HRW4MlqemRTHA02fzUoQs9VN/usSrU8nmX
o1jRCVInzKQHsSzFkUjorVUIkmjgEK0E8UACh9uas+94qnePX6XHrFkRF/rPF4Op
uWbdY2KwIALAT+v06rI8QijDEz9r7hPH7S1K4inoWyeZOOcUjWc53+MiTBwGi7ml
3Rf8AmZfZJqSvCl0SvVMDDhuzmWsOeuHcHkYLirKs7uhRb47DV/K1YoG1NngqkDn
FcNyhgcnUHk5H18oL16QDIvLAP+cnunV5c3yrqLMY1FaBpPYbx2fMx8+BkBdZY9Q
J5f7ECziPTvPcKe6auf+CBorptPIm4k8yf/SKDVNQRnyMio48UlSzAE9L1LiHSCI
uryG8lRsLv2OJETjl9Me0MGGozb9wq2HArTKlfBlbIl+QvM1QuYenjQOWf/3+c1s
UAsyx7FnfTSL2aIjCceiM+w6LzA3ANVtZHjazlqkFOtEbkrRgFEafQOSfQj7wWuW
bEIfZBhCaXIPA5cyPFC7Ex5yWbdEqZGsfGPWLuz4J69+lfFjo65JpLfxZHcrVQRI
h5Bep+OLHMPEWrAgm0TdqqDXqloHJwFYZGyXJMafAMm0MgnoTMnh4NdODLiMgfpB
pDdEPwLU79CTISED7dMXerrmntGuap5JwmKvzCr7+a/7TS2k+qdMufzf5x03iOYn
rl7BwNh9Jqla9gh317pD5et9aYdF2mG1yE3cpGkDGF0uA2xMMxRbox2yU3DDpFGF
Ye1vN0eIavQGTM+hNdQo5ABYchIISR2wqssdp/Lx7DFmBxhkAJPF2UgoV9tRfN+D
Wrgvoh3zaDsvSrYmQCW/Y+Z4m6Ee/+8jdRqVEXF1vHdy6EXVhOcQCHjZ/96XrmM1
TSedLL1GsUl2bjvfAheRImiqT7jGUmMHQU/56dgRWFpfNmHd4kA2KyyKO5jVMjy1
FUv359QX2+1QWJgazS+jD+wmCkbHVVpd9605JR6n7UC29FFwnpY7Wk5WIkXIoiyQ
Is7zxOfhN6wS3WCkj8Jowt9z8NuKkB5OJ5g9Sj981+CbubXT7jqBrgY8Plao9S99
B9B/+HnMbEnnn6MAcgkqRS3cxdR7CmWIheum2TJ0MyMoUIdIyMUYsqh9eKaj7b7x
GucnI4PLSa2drnxZ6MX+HBCr3plfGJSuwmsNfL85DDsgLEGQbJqMUlxJd9YXkRZd
oLehAKbqQ+EmOPi3dXsj/ZzCnJW8NFFUHTbydQWzJASXCiaJ8XDYayYNk1rbqvts
JCwjBiOc4aso52EfwZ2Jc4TSQNVlqR5q/dcSMFD7eRUsdV8yUR1C6FRYhInTyvYC
eAegXSQ1knSzP0p3TcdllwUNgpdynSIRYkNMoGSvfZwQdxtMVXBRO1Fkd3MiBuz+
K+rlxpaS4o+uxZt3cAF8DQFsCli9h1ADLfZ8DKarsyYEZl1D7GL64dpXndKisQnb
LPLPTD38Jrd650BWAOioQQKeIzmz7w/Uh1MLyoD2yuuqn1eU3mknw7Dd4Zg5ompz
M4ulJ4hkqvqeEv6MYBvG3dn9zN8HzUPfhxdn9WcG11KlP8YsO70XKp3BlX3Obfct
0C8CqUp5MYf+wP2naslS27E1Yi6A72xb2EZLFZ3fv85PfZtsHr1BeY2XRFvwteAK
e2FryYNi/GpG6HQAL3co1LzRIxnCPPOdea8kzGG3+DnuXrDFVUSWvoURRCN41KUZ
HXT9lmKc5kLG/5aGV5m3vf7pZG4lc2OR3Owj/0LnVX5sz0eu7rxMvRVWxVYTr7Hm
Y+u3xs6gqxmP9lBeV84tcjvVZAm12og5Vk6cyDgeiUbFK5eQnpeg/EWeJLMFKKvJ
UyKojUiv4/KTyNr/6I55JBSMhxW+AvFIYs7s1U1pN/SNtIMAs/6l9oc0g+GYh6IK
CP8xdxHFKxgAjQavw0Gn2/JdJPWtXp7u1wBNeJmdHr8c7mWd5txb37QyHjicx/vH
43hVAMMXBWa2XMoughn6xIIRlMLnomADtu2ZM7ZVX9mliEGo0vOzuQ1nUBiqwb4E
dyXW8OCeB7zIGO5KjCD5Uuy4qj8o8ZNr5CM0Xs5AiaJE0j84ZB/4Yx2pGhZnyTh1
1QC+L6jRYTpsjf5DWfiyPtnd6BPdzEHSXq0ZHQwC23elSzi7UD+uHqvn2ytWww5w
aT23r67mEyoGkOMa6IxMmRW9asbeRwlvcb9l3Q2VIQOocTmx/R3fDwY5DgMmxPtb
9QJ90H6t3sm0KIDBd3byQ0uEKdKCDY8cBeMiaT10KlInzbcO42yzRG/Y/tZwYnwi
LU88rJaQaJrPg3w5AQN+qX9NIfZyjceEXBLvZHpG5s1Poefc0e/EPKLIpttDSXRA
/zuJ9qX86SE6Pt1Tm/1g95tgZtkuDs7AyvLk6U3C05aSuGUG0bnpDTee+inA0ucT
DzA4+60H5m4ZEKcmgtd5YaaplzppA/7Ev93NfatkK8UGTh/Kme8u2eYszwgQq295
lpat0cL/pRx6a3gowOe/EFzaQ2+twAeeM1nG4NL4nyzWlPnQ6CXxLVbzbX9sewaX
Ra/dLFbtvfEHYcCKwduevQi3BAnKMEJgnBeKPEmA/CuthqfBXl/Ytp40KXVZeC0Z
HlQ4c3EsSsUaECOgMic+LULijK5HkF24QCcg/jzaCme7Zrpj0NRMoQlkYHLIL53p
8QOG5TzWvlpL9SOaBDC0nAUatXFmK9IqPRm+mXHs1IlA2lPEgJuunU/RhS0d5LzN
gTv6/AMkKTDxCftKVXbzJzv6s5dPihMh5zGLLfvPSlTw87upXC9z6GB9npMx740Q
Ho58ZpYUp1nr6Ege/eyq48Wg+Pf0oa3GzGuPx7twLv8rUKfZrcrNN2ay7nw/kybP
4ZioFnFfXCdyFZIXdLJySxKm3k1OOrvl3FKOvY7j/mslPonkTUATm4/Su+n+4gv6
yCeRapxPfzNO79F0VCmIxC7xDUfLHAPlveDSENW1ljpByf49ArG1L3CJWw+dlVRm
crpCXDnGYMJUDXxkG4hymfT40X3d6iCX2LmOMSH5SyuppwBFrplpZ84jS3fhsygO
KsNSmbHPdsIQ7z2/iBNPdUnho9/6ESNQlT562rbM4em4CWrs0AbAil0s6g0JAjk+
wzmVC+q3EA5QTTG6J5jrCtageXfSq/u0Jh7T7BNWyGEMBZcxKVUTaEBJdoNYcIPr
lvnVsXbw1VWNzWL4b/499nSamd0CH4OobLVYpRSKkZK6myHH5JiRmCQU154vMhMi
cH7IO0qmfsaWrNH3GRj7xD5bnVAaXQQCMIN2TGcnwgQ1bB6Y0wXPVi72RvZnVYTG
mJCByCmYedJvrGOZzyK/9jwsf+T+jqH3Ah5qmrONx9qjm/FkY2x1Xd4DGAjws6q/
LmZoy5TqXha9+aEWzBQVr+IriU8/OYela1ub99xjlLTomzfoY0gA4gP8aIxTszcD
ebhF1OJguZKN6dFFY2+NdtvFtGtF0QjaKID38xkXYy4ywVXIi418eK/WljtFwOPz
r3idCYxl4/LTwJmgZ2IJgCbAhOhJcRxTYAN2253dLEA4PvfLWhEef2KwQX0KSsrM
Tr5gbsw0XfoaKCLU1rsQNxy+Lc2rz7nb6NtF1xYhOMvWSeCoEfLL34kd28TKfBAV
dDq7NfUgd7lArxGowS8+eEFktvnWEn0qmlcdpzs9ZTfNCuN1YTCibPd2RSeeFaGf
GGmHp1b8sHUashiEDcN7hXpAatIKVRLuh1tnNFhP6BFoePOGibA3JgLPpHh38wLZ
D159INGgBDgLmyC7aA7g6THE5R4Kw9prZAjCr9RzqTD42xbLpAoIgwz7SRyKlQus
Cbwh5f4eThQ553eQuRJ4g4fiw3zdzMtYk+O1hokgsDeB0j/IvN6l1VH/8YBBVrMC
94pT/RaqVHS8dDxbs7rE35YrEKfY0bU9eXSFqbDvQw42V3QAXCUJLVUyQoHHMoNy
HbaQfraPVO9uE/SaoFyHbxrgFpwtzpl+/YoR7d0mi+F94sF30RVUBPqrjPh7IUkU
DyfgtcwJVkNLq+UACLHnmIuSdFbUQvhIqb/F7Ij0NPqNo4vAktreT9WaEtdfQ24c
cRnydbFa2/0CWVlyCPUTEuER0HcknaxPVCAp3twBJLPjk70yJJfc3MfbGHGpLoMc
DKZKxTK1J/KDNnSZqg7iqTcZGtSHHPSk+qsWa0tGuIaFMmkuM78ezxnd/EjvaxAt
NYeNiWsspsRIGinkAbiCN8fIQCFrn6P1wUVwOGsAGYHznO4+QNaL42mMnDOq7ftD
aOt3jY/wj9fqmnHXQnEwvdwhrvINeI/uA1ErDutIlyfKmKskng5w+KEQpaebhyHr
dCnQYxnBKTFx3kIU0zt2qX4QLdIrpWMebKu+obDQ0aQCniT63M67EY9np7sFqxPe
tGwoCAdHGxF0m3SWyzdsYqGS0IQF8DP5D0CZzoW9wMj0chGnyupf51HvnHWp99M9
pHKSgPklyxn9QDzSEzxRQ2y02Zq+OkEwFjXDQmESjFvoeFVdbKJO6Mlr/umJOtGs
7AYNk46FavILkC/XhCC1UhlWV11VnrFTwnJHj4NZSRkE6O2oLK7LTuUVUxpnwYcO
a3mwiXhFEKAOg87KmVuZmDAKhAoE6y/Ci2b/0ilrORL3It71vQXkb6aiLxb9iIgB
8Esh5JxAgong9E+7AeYFF8YUod3I6kvwtC9xQ5Fz3wz0m9NqxeOXjM1o4mxczv4n
MjRth+FU9Shf3wxiPlfGf2GcYjtxG8jOzLb0tGXY6ntkA51XAyGB+v6TgWPZKsuG
iHZy4q54kcQfZmN550vKOoFZKKDT0XXEvm4M94i9m3puDfLgO8Suby6rwwqVWvKT
8Pow5WtJA3hDEJbgwaku1xUz0WODhsS+I8KROpBFffcZzGOLDfq+1Fz+DNTTF/S7
lzsbAs30ZmGI1pQKAye/6LCp+ihjTY/ztIa3DsDPKsPBs8WtJUNx0QI/J1kbfYst
7LabGpjjh+Nwo2+VDy5C/OjqdoUeudpGCtG6EiHdVX4Gt1R3fSiQ7I99BPHrMQ+T
MdXY65KYXSNHr9uPZ8iCOIyBXVXxuedSBD5diemk8PuxkaSUONji4+tFZkqtcIcK
3+sh5uqcc3h4sh0CQsO6Dro4KBwBfrXU/5vmnu+b0aN8hY7iHcVrWrqlO+he3x+7
dWqvnIVGSBM/s8HEpteVeIyapeoqKq38qc7xQlF3jhd6sAQ72NHq/zzDzzbR7nwt
Hf0nu12J0tQrkhtd3O9CA4yTJuZXQgaNPhcK3nx8EvxyNgpatCoNFsx24jEkYgIa
zksN5tVw/oPgk0nUeu6jOJ+xaQTLIGZjpT0v/zRkOqft63fc6Q6kS+eX2+7nm8IK
+e7qJzHDtBfFH58B1t8t1bSK5iIfJhT2e6PMVUi3TSxuJo+ArQ2u3BPTSduCopEq
3GJgcB/fwys6RHCVsnDUi63zsyj35oPU/0docnrnU5009jZZqpJd1e2y3NwzdKIy
FhU7TG5b3JKRklT8OGoSsTf+IlWCp2tluOlRzkghUP5b4i6i950unBFjB0xYFOcU
/JPhCf12FOhhPKsDh1BTcFJRmkImPRRPYQjpNU7Gs5NTz8EtnzTCn3GDKwz5Q+jL
vXglEn+hfmT7eQ+S+rWKrFwI8UVNkFhB4eD9zJn6+IUWS4+s6MZ5U4qA23lvlzXV
hJdz2CCnAlJYnU07uKGdbXtCTNC8j1jlu5EI96fHBWlIaWMHjo4QEsHe+jhwBT0p
jujMMCv7X2dSiIF1ubo+naF3nRyPTTxkbrfCNuh1Tz0sKx6e/1w31MMsIfkOb4fR
CS/AsCKoRk+h/vD/A/grDmmWeIWn40/aONuWFDm/iLx+nFBAFwo9E6LdNJr6wTt5
ggPpBXSxk3CQpwD7B19gf5QxFd1AswgPHFfnC4KughpQ3lHYBRIV7LIx8N6LapVV
T2f+k4TS6W9fXl6XhrreiLckK4AMp0ntRwvsNtCfx7jC0i+3Vbi79AZ1rKw2nSaw
JfpWvGI7cbbtp9nrMSb/EsZUPPUtyQ7n7jJ30E9Vct/0w5hUlWjmqGG8QUhiAg3m
2zL70OJ/gceyD7tTeeCaDnViylcS99i7eoWuIsYAbIvVzCzDt56w82fhSjdxpg/3
w0z8JX7iTginkxo+mwvV3bGvD17Nr+piNbnSVav06qyOCK1TUUXdWMjlAds8+WlE
+OrEXqHo3citFoa4p8skapR0qhG1OtJiLl6oeJKBhnDYgm+9mFCwnQgQMvvun7H4
hASHaW8of0KMJgOUUbX4Bhue/gHWPmx37uuG4eI24GNYaTvvIt9d746ULqMm7Gf4
IzTSQe8EjJXAOoDr1K/sxmitoThaUoS426Dr4grqLqetVZkaSrkkQ9JcsvJuaA1t
mVzWGq76l/D4+XcJ2aI15Bzf0yv+OQriD60Y6rxSLEB+1GBs6rooc0m0vflTqlaS
r0QGLOU4QiFueK2nHh8yIf/fdzCj28WbgXZGmn7XjZoH10u81Y1rYHdusIF6D1Io
pBc2zxZq91+pDTcTh1q/P/3Y/kjlpLJ1ymlUfUGiLBppPzetJM2/uwu0p+WpQRs/
koXDCgMkNAqlzn7GYqqkq70bnBRzUts3+G59mrMaMezZUjN7pQKs7TWoAidJvCmh
+D+eIvyRVEzAM7Khu+00NTy34yHkzQ43Rtw30s6qZn+TFHfxxpCTrwsp9tW5EU7U
pgXL7p9o0P+5EBVArA2vUzNuF20JRxI3L/sgF7LSrmDQPI9v7tKqpXZJusCwOLlk
aJMoGQ2fEbRcsZd9srli+ruvq8oz1lGl2MrTokf1VjYqfiGh7qy7SwkCJ/zhjCbd
MpYWv93qnTFHj1IJrsM6C+jgRCXBjVfh4REVo6iNYyKxFzppIughs3rgUGmzGYPm
HYovw0B+6GuHv6Em5/cflJ1ebHRbrjUCg2XV56YpceEJ2ZMiWIroeMh6RSZHub65
r08aRdBNKgqaVVp5WvPMlyA/YDM/OVwj8Z1g46kW7aadCrNfroVj4Ba73IWHwyFL
YXIZy7JOC1PqrrurbkmmRDehpcIf7oPSHkAvsOBIGIUlKv25/ilNDh77GSOAXxMr
zd0B0yQL8yA/KGt0J95wlmhfNCWB82kyNmlpbCdgmjUdL/CJ5cpHsD7tb9wUkXSd
6eim1HsemdMDzee2Hei6Wd5AwBxwlyTSgfEEDpimBinQyOOmOKmSriNo1X0Z8Dfp
lDux29jZOlrWon5j/sx7RjyoPwVAag1eoK9C5QObVMmtM4yV2GbvXHqhXFrCjlUK
D/PZtRZq4PMkLnW5pmxmooQh6ORpbaUmW+0YF0ShMty27mqrFteJbHA+R2MgbE1o
qBotJLv6nxYYVHv6thhnen/+N7CiqpmY5KwCB5CGaIUeADrFtt/911AWRaRsuFqN
OkUdcREzFxVrUyrhxCWwuD3wSvSThAB3GUV06WdvTDn6w4Iqu+RpIXAFQZFVbPkN
5mLTUG/BG9lLGL4dMvKd/PQ36qd4kHzciVDkSWT/tI68l0bn+88+wY3KdJFxTsIG
Ok+X/whqIHbrSwWClrrHmwf0DfmRQLGTBWcMJupscEVH9cLeD31x+bMxGODZUlgG
F9QTDHquC56WfX3VaiOYgHxYUWZpDKuUTbbGF4boJgQlsA2MkQE9I8QuqIufgvvb
/HWYDxPzX8OSHwK4QsAxZkyDlAjYdE4MItgngod4Yusw/+bB01UzoKFl5FL7eWgg
ME/Hdv0bd1HuPwF68fHkHCDz+jvR/rSzc6Zr1LF90Fh2XrKS6swJfyDOJ4Kwz/6e
caoiCKhxoatHjxCK/5wpIe+bBHRQXxeZujGUb7LOtf9dOLVwkYfoZ1tQq1wnTRRS
TZJld2d8Zq826/+8VAHrVzhNDxFVvrGm4eHobWqyISwLLVNVKswZ0PaYmCHipbII
7DimYgrCnycb/TuCUi6QBA6zWKMe9aCqmsJ0Rk0f+dz8Xcc1MdVRtSkjCU/jxCcH
8CXgyLy1ehsBt/qjA3PyY4jxCSOglLFSvxE8bcU4pptcCpm4PdKdoQt8BR2nnJJm
E3w+iLxHrIM2YJa2XPBRrm63yji32dX2vyFOLtsDE3KbDIZs7BI+U2vhcDwlq2MU
wx1To+nW3z/VaqnrprQOlhyhvxR+p0sT5v4Hz3dh3uEHbT2INLvlXXM+ei2MF7uC
sKzdiKqY+JPbIxVRLcXltZ65gOWFZNzAHDOwBZjLdbPlzWCYqvN4Csb4Q+881AM1
WqhVoocRK+QiSPmRVfP5G/vBOoQWbip9T9fLtM2dNwvkPUWRns2RJMenfWIvOCHc
GMvnw5F23Gy5WPCzMZBHM/pK1qzlB6/wMbuvFXth66SIXCnp4N9up28Su4zEpogz
eF3GQSHNXNiFQOBiceh6hn1P0b6tQoa3lvUGrHGU+v8OWa92sJ9C3OJ2IuE4rp6K
beT/nyFvu8d86Y0tGwKZRg/xpXmxT9zohpCONzqlJ+EvEM80ggTYc3wei8r/TDsI
zluEN4TgX7Be2P0qU2WVAPr7rmA2h5d/v8pQ+0pp9SqUZae5alcCzoOF8SDkk8Ci
+HIOJdgMYiys6NlKXcc9RmpYa+NY+06UoHp3D9j6jqgsIR9DDV+Ay+DRSkYn0QII
hJmyPwf1TU+hfJ6J5Q43htsIwnIydyT56A012Piu8QPnoKQB1lInGsyUhX49pC+Q
xxnZEfV+mumTrhyT0wynaLogbqKufQeUzl6MO2dE7N3vhMOYZ52msBzg/nWiMTnk
58oQuTN5KGvKvbLcvtqYzhWy1wZskSrajDTrSHqYpgp2nOs1DZBVUfmFnAJXQhoo
NSFYTkHMk4uBtqQdDE3Jp6YnZwAgrDQuAS1EfY7CGbnz81AAZ/Cj/9N5Lyllg0RG
puYwUoWBbWReLv61LgMc61B3gI42S3wpemMArH1T/vnHTeHgY4xbvfly7K7kudQH
I99KKR0XRCz9pI9YaLEuShnQqwW7Qoo1LpyAWYDHD5nXTPebx54AeFvtEoXyUgK5
l0u1BU/QzDiBq2lP1AM7rolcKvyL9RHqMn/wmUCnYWcBLRZ4UZRWARB2bTlm7xcZ
NMSE0PFdZqYNB7GlazSWmlzclKL6z5Q8HchjsQET1rKLa/gujBOn2Qjyi8djVyoX
0kVugpfUadBbj4K8I3FcMsuz6ox4SkQGh3Gu8ZWu5HCejeqt2eG7jPt9mFkLiQjt
mGp73GUg8m2fN6Dp3T28Is16crzH5anP4atwYcQeEokhDGUiZKXLAOFl4cvsKVHh
s+5bLf/OdZwPJd/cd8ErDpUQj0egHq5GWgIthmt4u5fA6DMzy5LNK3oXjeyEIFst
Qda7qtE712eenXegf03Leu48WIUQR5oHO7+/Jdcsy9QGJXy1eHNBQTiKqK1eonWO
1EX7X2xxWQF0c0Rt9sTguzM7zk9cFVnsiJrnhJOW/cQ5fUHgzV8mENgsxRc5GjVg
5mC2+yjMOP9dj462SUNmZwGKZvAy1D1mr/JAaF1WuwxFghkcoxluYmN72pFfLAGi
iYjTiqE0Ke3aADPznSlAE5NTV08ffT4UHFvwBzMqoss6VjaJbJU3vtYwzWJiIT6N
ZakhD83yr3yncnI/8ILUNInNllUsFTrwzGUB8HxDAlqNfNQ24TrCEfGjnpqG53mJ
oSHFiXCu50NEBIHqayLfvUhkKz6OLiOpkALE6RFmL8WCmNDW1EEMEH4+dJzsjOi0
UCKVDTM4ObAf59YDR0EroZ0FRqsi6yTuETFwIHbcQtT4k7sF7BRiQ2gmKZAuwmHU
WXlumNiDjJES+KUv0eO7UNq2NtP7tw0VN34exqDhUxGv92342UQsRMMNKUToIx4U
wfvqGo2EQvrQZN8LvqWb6JFDmkv5TJW0ZSv+lsoiuxli/3O10mHa0AoxrerdPvLr
ngEMoQIiI/zNhzDplY8qP4xTjz4uMDh+0I+SmiVaulSB7TYMWqZlWhJuYmIYAV7n
Qrqfy3/wAbIMa93KCxX86CCapd2Xj95LXTzHbq4X7EE5i9DjWsZZ2jaetXBbzlfO
YL3hq7PhL4D1/PF991zvoDIMzQmQzmCWQfLv9FVptMW7KsuXCxWZljCI1wgkb7s5
eNXhvMMf9925EXQSHDT7OCxappWIVo8c+I/ZmohUEHnyFRGruoPyKFqq2jPU7xvh
Mspy9RK+V3d2U0qI+SNeSLuTGrdUGQDGi+1oFMACJFn8gZ5zsAet2XwJqLm4mWML
/ADg+q70GnDgbSpHmGIvpK0pAZbYiOQltm/FbuBLgRi8i8cfGx6P1c/DxSI6O4b9
pYYDADw/je3N3jQbldSL07hoEQFYPer3O6Siq//mhhy7kNDPtJE35/NpsGKC6ClP
qNj8cLQMcF0J5O6FSaOnmnOtJGUBI+J9eEAJRUJh9q25XmCscP1Pcva3dFlCpnhK
kePpyXtcEv4E3aB+kiNPoiLwS6LplztqFvh2IXE9mRcS+TxSDsqgAZMjt75utee7
XT4g61VSvc4dxh4dca/zJg80tSKqsZLp7YvueoaHoeFZEFfUBBIYNcEklXBJfn9U
jVbu9X7YaqaF4dyE5yPZIMP6BEG4A5GqWFQplcOJZg+Ey1zXwYM7nWqdTsP/1cyS
b1FPSkdk/pPkRHpl6SpjOrJ0KZAuDUU5/ehQMI+by8RWqej0yQpPJI0sH9IjL/aP
O8uKLIzFoFknP1PgCK2AbrO4NMYI6cgIg9RdmPoJscrEXxrXs+ISWjeM6ohLqaLn
/bmpJgI7c41ppNvw1U1Lh0JbDQ6PDMxSxdwyxLW5O6RoX7yeevv0BTSVdQKu1V5M
3PHIaL2LY9SL9hvYTO2hkg3Q9ZV/qhPeh2qeeu1eriWDFzkzzlYDmK2OIOk7Bswi
9m5oz1M+CcP+kZMtUGAnk6J2tVPuFtyYXV5RCkEL0rkeXJXKUJBeiR/6pM2+FBOX
lTIaMQ3X731jDif0Nmo6peZ0QY0oyevt8EquptzV9W+gkt8y4BqUtwqqtsGhSlAS
NIpWGpKOJYChEkBRpkVlcmrYjoPo0gvNB9h3fLAsLvIpd0JOuwGHFAweo40hk2++
9tKKco6aljNlHS7H+vrti5+Mgxy3Y/0UgkiZYDSLuf4hk0XBBLRQXnYzbZqIRt0Z
r7mCS8Y3kQOTiuVh6xDTavYJMH8tk2gGaAj9ycVcKalSjPK0vYp9qS8zKjf1Pe9l
ggKDVW5Jas1Cff3O521f6rQKSGmBo9wqGKQ6XGP+9UQKXZtWHYqGTlY/ssotQwhb
HTXH/5PFrurEipXW8p3f+9L0VCbo5UgPNNMNlvAaoGlupJrO4+yY5pxtEH6QPCwQ
5aL6M6THcMVw/cNydPM1rzC3C6uc7ayRsPlTjejTdbQC15o1xrhxCeH1bS1h34Np
1QuyKu+iWWc1ws+mpUeaPF7bCBBELr9OyMshkavewFnnZMInbW/XbTD3hPLS3ym0
6fCuUGqGJh9/g1DnCcQan++d+1qs4Y6T+yidOHEDHoxPGFAw0YpXNtAPoVzwRR2p
Wp5V9pHhTgx0T+tOPhifP6qD6VUuESAZQPg4cbSg6gMNh+cwGeCLxZyAxUe+j5id
8J49yTSTjPGcBgIbyTNHU5pIYMkmZORkWHc1+T2wcSPhsnvlPqeH7sOG26bui3pF
FXBibq3phYpnT0ruiqtrnpHbne+d0S5OIbciMl9/uA6q44BJmtfCFALK49RroxJq
wgWU3jRrbdsmDshJOvJGBProbvDk/GKK8ERodDtf/1uEkCpvg2gr/1x4/Hzn8dnc
OtRtRuwy7OVo3GRvUabnbVenEdgAh2Ar0Ui5yNSMdcvn8dvndujcPdtS+s9bkJ41
Bkc0AZlf1XVxsk+u4qvarwkh2jM1Tn4rO152Q6EA2dqwg6FF82soDroXbhWldghE
spptVv6dBVMrx36w62a+ZTmS7APHyDTPde9+tWlofYATb/P1orqd7YO56wQvcwyS
+qP7YCWY7LgVu/orUJzowghYZk6TRFo08/o4HDrM3DF1nZrPVon+UHONt0XBHCaU
Pz3z6xfzWN5zBwoqFkTWwnZgEju/fC6aUw2JYsguhNbntN0oGU1MrP4Zol9LKaWF
jdIBEnFLn2hdZa/GXfEis2vst4toBcUOYuE6ZD0Ay9gGXSRrDnuV4CdHInus9chp
a+FwJmFthk5qjS6SCK2KrHloPKctwACIOsd5/W9cHBz/AKlHi65ZtSBl5JN12pAl
3Uhx+DmButYINVlt7W+xof5XYiAMEQHMfstHdUfWHJK6U6lr9+DWWcREm9y+SQ5E
qcMaFiiXWcBC0diOUQPXkl2ZK6RNRM3P7MYWlN8JKUvvqz9GAeV7CRhSahRgyJeF
Mzx6PHa7ViDrcMmQZfvzukk9Gxb6pX28/TG2OBVhLDvPOLBgx/3Z0t4Mfz8gk5eu
LGp+b06EYQiCrR3f9VoXng1273bwfwg06aNT+8HbnUNpzBOql6OVd1c/dZGsMJj5
XDFNoigyhai7LszPFa/n8IybW5/wXqQhruLZL8YP6j/8p9jBsi3h/7dik0Tqb/Uo
rcvtd30zMGnTLgpA3zWZZnixpj/zZZ5Fw4ugiPISpAnW11ZRQEVcrf5hhwXFxIpC
yExm/Mjl22JRFI6k43FNOwklIGKbFlTI9uk26ho69ajws1VMyQfIsovog/+UpIlr
22l7uEX/KPklTp4/3/vRa81HjwZT1J167mIWXrHq233lvVj0dNzG68XYChqA8peb
tnoP2IPM2hpGZhS2IEjwQxtdGvxah/PztmGKMMeCbepsMcMK04oifxgrV4MfS+ZL
Cs9cyvgfYR6vhVLVq01ADz09O/+Nsup3+ehO244zSCqDqdDSx8dcTmTQVolPqkl1
9DIGOm4Ooizaa5NszDnlN8D4K8SArZfJwhHuNdh4kokbEnMnjXcBALUBw+TIbIly
JQoJRyfjfMyjZEu3sstEdBoxdu9NUQWUcAGNdzagHwtoekXmjr96t/eqT12rXLGX
P4xBVZojHFJav4JP5warkMmTTF/oFwo6d6ahh3UN022/QFCule+3a9MMfVwqWRsi
fFYu9wCitmkILIKHJr0L0suzCraf7qsXmj3rcjL7LGcxWDesKdPkfyipAT0+7JCE
yT5d7pGckPjDFztsZvR7wk8hc6E+0SuTbbV/NJeAt85YI8r94rWqrCMljBy0fHay
hJBb0nevypc44/e+byzDtbYD9VPya27pbdoZxu73HyPybQxpuqLFRLIusy4oOsxg
I7u9st5Tmq7fzmPOwDSgS7qaKXgwDrvmooYF24ROZpvyZczXCI+bWsMYrGBm3+YF
yBpm8SbX7xHnz9NqLv0qmuCuqzt6qfA7lBBU/lalhxGWaao0MdqmvormCouTTj5S
jIRVa5W/HtEBpE9rhZwwO0ghEX5LU407aPT5qPNjtMGFbB9YyhpoWPB4nckjUpgI
BRk874DrliY4tzpEHw/X0M596leGw8QgxPzBShBmcYa9q9cHDBEd7qSEhcIiBDf5
8AX5qZ9zdPfCbSvJCUxtRr3NZ4OgHhumlTHYLgDJ4xFc0M8BpYVCcKRkl1S8hlTN
sPh8j7y7NAeP26RFkXVaPkB0BXolNTAze352XbvRd7CbPEnC8QWj3+efnIxc1oBW
YqO6go+79tBCDEHytYBGNU9Vd7CTodWScHk0ep++/yNB0hT8c/65fEUz4mtDfqTO
FHJRaXHSWwT9YmYo0PH9jS3SPQPoFmvBQtVByL8uNeQjVu+BiiqNXIYqT4IQdwsn
YWzOVBCGBPxRLyiA8xkH5cLR6Dn7vgiw0WzbpXWCSMLemIaOUY/3Xnh+esbqpJfM
RsZiF1rBFGxWg5N6AU+cg4TJ+mPjn39ooCxeL5QLZy7r5+5kxRidFv8vH+syDAzZ
Wgw9KxjdjccRiRYWcqjVyj3HhWzH2TNjcvgeY1EtkXToZHr351YQTxRHaOcF6ozN
HA3P/e8dUbuKqA13H9xHs/VrOf9sULXp24R0GnjkXJ4eOAFh4VhRNi+KpXpqmPu0
UQDn8U/Ukiy+XrhpUiGdPyECly+gDOYktCzotSNPUyieVnERhKvNVu3dotqdqS98
9QLjp+P1wSh2ly46PQR/t7Cc6QGMOybbgXww5Bj07axUQLNHov0MlW9h/25WDFdy
YdKCcYo5pOxY5ahBOYygBSCxUl83HW4UgOrXHYlH8ADNCsUa2bJvCshPrWrmbbjE
jmvMoL9BrH702SjKLkQ6apFsxifVoEqGaUqp6pRnqBvSWJ0WG676cAhghg36FXec
Y1bXUbecfERSq3g9rQ/e4B5iMuYBX4SriaL1EFZ68pNIA335ZK4k/j/KMapQKSKk
zlqC82YQ5EZieNF8wIvohsxq63teBNVYX+Sm6QFWPRhVSlmNjKRinLzXnzx8j8ux
nVBjvswuw9f+qg4hFHA1TBQlUUhtyNwD8XyKlUi33DtagX2LMrWMHyoez4DX7G8L
SMYf2n1qetJlJD0POOAaUpknVtWwQshoiVjBCOhpGWioeQ06LmX3gumQ6pVeZlal
HDLbVG2UtxWJ568COe4lL/2IJorYx+KlcSmNNrlKZsfuq55jHEMVG5RaRiUiTmra
J66AsWz1YNapLRG85nqQdjkFDIG9dKAC3FLO9H83boVgXC6JwXish30QBEYbiUWD
C5MxVS81b93kuj6yYl2ckgvgNQuFYJwX08u6QGR7oujGJ3qnNtB4qi++ZKvpAwsD
U7QNS153006C/mes1G0H1Rl1vxJUlbdOkBcT7J7ZDNafzhIXa3CjfdBCDM9ynO/8
GyT+iZIBLPiWy+TSgsTQmeyUz/wXyRx8uVSo+PUbH9RHAcC292pemmB/Hf2JsOk7
hk+hGHWQe7+2rgnfJT2GFbzDl5DVU/v88QjrnkOOkHlVByubQUy2z4/TtWOsArBm
zvG/PHM17JAcscw8Fn+loJMqYpA5PQru9aTp7qz8YKjeVYfn/jYyaVOUXAOsLM+S
MZ7bYq03OvthUFdTVEHsh5r4L/YqTDIL0ECD8izp3igfcFroWwD3eTDQzdPjH4vy
QNztLzZqYoeq9uRok48pivUalpvyRQT7oAOBT7DbWWcZ81k4THK+AdJpdiUzqwff
NVCwjY1wDkJ+Gw6siCSD+j13B1MAzdRddey0wGvjzs5hJ3T536S44dpPdmCKmalQ
EKo7kMLiKskHHrcCD0tn1iZkP9RY3yLijGUUiPIIVqEOOIFtbylg81gIIsJ7Y82D
sm/csH/3gOgfIiGMW6kXf8ZOsTkv0pw7evRwuXtM5rnyH0+qQkuyMmee8IZqZyGW
wJtzJFVxW3qz4Fpcvf4Qh5gwjK52cf3QLPq81JsD/IHeFOW+AHJbfqQN83IhZMFJ
Ac1YbKlY/IIFqGkCa/3HofaDwUAHyhc//hvkLwgeTmIV9gDq9ZBHmbX6Iueb02XF
3Sfqv6OkcQ1tAR8u+YealTUlGBSYfPtYjhRHHFzojngdRo/33WIlxFza0ySNP5UP
I+Ci4o7olzOdiEMglSLGLyMOzowTOR456Hlpq2hZltJmckDqwa2UuH5e4YEPyC5R
dVy1w7qGmmaNht0b0H6VKoh5iZzlqv4I0GUJ8mY/PUKynQPJ4UDk5wt5H/Cgt+cx
Ku09oe0qtJsY//c/jK2w2s/QOuSYlhEDG0vMzvm3fKQmy5nhBaTX4r4uJGtzbKlx
/b1k6pt2WvoWqzCLAGFlxl7JrcORAUrM9dp+HH3ZG8S0kj2F7S0e3zzJjOfSHQqE
nH5FmRhU/zW3WYGSz/NqKb6HkuK52PVgFaXMkg4pNmNeIQVP9pgV6C8V76JrFT5+
XK2WB5D0iJnA1/Oe3s33jQbWvODtQFFzUqk4Jx25YXC6Q9XMZ7Nm/TlVVpeFv5vj
v/NIBhAcbj+hqQJu6l/hGUy3sb3syD3EeHIECLz4s/DgS/n8MR87JoNwRSpdBb7S
3h6pB1qj3NEiad9cLkvoJOWw2IUFStp1FqLP1UWMTTcolIRt9r/pa/TjpQ6CbaGc
A9TOVY+OmJXE0uemKMJQ8DHhbOsP5fvJ4FJn9Ff7K/aysC+t1OZgdJ86K/qVtetH
pN6aBYa9DNPidIvD8+1/HgeKTjODZqQUU9HpdvyiZVAeFCYAWAJWJRyTZOQYrfyW
nHeGwONnBzLSpOW1LlE0j2tSU0uUceEo3IUbbVG/I6JniICQd4wY3Rs/TvtcpA1k
1isASXo7mFoBdX149O4os0bwQ7mw24UChYDMciFF/Atkv4WR2NxlTT5rBCWBXcwE
uDQrD5vweOJOjUnoxYMR9csyJzH7Ul83JCyGIOBeJheADat589DEU9VTLoaQKyKt
dHuPEhDcWGU74a/itGoOhhh/+mvHas50SiUvSMGpQtXWdVHv+HyhogjDT9x0BWWk
LbvTZH1ANa4IOCNi0/E+Jb5UH7sCZjUfdQ5QNnW77gdQeoyB/G0jslLYdaaJoUkq
Jh+gJtlW6E/kkatGdCZ0npgPVBiI9DujIDj+aQyX2C26ui/crHCapMsrhtetsEQA
x1qW4BH3q+rUnc91i1joI9Xp6YVpDLeTYfqUVOkVYhQOsvswdmZ6IurHo6OSVAJm
YwkqUJABn5n+YYfIPdkCfvjbcbSXPp9Yq73JUXvbR/rSzTbKVUw/szQCIaRl2k/t
D46I8IOsa2jl2DF1xx3Uv80VbwoJrpqQDf/oqfwf7lj+TF8cKIxIizpjYEag9swm
JD7MqgKSxxAGzyH9/u454JlEUzW9mxgk0G/MeiWzYCnOT6sbIpinxb8f/1SHtz8F
6LOSufsGPXT1UkdODxONEHFai/+VAv6v+xtGfi+VlZQOGzOE/mNakaoz2RC15h6u
WTFFzt0LxVPCpuyNZmH29PEPu4R8/hMCdnNNUdo3mAdtVDnbSGVD0Qqek37MP4T8
Z4qtCu2CRwbrXpl+GkviEmp6vdT9qUa0kFJ8xUf54E9eBjzcL6U+VP23ooNegwpC
iPIg+Xkq7GAh25RB2Yf83W2yJuKFYEHV01da+aHT01/+j3nVERVE9j6/voig/F12
MSn7/0jTPemuxG9Fd8d+fBrt8P6MC1pvpBYQL/sq9mCN1g+zZUSOU0Hql3nJami9
Ezq6CwI6i5KxHApotpSya9i5f6FM2u/8VzULHsDwjMNsnyad0rkBAW1z7iAnfn0V
e0Wrr1GEgzLrmCoQya8dCFCryV8pSmAP2dwLe6fu109PVo8pvg+bm8H4LOxA4+TQ
H0LEpwJ6TYR3U9IW6jLmDjHsEIyF1X42SbpVdjD4uvKkB3eWQKwmb4nIt3lWm2/c
StxwLIw2+WoI+tvDEe6gQokFDSRZEHJeTeY0mIWSd9vwpfyz4eQ3cVuI9saRte9e
0a7BjrgpyL8/Wgz84UTq1r3VNooPu8glfqkDTU7kGInak2QIL0xT1wNkEJsbV0U1
GZEXyKwrnTd5mKrVok7mR19NOkuCoGYnX0/PzxkjpMEDE80QmwXNrw7yFHUi/lQC
gEHmyzhYnA02u/wMNE5Xl8g/YHCLS/R84HF/5WbjN3bZDTN3G8tFyPkLZ0/mIWtv
OLJZt1bATxx4rfywJXcrUnJCDmT3vZGAha0qbDdYm8IaH3SxlHEr+ZdUXqujEffy
ivyoDIQJWpZWnXuP1bLmbyDzCx1BBjGS3J/r1AMYSgBgulqnIcusceyjU/dc1lBP
4XD2HOH2OvpDSApSCPbGmPep7nPm356BRzsT/iPaeklelA5S1Y1Yy8tA2MQ+VUMg
+8FXZPSijRYFDtKo+5uxc9NsySX4dySkdFzDsiqfQX+/8mjRTKCUx/8gJQOd87I3
idWVE017FIEbQih5HHD0UHXL/ofggZYltiIaYST6Jka57NWE3V4iUoyDbwA8V5mm
JjXmoIAU+1coaKvz4daczT7fk1M/RmWnTS79IEy9bGGoLUHxVXwtdAQa7lIsmOdy
Afx/oCem33p9cGgIhud4w77InYIsNJYKJx/1+u2eqi7Bt7UJ5dIEFb+eH7kJZbRH
LlmkVJwqR7phHq8Nf/B+wYcZwDltHCSOAA/YulrYviXdfiUjr9vEhdS9axrRJ/l5
PjjFk2PmK9CNYvdff04llcfcnFria1/qYgVyh8gm+LaWwG3Vo3YBJFWbbFfthEoO
o5kxKg0Jr1EhGzFq1105W8zSHw6tViEd8AsAUDqADggyJJtg5oB5oxC7sVQWNr4z
F1/DpEpuGm2zwYa+ZyauoGUKOwwZCxgU7Gm0gDLkoKbSClC5obMXSCdeJ250ldjS
gSYZ3Os54m9o6rUjWayBSI7s7ePNdKLPYRfkt3FkceJQQoUrXjEL9Y0zAfwsPAxL
0qQ/LEnObivSgLvxx3C5HutWufqIYecMb/B3AXavE3sVwytNYnG0fS1nC4VF7s20
r610+rMh2j7eVZu6jq6WRBCY6eZyzb79OWJtO2JcE9NHeZrYQ+IetpwgWe+0Y1zz
mbNlHVsF0RvwsXtuI6r6MOE+Az6LnE0RdZOURdxSa5z0wKXcdbhSmemonPV19Rws
zppIMlD2+PCkzw0iZBo3cu4nbeeQDtnCUPTTEAojJceNW3Vl7XBSALdryGx+3b9I
td55epZS5WjrgppgMHtI2NJciRBeZClxI+Cm+hWKO4aDaXkPOLxwF5vRH85/u/HA
+9HHSU4xvtfGMyRcL4ntV69gsjhzjE7mVHWe22zhrKqgq97ScIrOYJguJP+8YNNG
ek9ba5Ym4NPZ7uDMCjAVWaoBjsPNpT+lw4d0b+b5tZtdOa9diJlAkbgw3tMc1MZt
cuiDIT2VDxKPS2pq9VIdpxZtgxQfsiP/6dXiMIBHMcIiJ79YHD/MAjmJ0T6nY5/7
XqMFdTGS7dQiXKyAKONVwaRDnw9VTNmd00LdpJpqd20XKSDs4eUD9apaPSXdz/fq
vrThTNSQZQf8qKmBWAqDerpE60mQP6ePLnz5mSscsZwaiqfGFYZgQyQwtU3T9Gb0
D/reJ4A4LllqCWZS8y8Gmnq8f0luJCT4xn2yM1xi5FQQTSzwr9TAoE2ugUzsMSNi
Rvd5QndQ/7k7nK2cCnqKU9o8XJAGsDZlSZ9B0fNcLB+/IVMzy0G0vTVAjndBa0dC
pNPOFWOhKtpcfUruJlNke61KNxCkCfI+ikNd2ieFt2aPugfVy1IxiiWheS+/eYCU
+uNyt2xZcVeCkCx1d5zKuO4HFYA/KkyoQseF65hkS5qlso1UoVPqK3jQIQ7JAFwA
dIQYBY+rGq5NEd9uyqJq5LP72QQb5LJVIFIx5C5JHC2CUOmSMOGKNV5Z6dq1DaBe
DKGM2tWpwfGQ6Qy90f9NNrCZ34NleWYZ03PpxhCSTw0Jq9+zgVH5vVaWsaXRSv6c
8oBiaWaBqbRdsJwJqxupFRpc469zi1gv+JrLItZa2V8dDbdDdTf3A1D0vDK/Udfr
NLFYQy7OcNpsCcHq4BJsKPNO9ZuprLkS1YMRNjlB0Dzie5ouf1qcN+KjaH1btRTS
QqBtUJ8ydQpJjk+uy9oi50C+6ldX8kckb9bD8ToT9wHbR7mkFpr80PKhdpd+x9Z5
BqlAA4hK3j/O3FTVdt7swyzCP2Evv/OXM96AjxmlW7zOLrm04TIi9RMNtIAJ/r1S
Wa1TsMDURCm0xx0VGy0llS8yo9JSoSkKddcft5HxTHMUyZwHrKID3iGAuTALA0+X
7E6JeEFpuYmpzttqAGHJ4dlljUxa8TOCRYg6Igls1jNW4fGyloXEeI+B+Yo+Upi8
2ApUzCPK3cBsuXLZxiCrl+8UskNDFtlLZwfki1aHaSaJlWw/lpXrrl+LOexnJ+ST
fWAwsrFBTCuyUmjxa7aTgLBCsvvuPqYTx2emRIOpe1nXWbrsEq7FG9YFjeZUCQEj
LpdEwHDOywTCYpmBOHNbw+jKaYxMmWLdpIkO0bO2vcf1mma3Rh1UlQO9/cyGGuHQ
vtdBD6SWVptKJfL2IJtMdP7hVPfMjety7crectGI0Bg7kUcjOuytkW7KRFOePxpf
+3r9QbGX56eAlk7e5TR2h0XNt4IQkwinMQr/eKfibNFZR4jV2xgPWfO5s9FHG2OJ
UUZRne+ZzKPOMVhzb425RxdYZzQ/lVdoKFISaKSQgKsQH3oC97Do1GRAWi2/Inai
mYg261cwiFjNMYfTXs0j9h3sEkOdXK33zj4Yx0Cje+GUzSAmYjnVzL6amu+PAm31
coBJHWvf4yCBR53bYaCuoHL29zSLqj/e+EhbsTcYMqrqFGt+SkB8zy/SPVBDGf4Q
xMYowS8KFOqXW0/ZYIeBzMRQMm0rD8WggeuyXOyaiztrU858u3VcLr0DIH/GpitY
WNvEWRpESQPYGfqjLnZSzSJqqecIhJ85yaL4I8z8fZjqXsKc2kzSsZJYdkGKJCjT
xgrRfAaQkzdkDnSVaYwmXKOBk2q14OiE9WNOYnV91d2NLfaVgJXud3UM1ZiJ7Bfo
+jS9Tt0RNmcd/racjqdnLIH7/bHt2lqFzua0YgxfgzU/M9e+jiqotFgTwCvhf6Fe
NKY5zAJWY47/fN4yI02jt83y+qKw8QRyHAfffKXqS0lWuaubEj2B36ZpZV/Zt8my
ksDdDarWiPn3XRzGhLlsSVvfROh6Uopp3UMUvOO686ZjA+eCapY4FqiSoxNQLQm8
cB6ua6yCxwWal2C07nkzxDrQPa4Fdym3gLWD48A5w65d9s2kFHWZE5GdEQEBhS1F
ASa7aQIweZBPI08MuYMDyx+7vd1SViTkVhtRGbL+s+yjXa6M8fWrmRQGvvHmsLBQ
Bn4rRpwINVLEmy0lcCaKKIlQsn3RR4IbK5pUwGo5Q5wPN1H1X4YPJOUt2pZ61Phb
rwJ+TveC6fGjv1CDKzQN2Vku4AOC1J5/lziPdHIhokIQmNz6tXmTLlt5it9IFX3M
vHBI4D9kpXmhyZTwGbnpzCICyr8kFbjwR+hTKWkMfbxUr7U0fRRDh3p8vFgsFpbO
7sO1D0EFo+aeu2O7t4cTm8vI5WEsc/8jPWlqGfUvDzSmZ9GxYvRIFiX4ryV2UmyU
SrC12yBd7nG5zdAeodJnw7raF9TEdklfynNTZ1mJT49UWOIbs6HUnOKpUGBju+cT
jSnBIL1jWAG7sEE35rsmmcVs/onIPWds0HTg3uL8z4/SthctWIL8AtYae7B33HT6
AfqyaG/vMGYvRyACsBfCzHMj4BDjWy7g0B22agy/XkN8VVJfbh0dWtOvYZ82tMh6
8dfAY7zlksqDduu9+KmUdQ12DapAPByGE99kdeAXgrU2d8wJiL7bYb1Hu0jjg2Q8
Jq85xHlvqZelO7kedv7/Yi0fJnR2zBmabSnGsKJ100mXZJwpTMbAp6UVVM700dUt
kjlLKEgRpL5hIwNCDBzcHwrhK5N0IuCYAAvIhWH+eAGS9aatN3ExAHTZwBZWV6L2
bTQgj5uXws/GSWYJdNd4hOrEyp4WnWnnc6VKsiDMZKKoHBjC093Qg8RYMU65F5f/
FPIX2M8WjnwnC+ENIoEs+0MfOrE5OsCqyIbY4nJzqMb1AMPBVQAi5S+qWCZ5qC36
oDyLvHQ7dt7JJ8YB6j70AaV5t4b1hlGYK37G9bOpoC83pCk/TKj3j6udKfoMkcNG
6w7vPWnZ/DF5waSo1rXzrY9Va78ZcS4lBJ99kMpovOWXuT1xFRQyGs2Y1NAMUW64
aQ3g1nQdsIx7A9xgm5jMLNUv0xRknabWeAvnrdmSZyc4Guka9NJ/jxkPHEC9cOuL
L0tSiNXiGDxxfPYjc1PszzyDxDdg6bD0EJR6GTVZs6hiiU4Cfn3sFZcKrMCjcWpC
LfjG3U+EFCTPuZAMVLkYg7OdOy52J2CWb5WYLzGpL0BtMWlfQKQyjrFQEhyqTXRo
Dd7zdw4FrTZeSDttSwo3fj1dufA590SsgcLuqyH+HgBmf4IvvZEUuitc3I4m4wOI
xEdVW5PMBMq3eHZZwN/eKyzfpvAmxvA6BFaa1KjszAQ2C3dpLzmGQ7sO0NexkbtQ
y+l5gVoNt32273I+m8xg8RwTkdsg9CD9JmV54u4oc671FnTQ573b+5gzIoxQYmqa
ap7no+7X5zv6o35+NkMnJvJrsXm9pXTPRoEhKlswfZ2LvvQBFCIXJ3QDVDs9Y6ll
EUSKwUf/mzKaT75K0zCbpc9MIp/Kl+7Pxm/8ey/gU2gSQlmbe1PORgvq4nW0r2qT
bNl32hPNKb1yOV8MusF862PsT0H6ZlGj2eTG5RxB2nMpH/Ryc4nOqP9yNZCtNIu9
jQLJv5rAbq5TqD4jlr1oO93gN2D/fv/llGvWgm0KDUmxXAyFPgg60kvQZoRTLeAW
2fae9ewJDFUWl61qwHt46re7zUkVqwXfJBjuuCfcHvDxa9kVSS78l2aYaYZubtym
j8whEaWan0LUtmK5GkyF9czJqQDi20OogGV9Y7QaZZ5B3XnQ8N8DGpm3kEoY0kfR
PujozWv4n8WcQUj70N6YBQv9rScX68hJKnTbPrPWQan9PgZchVDT28dL+YqxZE/b
WkqSO44MYgi3gRiHZsQCufBpMjR6jecWQM6QUzIRR6tFCslm59wRYoNn4JJ6/yl0
dziyGGm+gO88+C7K1A4iXqxYoO7DonPx+aTdCYNrMRGJC8ntpt5MTwZ3i9mFsrpt
uSdeHaTDPQlxjKeCZN+Q3u1j2hx26/3oBYCXFPdrmoLhWB8xZtkmoRr8B40gglmF
MnKToAxtsCcbMtGFgssFM4v6VueqPR4cSwm7mf5jPSYuEUS5iAY74DWbHYCG2Jy3
5xpVR6Itiir2+Hu/mEqIIqpHWMAe9zF7pSJlEwbdRxS2iu2dXYFH2C7Iomp98PVX
JNd3rYcUAA9kwPH5ZWQNlvUd5//yWw42DuvvJ4yvsG0tBtoKvat/cSb6/qh8OiYC
kV+D84JEBupYilTb1ypoJsUtwDw+aIsR+LySYmeVNiCSmgccoDn4JcVf8FdyoNKM
wWVVEqhruEf9lp6TipZ7zDD2lhclQQcoWePSV1H2nM5BykndIyYHoW9MnvhHI7PI
Cb7nM83Sc9eqJ/BfYrlOZV9+Lsur1UjHPB7yYslTG+tYWDBg8SGOJTanIrR9QMpu
T8cy1GTCqR4s5D8Vltw5u7El1hZtDXwexmuewSiBtdth33cJCAEOCevgsLwuSWx+
Owrmvy3NHMZzrWPM5vTXSWcDInfHxo1yyXP44Je+ppvAY6SsRGFjT1JBYhtGyofC
0sNowXOab6jdtKZ3QqwBPTU0UWGQhbcR2F+O6VyHaTKNiYJbB6CZP2mZfzFESRCp
XEcWNy5iLKkECXmqb26tU+KP/M4KEaivMpeGDxNQh36Yv4YibcuaNYJuez40o2jS
RurRynuhuZA0gnnZI4ZL8VKz8Zg3Dhn2U23bNJQpq10DwjPID7YZy3R+Z8v4ZohM
JvLcJWOqdcqVdKvi4/0KggA0bRnYtWW2rD1wR339XwSs5QUubDLV1HL8a84nad+K
V1QFyyqK3K6m/8uWlNqYWYPepHKck+To2y3TN+1qH+4RLPx3dqTeH9yBP683E5DC
OcEotVO4oIR5iJtRHBuotuo0By6BJnScOqja3s/9Pjw9x0QiqxyU0+YDwczUMrA0
J0YsZa1B4+9GKyni7RgPVtlz3rskNxplARTKtVLlNj8Jj3vg7PNqEMA0xqPU/MZc
W+4G867ckJsoZ2CE0gDxLd9fjkxDzwRBlGEQVnlfL2YIpc62yPoghvK0v1WOwaUA
qvd5IuU40Dlu4mRGS/WtU7qSEQO+uGQHWW8wGq/QCCV7z80hkwS/WCaolDyp0biQ
siunxi9GXgkyQTNyV6FnaKPS+y7GB6EhyEvzTr1+k4pGpX5JdAhdQaEzr7W2EEk4
EyhYK5L3XHmvQTkCzwXTh8rbw5xQM0iAubKvspDydV8zMGQ4x6lkV8511aW6nMxH
zoMBkotCkEclWZXP4AvkT9bWx7a48d34BogTovwYxskNnZ25GJwzqB8e5gKTCaRp
KjXosKmlTjRUc6feD8rujvCgNmgWCghOtQbQCP+GUvCBaVIUoL0WM+9h/Nb7FJO/
mHzmuu88bPxziLm7ubngCjJoOGz3VjoQtHiVtiy4NF/0Re/LwFo25wmprGhsbJXR
qoHT+jIP/Jw/3141BtX5zrOg+PsY8oFz4fS1o3ouhiF4W3uXNe4WPzW1VMQaQjJB
XThRwICkoFU0SpjfsAp8CHwAo+LLKb1V3hY4+lkZ0GqibjrrApjO+SaZJuhrMkEm
k1mrUn0NdtJV/6h5RSachAX99eOd3raygJ8V4AM4OgljajbV6fyeE1kq/8fre9yh
/NbH/zUSormeRzBwee8StigtzGCTfNoDCBtgOw09ZaxNr9Pf2PnHoFQbYNpd7v6p
D3EGuXMB6fFymm8/d4yCSq1u0gEuNwMQzBEQ+1BuwG/XA6wZDR4olctnGPMrcFgz
6FWBKWiB8exszemyrv510mFQ6MjZ2vkzGlM7jtxNxoYjFcG2FCkmWSl89TzM5xOm
44iXqX51k4JZwdH8T1nVSwp9PaRwBUxBd6qO2GefDlC4LsFNQp4WhzEcx33rXpBC
DfD/nPECoe5SbRXIR3Axzd4UjQFBy+a3DVkboUxZLe1H9wvhGCu+DRO+rEU8jQlG
iq7icBbteb7y5Lb3R43M7/ZqrZsWYa5Cyip77Xv+RG0z2CsirpFNvJK3BXMbAe6u
e9goV9oTurmm8MONRMY0TQkVEwdb6K4FBPCi4x4gl/4apcaTifN8T5eKDaGLXy9k
aJOQ2bjhZrhYXd9JkpFR/I3uXfKJIC/y4MmgH+Ejkguzd0CIXLBFhn/wfoTvwPJA
+mEnvgURVhapvLqOCmS5k6ol5seeN4ceBNH7InpfoLE31rZ1tftxj8/AinGJj+CA
+5jcnMHZDh1eMX4i7weWF5/YVFFr+kOEv3ahnscv8HCh8FLdBnY8y2X0bfSGNPC9
jpXSjuoKYkZaqrEwrOIvsutBWvdXvzaZDYsqMKvWPsZwx4nuDySQyQGiA15S7lG4
TUEAjDNpBHeJEM6B1x2wyfjmfqf5w6azpgl0UDC+NriYcSRMbpm6Ah5dOEQDSVR3
2utY40wMa1AcIlOqi8YB+xXo+KGMWVpZN4lGMFjIbcGhkcsvB2HymnvcFxwizeNd
mavp8UVLhpLCYmgsTPPJ6zj7lPhWe5Z+VoslKyoDaC1dLOdKO1QmTpcq+VXSM7RX
jVgeSNSrcxDXUGFmJDg+fIWuTMn2vtI9PE2h4oD92wvsZRzLLOrXVIuq8oU3lme9
BIpLXgKhRkTdo7sMpHQBtiGwF5GYasE7srlO2dlscB6URPyCkzOQz6aL8ZP5oY2c
V8yxAr4p4LbHvBsUGLZXSGEXRigdbd6GQ+uZixcOr1h7mINR+GjGgSpnqMkQXmzc
/YUQWyj+QNg2x+DbQNe1LO3qvRfNYBK17PC4i2dozyXYWFwmhjylE66MSKbZ5rm1
KQ1S3J7C2C32kbngGp51J7Z98YDFEa5RulKXgwT607JZBWLbBvcPWnvJk8/qr00t
4J89b2e8/fKMAKCpcVZvG40msuaIeUlFty0OmDudoJd0ASIN7yWo3ZXX7KbzB2Uq
2D5kqbtjmbybUozN2LbDQMJt+pSDRJ0NcupzCklodykwwHaMtygN2OzR2rDBtmMv
Fiqsv1/LIQS3kSLtTdOg/IcMaeEoVY/Vlia/wiorpP887eQIhTp5w9V/RSP4TyvG
uu8jEBD5VrCmxlhU53y2xodKA0g5YRVLuzKo8KQlXN2p08vP19anLYN8L5fK0L+j
C4j0+b2mArlW87/+r9jYuSEVzilQeSgFSO4DQ06kClmgkNL19QS7Wg81vc10aOlq
xJAbObB3y+7ofFzarBSkgJ+Np49OeaHHOWxSpKNd9Yk+nB4J5pMA+txjB9hZDfcH
kvuLENrc03JH2SU/JtJ5fBcB6MtBhi0MoxUv61gduv5+nWVtMBZ+dStOMxO4v6Lg
A/3I/tLkzu9zUHTsTE22NShxqKCLmVfbcU+YhcFR7Kj4nNPCdiyQ3M+CKRDLK4hL
HyTbw2eB1py0Lc4B5BiozDtEYDXte5o7tlqnJ0FSWL+yuZ4QjwmImDd7HsFCGCST
R/8PFbMwUeJCSSQvl0cHXBK1ozulFw6jKQ7AuGRSvBiJUDs3fSbLXfcx6ka4ouKu
LZqLa4U02WJTtAxSd1ySwVJBswDcVLR8wrsZg9J+66PmvlA8TO8YEnOhSZxruHGW
vUgtuVK/GefWLg0CrIzpE69OzjruvsrSGuOoARwuc1tVSrYqDmCn/YGaVjQQfxAs
DTVvISIVI/47yOW+iWJy/6wPhIyA6THK/JB34CT7wwe5JkjHB16f00wOdnYGhXCB
a1f/EtvhlB78Ol+ZISJdYeLcMwz6YXvvtLblUE94crahQeaSCh4raWRL+X9Ytb7+
7dO/5WxqjCunLs7BlFgRneBX6yjUwPGEbh23x5mMZeDMelQWg+wuNCfA+dbFx3fj
7Fvu+5E7AZLsTxu7zIkwLOlJeZruGpgBv+mtljrN5S84E20i5VAo4xq9xGVfIX2q
bT/D5Nq1JTEUllspNENDRvsI/IekT9gtMXhcQ0afgVDnhA/vXzZKdVRAIqqu+gDO
sJU617eA21A8RrukGvxdFEtm0cm7IUJIao+hsq8Zw7XQYxKgKJzTJ8UInBJmA1S0
eOvM4SIdeewxV3k1RiRQFb5UZY2ecIE/vImpMZrlCZnTX8Ugy3i8lhIvRV/6/GUj
vnlrzQgTl7DAOHh/Efs1r6DrSS7dWaPGXagjR0poRTa7QQv2gIFCHbE7tiy2fGmb
F6IuznanHrfbYndqmUi8ur19mTK/qt8ZpTW2cs43EXaB01qTdpL6qCrw0Ba7ALRp
jqyyHNRZWng/YfyQ3TOvPg2ld0RUP9yI/ZYYZJrXZzmoKX7i1390LnxmQ6geLC7k
mMv3HclPN+CzTSlcxCy6e3M03JxOdrVlPco5c0VkMzHdrtau61d0K4YIeaHbd4g8
XPInnlChf5OGKY1Qfu3CrlVQ8Fwdl7xerTBawpxn73rNrkSTS7JpW8NJD12tUtso
YOU0B0zhnHrFT2OrSJ09QYtB5HhR99kdEuSFZo5MyZ62lis6h/+76PcLtkmlGLFN
b24IXQ87LGeMP5x1Sd/I0wE1mSQMdUF36+zQJkFF/ZHuXY3If5Jo/j0VCx3Q5lN4
tp/ZvAWB9ew171FnV55VpKx9Np6oTcXPf5dxSCL6cJNKcnnnJxP1QeSYxwi2KFog
Hf9IbaVWrtYIlPiErDe8wHVqe0MrJDkIw6riGNgtvJlgnYBgRuLKnHZyD/Kfxils
Dzq0liEVxnUZzyteflwG+FsSvZ8M5EhRCKhHN2pWp6+0UjknOZEcYIXDwabn/81G
mz+JFJvKTqf70AWHh7ERXFq88PaOIdK1J8orkFergvNpI2XuWRGtNjvcdTwHy6OC
045lXtMAyELYd3SMqdbx9o1E/VfjXn9jrAiteLKk2ukvIqIUEHN2AsM5WQ2RIVKH
IzTkV0uhK+eFomonO9QFLpbzw6oY2A3b5uzEGgPG6xohGfrH0SWf9apkzJdnT6FV
XgzNRr9icbXVLzVklH4itRYAHcngQ5SaPAMmIcXdJHNZelD2EJta2FCFuEJUJfMx
2yJwPno5pExyCCMPOY2FKCd8nOtCk0/iNf9VKkuatvi6W8wyQUm7DDysDfg8otfj
dmUBX9C2p72qmN0sTjg3FT0O+kq5UHFPxWbmrA82ui/ca/2GnQj0yz8ArETxL7Xl
3ou5F1/YUR0NDXGrEKrzsadiZo/eMQ7o9Nda9H7UQJdzfN/lSWYJZLbaCZjjs5A7
dVEy05plV0c3gXVoPqoxDX75yAaJgadZsBaE7iJiBWWJv4E4aFL3StmuO3lqPc0/
AYpaDVzeIswQJcq2dYGl/KU/5E8Lcoe3hkBwsTsn+kr92eGtdiD9f5ha0njAFgOH
nqRIHasf+Q1sqZniaIpcMX7nYL72fzeqcB7ikJteHWQ/a/O2S7SJVPTtKTJ2UqR0
UauOPyfJLGMnYt51VPiyR3dZCrHri7NfD9zlo9gcqw+MVD9Q9y2tS9BrcNI9727c
EKl18cZ0vYqD0zwKv5lkEjlC9YOnOEdO3zM4sAfbE6zephWtzDyLf+yFbrYXtzv3
ituSusnRfHHJ6EV/OPQsx9rf867opFibZaT4RvISBcCPfyIf+1H3qEzhoP1PJroE
0v9HGNMivDzF1yI5EVHfQH7alSTaIIjXuI7R5RRaXo08M3qBGkBmXhWsE5X6X5FJ
+3cMj7jLunHxJBGswzhYapvEekqmEuGYbEnUkx5Jfpq9sb0uEdGTc0jx4U691Xyp
x+zokP8dEzjuU1lyaLRjn4oFYeY4i0XuNZt4M17NngsUeuKR9oTNqY9saTVrfDJg
S8fbhVIVghop91jXQudYyX3MafPIquZyHUhyvTQ5uQG43lGDt+XOd28e0z3Ic7ji
j0snWJkbdcRjLQJKLYWbqIIe+EFegZU7rTn/3W2hE+84j9ntCGFsTlVfnBSqU9To
z0Hv6Ki5adkbbz8+r2Pmq5EJ0k02KEtQvyG+J2F6QxgLzxWYjY32QlgGceZ/6+/5
3bz3V/o2iAQ9AGp7TADTfwVnTXA+Awf6dpzg3qVqj4zE7ZJrSp8ubOvYHePkf1so
yt3VsOn/MsFuiudUabWGF0JeY/XBEW6041NSpjBFc62yGqlgS30mHq2u4QBw8/PB
cyFqJTwJqznC8lcK61Iz0imnmF4Drgw02FRMz5TcEMzcNQCH+tmE1c4RKNQ5MXmW
YrjyAl6vrL+0PHVEUpXC3XFyAeOV5JS1OhfgUpnbotFIQpxVDf152Ow6eSVJ6Fv7
33XBa5/HEbhWu25x+oEHANGRu5DpXQJALbC4EkwTzKoNbTFiDZYxi5h1AJcwnRpI
ZWfrGAFqJIl9vzkX8jZ5cTlDDBJYHMm2aQIdF38LgpN915Tyx9qGDmKcxvZMMmWI
i+UJkOHXt1jLFVuLXAz8K2GreQjJDCeIO3mCJ9KmE7CLwLqcqZ85tQ7tLS+H2+LH
qO4uck6NVS99ML+OQUiecdavt3jymfgNRBq4THggW1y6nEWe7kz/orNnBP4vrWOo
D1qC4pGHxQfHmyK4cstPUevncYiOTYFuQM8PedGyZpY1Oly+mUMSSjlQppdP1Ezb
J9DR7Bun0H2QTO6cL+QPckuRQb0bnYnrzF9geXm6EJKsHfIiq+YcTG5KT230IURY
byuAEMcroP6L0WWPADq1kg+k6BFRcD//jkjmF4C+/0jOGpEl29MRmLYC9bsHzseO
5vV32zK98KDKmwgNU6pukYWf1J2s73VFbmDniQlL/VKMFaxPAtpKuqKLjrpxsIKF
SpJmlzegaS3+D3TtekxaUEHiKqQUDwEfwYL49+EOsHV9SMi3kE10SAmTg9efCMmE
ECAraOvM0i3hl4Egddz1XhtT+JSMj9+EdXZRUNL+9iJvpW6Lco8rR/jgJjexVJdH
nA/g4JkNvJy+gFL4kZXjq5W2C7y5LfKXHkxKKX46vL8DldWtbLDAmKr/FjQc1biC
oz6CZ3VWD5Qkgg3wMFFAMe65YK0YLDC2aHpEBWLoXzHvpXnaQZzGDJ9JrJoGEiN7
4QA///JZY7KsoSIUd+RV19KhsNZLktY0es/gpZixqF9SV0GCM/Bqoog+G9cqPoOx
25FJaxoMJlggqZXrgaN6wZbW+V5TyvqdxxkJ2bmH35gPTQ+RsuAMVKn7JcyxU1NL
9j7mRIqW57G0IS/HOaoisVvNDfAya1o8Xtx9y9BwwY9QTszUIyy5YQmb0yUDljgb
eXkJqT9Y4wdC/H8ZeNjIyLY4PAygz8U7h7EP4cVZ+m5z4t4qL5CdAMvB916OEqMD
4HPOZA5SaBvDqbnuHr1HsrjILsJzXqhgY/fU/rtJI8ZO2OKuvnyofWLqaS+5E01p
i7bqy3k3ykiRaiJ6kuKb1f3r/GnoBqqsuxufmTjlXiepREsKO88ohjE8nDhehYyp
4umbE5pWxa4gOKA4AoIrZS3HdCW0C1Zs242i3Vrw5rwtUDs0KBLYxePGHQBpKJ5V
J2ChQvTADTLwnA9KxdlLyLRSg6Er5vtG7E2DlLmvXZd/yGJeY8pD2jYPVB2332L2
VWv+kO/NS0ufM+oY4T+XNR5Jr3Oyjod/0DAXk8fPeNwD5KwS65jp/chLHYpgP8EU
LOD3X4UwpVFlhoWjhlZaZLyfRTXDdqVPylZSYZX83o0HcBSPOAFkbk3C18bSrc16
f8+B7G4vaodG+Fpsj8WTFQyTQ1o4l6NhUk6jzSr9kyBeoJtzXP3ztDE+H26x8/RW
Xm+pha/ZUmFslXuA1uAh/blY81TdbQWKDlAeciEnDrYcyvSsDiwO4scVHZfj0xaQ
wapcvqgF4WrK168fy6ctz4cX03IWUMTh/hgcfuThjTU4SV16axYo/aRSD8+nBvlw
AQWM4Tn0pUsOFTLH3/A7xTN2qtY9cHtGRbRkqbx610DYV/lTpl4XIxMB1VuxhnJ3
r0kAFDGkoEZJH42yiSDt5lyuPHKjQ2IQdi5RR+COaFL5UQdC8HKch/nBCZVB/6+m
Cjib20UQqkoAil5Pz9NTGOuXHqOeADkaXtRdCZ9uJ2hDT57CY29teo5ufJf9635c
rZUHZvO213jqf2PM7ek7w/miwigWV2smJ03La8A3vfEUn7iezoGEu6R8ZHcucruK
onOciIYpxczBBP/az1znjjojctvssg3fbLm+T1KWpp4bcusgYLVpUfFiHPXDfkDW
zsU3+afHJH6aLTe6ncDm4COpMnhZB/WoGU4R7ScbiEmqzAs8lrug2jqwj8shtSda
L2GX0/oZq9NlDlvW5C7T71gMfd8FDGZNNA0b3nVLjWE5chS/8tezqC/6D5ey3lOG
uRTpVnJ8KTrl29wfR1Jz8bjS9BKyl+bM6rp73O8lPanLu+bAodXsOy/Asjmw8wjt
adQEtMC5FQcktTJSPNYr38TcZppgS3Z1OkOgSQTNOljE9NJp7Kg+nnd7cFcYvMZq
mKIZxSHiiFwPFJuRtO1PeXMSIFnrXjQaUQuMZedvul4Z30v/PBB00ulGOQSxxPeS
uwug2F89fM28iUBrjzK7vDiQAkvUy1aaRSdg/S/jaEKeDaU9xeFKNZiOdr6H4re1
iQanlXjuNVIwmLuKqDrDbe5ry+mUgPaUkVBoqYk1NfsARZupmJSwX/zdz5VJY5kI
Dp6aWScJuj6PBoIzS51NdwM7xXF4aLwwAmG118EousgovWd0mEU6wU+URXMJlq/q
wHBui+EVij0AElT+1b6A6Nf4O9Zv36oKW7EZtb61AhuI2AuGxRErLVLDkKa6iD44
1N7uXCi0+RjHrY4JtvrwEE42v/ynWmKmyWi+AZPYfN+DOmxbX7IrpAtRjwtcLPLj
bROQJO7JM+FHB6EY7a8512SHaWDr7kWzMd3T1HIppx7z83adRRq1Y422BAAFfPiM
94P8oyYsmmI14G/SYKWnZAgDBY0KhufybpJkdRkSVKqoUnCeXUuuCJbsr0Ofl/Gi
WhocUE4FJDWe8vOOyRphk1P67lXigfWp5OGtM/UhKrKRcICDsbvvYnjoYmEtiqhe
si9+6QQelbf6s1Nqa0NMT9bnULT28JvG4QA4r6Hgf3X9XpfDPzteILRbRTT3vZXc
FMoGEdRI+ua8rKMJBUsWjNZbyrjONv3xf5sCcqDZo+ACxOFbiO2laoFS7keDeMKz
peLkXgReyCPqwadp/ASAojUgJZ2EqVAYnmtvdyns6R+orxeHEZ1KevGYtRIPhEsU
VoFbqzE79lFrE3HBikBq+CwBlx2CIwLNaV1QSKVhSBtjWQoXObPvsSk+mh7R/bYK
Kl1rUSmm+e0ozeU8kF1vfIyE7hzjIUUKsix9gtDDmte4B+Op9KerTlOdH1Wjv0C8
MnJXMoTuIVke4mK5BcRhVePRLGf2rfCGqIh/6WwKrzMOVZ9vS01zcJAaMBdF8njG
/WE1mcnlUhVGLQ/HN8m3zXU2W2UpLy90WabNu7SInwFt6tZy6BVQR4mN3ydOsO5+
u85j8BY/hbv6jDsg+lIvn6g8J/Nj5p4YpEEL+ApTUzfCI+PXWn/cjH1zGmNVWN9q
zr5VzHnTcxSfRD/ASRkTYkBzQmuEUsDNhDs8Dx+Q/eFE17ZnWrLA0ZSMOcQOVcMr
6QamIzl7nJBnIJ/S5meOtq6ID6ZieJDJkrwFFuHmDdJlwAo2ATeoH/Z2kN2T4y/n
jZTuNYZqfoeo018OPoTSYPIPRKSzNdKKgNfb+dj0zptWReKjJ4WlYQWjDVtelImt
ryce3j8UfJ4vhkkG1bnIpwH8/JBxOG6OWLDu6Lh94XDmzY8zKuiJskATqKOl+E7p
nph8FUKFEr0TP4hikXCoxjl1uzusntZ6RkuTICuR5ysRrS6/fp3/xRrMsB92LByt
aKrLQA+S8Arb2NxfZKMMuTV3/AQ+ldur5FgdFPnYAz19SU+NhsABDqX7w6RlbXaV
bT6ayyTHYl7BAh+pWfMuxT2OyyPYs6oB23cIbQ24MCNp+fngUWFKc59c+lsumA+l
ysYOdt1ZGPkSpds39TwgEAjlZuAZQEUS7ARP/VhBJkZ2f+j8zSn6cCY0MKulsK07
geoNUv+WXRUFn1HapVndzJqrJmaCLVLNyk+Px6vXOMWL7Q6DSbdOwN+2ncqsfsZZ
fKK7+Tc7vY8dip+UTDhv+DbroKr7j5dA9iW8FtlkIJyikpxImimWfBBL9k0mLbq6
8ECKggPf529eArV0EaOs5rJiJAnDNBJXxG/ghOE0RBTfD5Rs0dF7DTpmArRlzdFy
unw5gYXYRRtWtiHhrSqDWWGirNARNkXuQBLn3uEeO3Ja5voGu+wNYByNWvgCMpvu
Gd8hSLwK6/7RVyZloHQg0Zg1bqQyEubkdhhVTBncykX4ThxdWDzEnLyHZTExII+W
VRY3vdM2gMhPAmCj77Abcg+Ni3JUZFjM/jTBp5ip85fWFOvhtd7rbl9Wg8fzk/TJ
dOAR1/JhXGo4kh64o6+OjWc/k6+c2g60ALo/GNT678iUwl5fONrDCk2y4DBlK/je
1V744EOXemawy3g11tciRXUKcmUOeufkERgzcMFjDFMyBzJDAtoKllf1GZAf8CkQ
oDUVpcv2TEh+gGB2W0R0gOd0on50OYGWf1G2yvtL3gvudforfh+33lo0hyl8YRId
bDMvhSTtGtKpx22BFLFlvUhl2WvLDpq5uY/A0+ribFW0pZjrmEEN4ktA6P7VLbw+
Blt4U7b+0jv+2iLPMc79az2FK/fbs8k4CbhFBMveaVne6thGkbaekwo9bqc9MOBE
WM6di0SrAVQKDHI625e5rBDUBraCRMaK8woxYJ+JiTGuoOCthNuaTa3a0vMEtJhr
NjZQGAZFayhbG5nKU4m/JaWqiCHLZssD9l7/rqj5qobB+qtvAfhfcp/Qklqezzjx
Up6nmR1aUpyuuuPI8lRWXzR5y2DxgWAS5w1lJ1thH4RQ3nZhHON888+ObLDNF8Dw
cGRXHw4ZM59frznsEGhvtOj41xL7lYl16DykeVfy7u1dSHPvIDMJ/jmUCtQyQq3I
mK/aHhQV1qgVDydj9r/jSYNjELjU7ttBGG4YAaspaTkh0oi6ASOb7QnTP4xTXaPB
DOQwTWc5VYsyeLBqHl++2VxHmrSd6SGw2tcFyl67Jdt6doaKul4XXUg69db/ZWoT
XDoKO4WIP1c72Z1xe7oKiAMqdWO6b7L7Sy50dCQ3PzBthy/TJKzLtc3FxUAxos3F
oO6sKQJD5r6i4UMsUYwcajudq/4vGJzbbrIcIM/oj4R4JFK+Fi0Pt/kjGCtVDl6j
r4bN8HMKkozn6REA//kZq0pFd9pwzIhXA6QYHBa86Lvc8+ufflK0YpZB/58FuYrm
qDBZSLHST1HMIs/M/A1iytbBBOOdWbRUEzwnwe/eK5kiFdUQpRK6bf4NsfbqJO9e
6UBaoBb3lK9WlQDeQnSBZKUXDzBisbEaLBab/cNYf9SYI9kV9f74G6rkKFf3Jnl9
oqzfC4ZAUvgIib2QZlGDJ09yELA2UI3j/1AEHGtsNm5Qvf/LqWabjk0R3/30LsNg
e63RNMwLwxFfQTjgppWLtpm5WhhJ9LvCCJzhLMFcmDGXuq7ybX6ufTmxIowLcyvR
E2W8PiWFgUUhzBEqPeDhwaDa89ZNHcskXXsZVG+vjSzVeCNgIEXmTWdOGH6EZ5ht
85Mh3E5ZQm4DySMUd5+2AnFDwsWRLKSCz6hGWOTOiAKXBflgwDPZK05WfHFbPqjA
w3MXbC5+HGFbQM4gaxfUrwMGsSIPBP39Xd/fKKrOyrsG1U6GKm/AulGL83rCKu63
D7+x8MffNXHr3UZUBuhi4K+A0ZpBX9ifojLtlOQE6H9bKmgMQgvhHNSiJCYRxTf3
TGUwdOyTUpBU3xMbKKl8kH50FCqHTMWUqWjwarTbohfgE97Us88cM5WI6cPCIzkf
c8WjiDYsZmfeY3x423T9GcE7TaSSTXfdszPOr16shwb7VcS/bCupB6wFXUs5NaW0
3rU3zzXiQUn5ZbW5AmIE1cxtc0CxycoPwpzgskhQnsqxFxcxBuuxuTJ1OwfkhfMB
flz2z0OTXxY/mBTYWHQj4FkBeEN5MJ9VNHkHck/+XeekCDa9a9XoZWG0q9uUAbyx
sdwtmowkVd88Aki8oQ48zKgtlroEFsq+Kmlvkt95UCwjSVWN1nZwwt6ITGNF4LdJ
dEOiLzloZ0RTFxhzr/ni4iZP1OqFZLoqPCG+nbSi3QzmLeVshD+eAxI9ixFHrsGb
cGFCAThbTJeYiSxKZO+YAxXMv3/tJ9XgPWQG/3oCT0uhXA8qjBnOMo/yTyL2w7Dq
9989hEDU2AFlWiqoHeUFVq+QpmErv8BbiEia4S/3/lJEsrdSzJiRWhCJUEPyEZ1C
xj54HI6pNdXau5kwzMMlcD/Acm/Mog9o0Cl2HHhZniNdCfw7lHEoEqWp/0KobyBC
6zyEwe4CllTXR9h6mTkzyV5reIVUHM6xHElf812st6dh1OeILUxafsFZCyxRkOza
0B7K1R2zcv1/oyk67RTyoMogiGoZ2xXPuxmt+hX2Nk1sXBBbBJdHkauo9B2GMqGp
iIhr9SBNzpp71Rzc411OXWXwikDOxxdnAGu2p1l/JsnqqKUBdiIy/7GDVC2UR9Gw
Sg1d1PqQR1P8Vui7KQ0uBJoJNI590NrHpO8qOd8XhPQzZ7Ifo+bA7kiJZa21nz4E
wwyiBc3WRWn4/2JV5adb83frT8Jwsq34rt3t5E7CF3ecgNN55WYFjsyqq0yJk6kB
xqpNZGkO81t6IQ4kcNA0xf7gV49ULFG6W+x7GVsCK107guSTihEFwc7283PGAX+q
sFkQs+dsLMBH2Isf6TVhmVodaFaZ9eacEtxyMFxFG2Bthnd1bkgHj1YLL8N7ELtn
nUwCabQGv+7uLqGzrhAMLKRuJuQtzQml7xewewmeW/1iLEqLBgY4zXF+VzsTiF7Q
71dfHhU3NyKLU816vucLMx81y/xeNjgSIvNN1H63anKNO7azlDaVU4OLGSLCdEuz
MHuC6rTIbPkTYuTfXvYFNI/Fe06xZ4nSO5Ww6Hyl9eJBotZCIP+GacDc3ALJA7p6
gSx14W6dbsXodbM2XgXJyl5R/WA8uEmJw2Jd+yXgraNLr6iTMFWeguHfmGnCcUw2
VNEMGTx5vwtlluWWOwvWlZ2ixy6cNOJthQf1kkryc97ud4WAXqW5p/uqfmUNZ7oc
jXOM8ZQqTEy9q/FQAKi5yklAeuyBlP/3YgEjTmBmUoGO5a8DJVS/oabSfHpK4SKa
4QQYjqk+orUTXCExLN5GgKDsCvmAxFkhHR8iM/U6qbv1Az+NJ6nx9wNeGXR5ARfO
7e0kNeCUeM6xOzgUkQowpqr5cCZwPd2ChvcHmkYHDOmMltsqPlCuCUgQ5i6NNxHU
puhhp8pYAQHJFAA1tEBFK/BGnqSpDPdQGvNfaEhWNyyAgbEKncj8oHz9mgb26gcx
idnC6eOAYQfHpkarKW9Yy3GD4mNNzGA2aNJ8aqU4Lwxd3DZ43YeNhtJycis/rX6I
pejUCCRPZL5wT8R1P7Vl5D/4BfVKQUvXw6aQ1+1h4LLadwA78GYvnZYpl0KZg6zD
0B4JtzVQwOa0/PcePVKGVvAHw5oya11zbSY4dwF7LV5jA4PT3voW1ONXsBw36fOm
qbkObV3xfkTCZly64HZuXprjza/cfgLywf8TrYmJUSki/7zRHzn3lyVJD9PIdhww
FI4sjs2NDmJsy4mTWL2RqvMJtkOa5KAuAhFAvkcWN45fckE+DvNfq8BjAdBBydQt
C3dmPx+WOWqOyofMlZG8mC6srblM136aAJVEGlI+M7V8e0gOIBc3sk5SiD6UDxia
ZauGNpH6fcpWfxBIszQi1/Pp5JypU6X6gYVmkkI+O06NZdBQAasFNki51iiiYdh3
CyMzzpQurOjDAOBxOo1yVu4pr96DiVJqr+AEdP722f43JzQyPhVshtmCdTtpfcJQ
amcW3xSyLsYK7EqFUj1qvGLv9HEXQn4A/jUHGNLiNoTSSkUUykDig7CeviZJWnLR
tK0aZPN+vcoAFjAVDIlrlVaOxufkqi68SuHGFuAXK6rgWmevmgUjPPKt6Hwijqs4
6jqYJ9RCV1xvKGdXORORiooOoh9VJ6hvd5ov6fyPTDoH8Xjt185zGeLFCt11BEp2
OPR3ZYflz8GTUJ8WAaQNSKFtBdePC+8ZRfET/+YZ9Rx9RysHL3xt2Uc7aa0eUrk0
kDoT+ybgbEfq9ZN8hqkYqZZSBHwQJQicf4BbuwFAngIW5ssBVXQCRfeAwRMc6e+s
SVbReAsRcRmhKUxOeO4CA7ljqrNUZn1A8sYoAkXIngvEelv5iMihC2Q9ukhhZwut
6jJK/fZLV+KJz6oZBBUsZePJKTn+ErAE1dnN1C53RX7aJZ0lpFX6Djic5mT0EpWk
jtRuOMMnB8ihULrGlQVB7o5LSbguUPeZ0DEv/NQL4WXGfM2i1h8WuumKL0t5YkJz
jJqQQ5tgfGu8m5xCMLMOT9wmT2Qkqvr+Obw+W3wk02iy/5pNucDUvg6rQeZPg6LZ
A+QWlrDiEPbHn2PAxQuriAX42M3WvmpMBRSDVjQriaq2iHV0fWMpyPhOAlCxgXmZ
/hWj6zaaHEvqeaMBXCADLBEqORywDcqsqf749iDD8v7J0yCJthpdXVXxfVklFN9L
R3LXDiyBKPHe0ihgC0oQJmFiPNJ1D2nqQDjMAfIBiL/GVjTOkMMaU7Zx0Ujs0APO
PguOFqFccgQG/VmilJWtP+9szGs2JnHlGz/RWuvWPAYKJlVTXCxC00yXP7fwj/Cd
EWZbYVUvdrYktQavzfNqfLdBoddWAMbctX0znaqiKrwPdv0mV+Zfd8If6ervtVj4
/cL+d6qPrwrjVOLUlUjWLLI+wT2JF0ay+JHgbhR/lZw6qxMKoDzKImXUH0hQJcXC
VVDLddqlTKBxKqjgYoGdC7yJ55Ha/Vb3Gdky3uSBmT9xThi4pzI21Z2EHPta5v+L
ivOOpcX7Az11G2wWBIJ2c7FZijpIXey7zbvF37qQu2m5ZevXm4cSGKm6I/QhOnTK
WV3nO2TQiiy7TKmgVCVCgxml3xbBS8ZHGSWtrSDDpsf3jekXKURkK1qsjDaAjCDQ
cOuw8aHsTe0S1YXBJxvN+EiALwvNHjQ1JGVziZCqnvEIlJ5VnfUvmIHZ5NuvlEFT
cIuISgVvSE4v4zUbdhg59lfpzkwU3dUkpw6ILOqPnwcmGfouivh8lbcOBBHA8rPu
gJbnQkiP1dA7JbJLYWDcFA9UHSCRvyWS91QRBNrECS3r3cAq3OQJSlxhq50H5rpi
f/wq77IUk7gr4Qh/63w1GduYiRHMkx5S3s1NRmlADyS/uJVd+vumTDruFqOA8MEW
4YGZtPUsvq6lCQSh5i8u8GkDemj80mSqclKOQn3E6xRfXtc6mGwV6DweA5aK68L/
L4BFRQ9eglcgPz/EiKguxx/QY1kjhBiI3gphMB6s42NyxMSM+zc8Xhxw9iFBBWd2
Jq3qS1z20Xyru2RT6D5A8v0g5uM9nWfP8FfwemVYRYFmEnqV1ucjvezoUGslJRdA
V1bkUgI9gA55n+A3YJcEnLON0+/575iwq407qdKB0R8ORiEvAfacJqe165gSqiZZ
6D6nCxuz1vTj/ct0mBtFGAqcAektPNJ6jCprbHQfR1LSTrrrZmuaNIhZnDv2YaVm
uN3Ur3O+Y626RCwgIbivmCrPns6QeCr/tLZBlSjrp7OYJJdaiXj3D2i80wSRuNL8
Q2x9FzvkF4f72OmYjHTGj+KXPk3aHSuWecf0d+AIttNrrYCstadbQBlUKwaaZ04G
04TGgI+FBqZXuI/5BfgcxQHRQfmc0c/BdJsG2TE3sG9C9xarM4PFX32q0k+5BU0r
VFKPfW+NohLmFhtAX9HtD7QEHtTJMhcSMY5HC9lOtUAhKCr8qebWajFmzpxgujo7
5yfMpCWYYp2JR+Kz6O7peqbMF6JwZfCh0FO8TB4klOozB6U+bo43Rm9/e02EuOuN
9I6ct9SDA+hulCsIcHE72Ogd3W5UmSfB3zQfB7t0gjnaBiDJ5wFBJvzrPuE9OyH8
szd5xUxlL+qZdB4ELgtYEmuePT7j1rYfMbS8gKopEymZmRjTLnJNLtRa3LroADvX
jEBQBgudrJtuw/vGgCYhCFqHfurf2ZQtAJc2ivquwK9gysseVIvOlyYLYfQUyKvV
Hg5Inyr6LSNnYRQWfJlxPrymmgrgFAsU2ESSdJ60iuOY8flZEWZqGFCBUdtBI8Qa
hfByjRq1keswzioPsDASq+xFns7f9NHIloKbNtib6tjkZdyYlupyTe903C/9fg2r
j7xiLJRQKlZjowY7EgLoLkIr6qpZAzcv5jFMnXKDdmUnWTzKX4MvHc9+HJaGJMc6
mMzEGiAuLo2hz/YtSVWOUuIqGA6aoL0UId9/Dn6HTWDi5anMNVH7jALuoQpY4q7w
SdoALNGVa1Zy3xPcqWHPBN5gZ0vt46Yuic2bHv+htL4kMXxah1iwdybXMveb/o95
sWC1M+UTck05Zg/8qMdwpIx/2QYU7dKr0P9pBvi4pkXOggrMYu8KP4qrss9ax+7a
lB36wCwqamfKxvgVP8sniMEMvas592/f8mGJ44hXxT4dmSkCDeYIJq1zZq0EAyHO
bJ57hXJZaZA0phu5Hepguv72pox/v8zX1jgRmyon0AV+vBRNkj54VzCIAehXwOA+
XjG42bFz80sCEKR04QfYcHMtQ//QxyCxmWhbAO+7V8KPbnNG5SPrwsP1zQ70k7RJ
MPqDd/+ten/u6/vtzZojn4ZSz6hYmpLA2yC2hOrCZjGRBh04f19V6A/lK8Wz3QXn
DNHdf79ORcbwVjeowmNDNDk5O9CF9HbmuqvOGqEv3iGWFfVkr9sZp0edcWFnZS7W
WO6nATaEOcsDciVMQdmnxw4qaXai+huwMFBWJiUfVqi4xHm0n03ECGyQlwTy9ryD
7cLd+v7VfcOSXBE0tyQYeFCmEgiGxs4bXHzTRNCjk5Vhrc+E95wBaAzc/f14R9YR
7FYJ2Q2iE0m9B+M6xrhtenM3fksg2dnwjEOEDckvNh0AQFswmryDB03RpkZfNWV1
2cNaqNj/wFALaZaLE3dpNNb6ZoGs/yyGS/88S9o2m4IBVbEHU4u1j6mdJRpkq0cC
nLoQEMae9/zmDGcROTVfvUHBRrN4SQUb7b0FPMabRhbzb6yfIL1bidjnk6nxLV3P
N+delQ3fImxa1ToCNfa1ie7zgl42E66R6rxQ9V4KvVzdzzeFUwKmPK1Y/pw08ktb
NgPjrmGy0pYsXge/4hCiTDLjI3PfrXavCo24LCy+l3eTtywj+5AgvM+eaXbU/E5L
tq7C8sus+CTGgnDeTZkPisEkaBbze8X+XOLhXfQL5fHduAqnqy60LflVn0kOfc6U
ORzFnPj99HEHgjtxfCfVEKbiiyIuZ7mPZ7R4wWgp58eN2k1jzRcnsp3b+Fd9WgEM
vOZMuEYVJT9+HE9Sbed1AvclaITrJ2XQWniSzDa2Pli6upVOBQkpf193F8CTTW5C
JZDiEn0jgupidIxNPHsG2t/d0CePmlP7iH3AgHTYnhWHNKseRLlQ/XzlNgBcAzlo
hoqfnqx87VymdcYxRCFWnlgsbbU7LEG4Gv+oZohhCiOxpVc31qGAiXFBDBzu5zze
ASaMXtPjtpE3BtWfBS7oPzk63nnu9kWy7FtUPni9XscisleO/Yh3nGVMTfCUXcdy
Im1Sc7z5FOlVOUQQ2NQ0Q8HGDBYIq5N49jBndQF5UpfWAR04AHQRsAnI1kBZrvag
uxpVEqwfSUA0lT0Tk48ojBD7pexm16bV2/9IAgvmjoa8slzn506BjL5jaRr22nP+
k4XJxPDnjd5+tHs2amCDw2YzdZ8A+00HypQ8WPg1GEtznQ5ubs+l0Nk7J7IG5+cs
mdLxY5XQgeYRNkQVNnLSvu96HQoiY0UELWYnfjo5rd0G5RMLum3oTn2t8oDQytcN
clCYuqxm9tADxCtTYTsHKWyUStDkH4nXGjCaENuzW9wbnpScie1XjfEMavdLKRxK
7A41DXu+LhWq//aFIu77uYitdNdJ/5qooGJx9VOCPfPt7+CBgE4Qn5gpf3var3gQ
PNUd6DlV8x6BsiZ/DXU5k5bQnJhr/aEfq+uD0NId9OvNP5PR59DYJI31bg4o/LWe
OMJF8yHvJZhWCrFiWBhPpJmnbDgwikRmQ0l1Tvj/YpG9tX/n0+3RJQNj87vAHN7k
7lzmBuPuilUU5i8K6wY9O6azmmJgT7f0RvepRwThoLfz+4WrljQzjkDs2whBaSAT
ziUs/a1lFSAmsEsgg3oIj6IAM3KCx7gqraodjgIFQfB8G14qwWuhPh8hyhDxo5i2
nyUmyawHgRFYZqvyr4KHhVhL6yrhkIQEHKjlwN80rr8BqAkGg6Y42InF8PMqt0MX
J43V1EfHvHjTqUMl4Wy9Z/ns2doRre9FfyN3Ifg3f4aFvD4JBSF8ulVSdVOsrSY+
1jzNkXlINUX8HWkr+wcjQEAzd9nVi4e3zSmgkeSivPGboWG5u+chhOznLY0lTvbz
gVSQSocOTxZ/XrKq2bA9cne8OCSYPGFJZwi3kUKghyvUvxSeO5wxQjHEvJ6i5/x6
5nue4doR1S3V10UvaXws++tAjHTv8XVa9Nk614+euoALVjFQyyhhSbW2Wqax+peB
JzDFu4spBhBrNH+x8MClYcn0sHRZiOp6LmnwkeUQ1sPD+67pRZHL2TyqygRQzN8L
2ERhjk6/0nsNWo6XwNQiCCXvoJBdGKto4KH6/Nh0t4Tp0lbxLTSMli4mBCYhxQMp
Oe8b48/bCz3mBSIkrgbntWhD1i8hYjyrHbkXGh3jnqX0bAiXgOj4fLnHRZKCLS4D
jrbMRfiUFYCRQz2a89+TgSmHe9+eu5VsahZHTyr1omOsS+GJoG3q7VqEEr+kgWGr
f0bDzXaER1xrSagIuQ70CgJFYePYwFdRNT5LpLnolFGz+jotfPEnarIVRBeaMPSk
vV8eku6ykqgT9ha4iIClAwJGVD82D6emMbUHAXf1yTJPNApFGuMEU04mekaUJ3Pu
kkNshfzT0wAY6phHjpBoa5ZFLdLFUsws2OeMcjTLorYmITP6PPCQlsQGvehebBx/
qg19UA6CXVlPikO44XhC4Bmqt5wDkwuCb8u9/PCxcYNhA7q5rLiZc9CT/QQLoYGB
6WyOW2sGfHtzpM2ke5QvHtPvUX8i8KmRmnDOXB2zcOgCvdbjbFdkfX1R1mJoz8rG
w8yo1p30m/XFym64Ddix58pYs6Tci5UdgWb8YRD/sgf4gDKdr9iemioFsRSG65hS
2KuWee2jzXBYJqeTAPdY4DHeQcjRLMyQ8hzD0ZM7RsUgfOWmVBzdDREAc55gHI8I
Zz8OOSn1bjDMgjEWC7KIiozvDOj8g0Oc0fwWKUo77Tu+xCTn1EYxbulYiH8c2PUH
yJ/SkunehSIPoXQTeI3wHrjqTWmzawFUmc7V7ZeAXet8/TtrZOiRRtQBrwwmKXAg
OekzeR3Ji8h8CiQpflvc8Fhbp39J3y1xWf7X+jRJHrw6H0TRj+IqPcJXrRFNkYn2
TNdSzcOylu4sZR/1TYbYZcerUtcA0tNeWGeFr3poP7XE7mkufBcoFJffQZKX1Ceu
NSlCPUFprlLz1gaJUi/hxWFwj1qpAUU1Eq7NREdzJxSwzlps5rNrRXy2YD9BNkRB
oN2iM1u2fZMd4wtP+L7MhSomw+RD+A900UrkkHVXZhEYBbMMXxKndNhb6HQpHhC/
ZjD0huC0aFkbWErcIHsC8AXeQMUPdxlOhWifeiTkBkqZpghmWNX3CtLryzazIKNz
Ql3lbPeXDaPSpnEnpwAuISVoDn3Kny1Wt2NAI+P0pidfWnshw8JJczKF2v2XGgyJ
5Mi1EBToD5noUEKfitZI5eHm8wgBk1rqALGcVDEmTX48EuSlchU0seZ+j29KtcnH
yFgHNnNmAXMlrdXpxU+vj6f7kO2X5CogTAKzr2ZRek1N/eMatxxS9M2qCv85wsST
a8VJEJKTm6GP/wScoYQ5Q5njHNq6GfncjvsPnhK11IByKE/AOVVXxEBg/ghHJb81
R1ei1H6BUVumOrZ86ez3lSSdgMZf0wiUWpq8xPOLdRvqXl/NuTrXfFAiLJ0Yo5J6
aefZsJy5sNNjjwiA2V9o+qOMK6+iExYkLlIIbpXe505iDhjje7H39Xwhp3mtEhm6
WWVhWV1lMS7LvbQ5Uz515thJTECyqbWR5vcaTJd3wRnJ+fBvOjkh6MwMdIaTX6Q9
4uMav9WzFgK/arXUPtIRXXSDqz5YnNQaNRGcPM0rH4Q+2KRjqINsarRQvk1q6rSz
Mi5tCmxqvdaX06Qw5xPZV0308egwfPnSrGys/toGdwFSH4Jh0MoxEKcXGu5wjIFs
TZzzLAHTsAZ5ZHpWLSHNnsEeRB33osJejTdDguXEMQngGKjT1G8qGua0TNz37zIy
QPCF1knwqsjjfq9cabE+v69kLakC680qrG7725JisEIdgMu/HkDkv7QS39pLii9W
UQry3ZXfyBC2+js4aOAvJetrw+lG1K5xbKSaDr3S04gozc6l17UYvfIYS8vpMc54
6F7w9QZU2onjbskB1VPc+HuewdqyrgsOEtZUO7aJvHAYEcQ82so9eHf1TfadHlo0
qNdnsT46Fji5k0hEj8Zn2eigIgAXygPG4D2IyMKTaE2WFTocsoH0soai0dAq/XG1
vsEh++MW5anUfubwowOaErfBOzkfGVJwgOtL/wNeexa9YJVB4FUoV2kyQG6nxiMr
aoExRwetuUq1Yuyl9Ug8SH2yYp+APM/LTOC1bhCT2fAE73xKx+OUPwRqm/3ZCOl+
SuMIpji8WnJKCJp2RTy/mpA9skUuDGAIp/61LOaWdiuC513/YR66nLr8jl4Q0Sbl
cKvX4Xc1SKcjkI+/kVjEoKr1M78osMVbmjU1z9Dza/X7gRxX1H3XpNAv+yg7ajsC
S0ceolzEqOOostn8paYwN6l7++mUrM7r+X1ful2lHdhLqAi2LUCv71Rp+n0Lu+Gq
an04S/xjWJ7KQnmTtxGWZiNhD2zLTwa5trd21BgtdlNUdbSl+ho9iKnzqSlwk/4u
PdLpgo5txCTNIohbPHpjuSwxNJiIQn8TgBIuWcqWk7wkWYLvTrafQ5DOcxr/R3MW
5qFMEC8/b3NRoGwJD35s06I87Lrr4qSyy54aRT3yzrb6qk3yv354t4OL0Koi4Ogq
xakhrQy7vVFSD5uleBBrNE42m3rbsahMZVOqDEwcCqvVbCjn5yzYW7lU5om3gOVD
BS5pwAxqrAlXa6OcZ2RiIyVNPhfU4lVSgC4cSPjv33KIgZXqKyoPIhQgBX4foZHQ
FYcOZ6B5uhhNzOOMRgutBDBnnmjYwTHxfJbFMftctqy4fooQ6SCjsxwmZpnIIbXs
pB4Wbv5PDErMBdxT2i6BwQl1FbA/XwiGZuvUvsubAG29cCOYuldYlEx4YXsWAn34
+UDrHdGiGK+0bucc09ZLSgQ53dogOR5lDJd1P9dXZG9lBR9bvkQ7S5XAZCAFZoAv
+L2K4wBEZam8SXd/k2linXQAJCWmCN5GR9hZkmEFunr+z3oK2rG3fmXOuNdEwIj2
viXpGJ23WjBgP+fpV5f/FXe6YvjNnPsu4wk9E7pxHxaqIJ6VQ7UrmRiJrFcB5qeU
jqdsriV2egAVArGwA4VZg06YlFYsblLQhtUhkrpzL5TYDB8zFFt13xLNka3bfsLC
QaYscgcg+UIHt8VzEn+7WPyqskWUPqfv4wr1BGm8F1NGnnMNcwYXy7Z+gR2sU0/h
GvMwr9tmWiSBwrT8cn1SO37Fd+k68U+FV4E9OQn0v9ZDptxywpWkoQf+YhejIG4T
xrqhWA5RfTorogMbotnuQlVjdW6UqVjGIm7arzNv3IwoZxNaZDttjR7Aw96VNynx
Ym7rnUY+01xCP94ZFpSprdWqp/lcvU8nFecwYNaXOma7fBlP0PBYNzEqsiKfYh/i
rcaAQgp57LCTs9yOS9qGPXEowJKQv9YMJGtAueIasZci98p1YFkrRGLmJHO+o8lv
oXwxKb+Z7WN4D2ZvUjZb/kERLngD1aCII76N9BdDlLuHGgf4uvGRCB4WD6poUiUr
eTYz5QpOK3TnCo4Ptac7rXWX9Lb58lGEJVMcERKs5BF0Ak9XVrOwr3ZCmqSCN0uA
0xg2SA6+z3JyYGQgsTwVSJwVMlgIx4h+BGO3GKC7Stm12n1pqeQCS6nrM2JgR1Oi
t7k+Qq/6s2G6/8YAhRhXOfBWp9QJFaVxOaQx41xtR5itrs0XHmRSGP5PvZOCzIIG
em9Xeqlj/mEgOt+Jo5hR03M5eDd4JlJKDNcBlkv0HxyJ/VzuLu/U+lHBvdlOG7PV
12ME2N+v/IUTpwxxcxOQFNG/TDqtcUGxjgX11nznj4WMK9hmBDRUlwewKRhmY6ad
cjSiClh4vAXFH2DHsKD9YDq8p+/jv4CNwAXN9tDkKNSaj0/OFdtJffp55wsRNqRN
xYK8UlCHncFNwOhdE4WfrQYYJJPZFV4w/n2iqX5g6WvD8R38+eqji1mLWgiWSRLT
mJFKdW4/q0i72oi9Hi90+KVUWTU/gfbHG4jiK4S3tD69NjeSVfp1JEJqUUHWfC6c
TzKOj1ILb8eD0hwGbgf8BVFlBquCgmRh7a/sxxxGdmPvgCqf12YT209aTU4zRkuu
G5Wcwo/Q2MqqOPlz/8jYTGWe98MnpW3tDPGagKiJOD8nMlj4xJiw0OS7BMAsQRSH
jl6HLT3QqCQ09/IGMtceHN3iGoHKIInL0gstOJPkeeXgnL1Y/ncq76XHAAG8Ud2u
sBipqgQSWjtMglEBY90g3NcLk/PxZlOpD63CijYDksqdr0u2oWjogllhs30htNdl
PC7MaFp5X9aS/lmiiOHrlFcwpdRZrVvnfnzP4MvLQA0vF60gV0Z71gN/SeAkembk
T+xCBdbsMds45d9eSRmHRGPyYnDukBg+n7ZbmM8RXbcgpHP4n4Llx2vaAQJdhmYn
T+n794hk2R0/tsgTxFSFFS/IpbIRfaHwB2YswzDAdsypoL2CjkCOpVzNBKKS0RFx
IxSoLoPV4Dbf07TWCCns2H/warwpK1DhzE+8Avdm0R9sFJ/GCkTF9qm9Bpi2WEEK
QP9pNo/TOlbtNFP5mDfiYxaYWZwA49uMgpf6wFLS9apWY+trbI4xYWzaS/krbOYH
Prvu2aZrQxvhAm8tKRebvsFYhj6AYwCZ8qhDKRW/+lgi8nkUSAd2n6+H2QLfbQYz
cpGelSEozpLkO/5e3Dy8ODTHpG+9KbsaOsEoaoSlmj3pCCldAn+MByJCkwp0vGOx
iZhElFdF0r2hWSjgKsj+sxd1WTHugMXrD7kj8G41cU8ShwehDUcd2/xUUBXLLWjt
genAo/iR4ZCjIlE9mHNZeQEoFl0DAWYdLcnmSTbD4o4d6VmW1QkDnZJzASRJz42d
o1hooHKAIh5Xh3kcNczNN3DsPSAuuWcXS+TMyoKZIMKImj7p46xZtpEWat90zsrq
of/zJ7tONaBh9Ds98Zj0bRuuxT+ab+vXq/Y26PwTzmEp3phdReLduJ7DRtXqpXd8
XsoN9e9z7BRacAva+bPEMuI9pCawdFlhQq650HgxuFo9UoUOm3NzTit2dM++e4p6
XaUVdhf1zl5En+d0YPsjmljpVRKlthJLzVxmx7pOak+9adA1Y8PIMTcRcbURSwa1
Uy+OEwAGR2Zhg+ysLxHMKKLvXSFJb2oq+PSRdMfBgRJYduwWG+rRuZFeGwvX0QHD
KJIYBclgxh7cbUv2tIvo4fbhXcDVWE1KwxOhvhaSvpCwmA1ye2hThhDpfhuZhUOj
fkctjj3Q73kemzGjiJiMADJ4xoo1/ahvicGcPQ9QI3TPh4h05ECQNpSwgmV9JLEh
khT04Vvg8n20Ol5xQAzPYeUUWzDtvgaP1ROtWKTYhpwY2ISJ1ewg5HMOnYwLVMRz
IhD7mpxRXbFVi4SZ23lIn02TG0YV1CVkjrNJ+6SjEIiuu68G7VPc7eBL392G06yl
LqSgD3aGs8Q8DmjQoA2940Ut8hvvMi4mDqeZWSk4vIWhfYfEaR4iwv+piye7b3n6
uTdk6bqztGoRiji0Q98KHY6SE57xBNAT+dUUeHjki1KM0JO4Dj2nWByLCM5xD0nz
KNX1FQ2BHP3KX99oCynszWW68gj8E1NuwaZnUup0cmTbHBRTFDglwXvVc404jr38
EYkTaiZ/f2X1XFFIgqbiXg66FrNhQHnXJYTzjabgIuyq9xIAdCfaJgqn/6sanNxO
/dHPrc/beCqB4KeLw1k6MlLxzTQuK2SfkD2IbZ/NUVFl1/EbNQzQjPWmvINe6M1k
sH2YP6vOJRefTmE2ixu5eAbusCrCgKGPYzgE4bCpPaxutzoPbiNre2IxgbmyEkaF
RXitE+S9em3m4hy7gvejOLpMFpI2RLaNQO6byoLWncmalkoiaeudPr5uBYXXyeZR
zthEANn5JCKBOqgQ2ABIZH9dJN74I4/J0plx1hNaw/GuLCTCRQ74hnptX7so+19M
9M6kzyiyifeZJItt6doYVYjU+9+XeAyNNJoY312lji+APfOvbvLZOsoQ32cBxs4a
i1aqJduRMzNk/3jzszJyz4TNG4gm6nyadSJmrQpxPSnbQXqWLFanMCYRNtRRr2IJ
tiG+63qu52njLOywcI9cWALjSTclqK2CCcD4e/l3aFvIw2df6wn+7JNDsz1gay5m
aO06p2UX9Od+eosG4o3Z8cm+6SQii8OzsQ6ZN3QP1ABzvY6KKIhQ5IVQ4k7heo79
Ic8+yvyTVfeL9nBiSUc4cyNE94Us0brLXUUFMJPm7I1hyMYVfgDA9mpeN+YXKDz4
+EozZaTAp1Z9Iqyoor8vJ2Xk8OE82tXbb/JguSU1mpQQrnGgG2aZz8j2kdVOIKed
/1pM0LVP9zt740Ry2GhDfTVCfXXiOo12S4DkPSa4p9gcfD4imorpKYSsiNBSA+VT
yThfRCVE89Igmfm/QsrGyfglBhaO0eph3mNejNq6E4KnwelTwzWkw5/dFw0xQMCw
UY1oaiOC/QEOa7fXfQiFgJI6XkFC7Jlo3f4U1JtfjTPWpRyfcb7itpA2uhO3VLdP
EI2qnqLnJt9UdB22U1ck9m9/kbSrfG+j6au8XjGx0QkpalIx0EV6F4Yg5AlKQWFO
gZvJk8eOPXzvk4zwr90Wnb1oWAqcypr2KLAMjCnKAL8i02ILsVSW2946p2EBb5ag
aSyQUP+1DUIP9Qi3XaGwJ/vrpV1wcUW151BFOIlnCGfAd7W3JHkG6eHA1Iyx7pU1
g+0I+REfmOpdTp9RwRK1QX/Xc6xbSEBjcS7P6bUsg427Z8PspSwiVTgtjRGK8Pma
mCsNqluCbvqdNhYM0nTL5NXyqxcI8FMyjuBTLCGS0SP+6hEzhdNrU3wghs+fgSNp
ezeZ2UUAtkjh21oH2OaT+f5iDgG6hUiAywuIxXmLvVkhAL0zmjUjVmOiZjgc4Nbs
9VRt3HkwuCM+lXAaz9F/jTkxBIdssIPBHuFlx2cyAEYjWz2OMAVNGYKup8vCcQKf
HSlsljgzatOPhwvjB+fUkoIJTch9ZJSjaZJD6UBQu1iGpTTU6AtHKxUeGjZW38LB
QPBhZpCfYYVdsSLQVFEwsQWz1LEHtVzaWDYPuY1YoFCawFar7lNvus5xwJeZMBM1
Hhvi7jvByAD5il8+yi2LYKCCpfAZIs2acMfr8H4Rv7Ir1Ju4dQUvapm1PiDOdhmX
eBLaWKkmE+bqOZT6uVJ6y7riaxhnmHL+rm1bt0VcvfsfbvbCf+Eo20d3YJvEW1cA
2DLEgVSJJVjtv37teOUJIu43cRn7ky9b+n2Gj9roY2BYau9o31JMRV6hI920pElZ
QKOTnMmjsBhGpmCWkiOz+6RCzXhGsrEfjsmY0WzCgU1AeKaC7bmM/qq/veyTGnCl
mtRrW/RcIvR/i6iQ92V780vxPWbAz8KqdRjdvi07pnjeaMJmNlPAFizAdq5UzUb6
GXDCBmlR9arIvrg3hjaTyCS92cKTc3XH/lvHeWUb+5fCabNwQyx4lYZR1++bzzIJ
eRtXisF4+Y+oKJEH1SXVhsuzOFjwyESMNbPiO9XtGr+C2lO3o4tc4/wnBOZ66bbK
GfRKnXaoWrrIC06hM/Zr623Km+mILbLM1LmzTjlbUq8whNdcNSM/UnJsviB+ZzwI
zkmCpVFdFw2vA0US2y2SY5WX0zlcGOn59EwaH4kbt2Fni+tldNHj/eTL4U00r2cS
PtXJefBIzrsR6JOJdV7ezcX3IkIgBL9SbiKbwXQxCEHpbsTn5WVF1M303oRxlMb7
pLtcIwmU2Vmjo+rYtoI2DYtWoRB+7J2m2ZP3MFZ+ZVl+rAqBqRGFXDzuYOk8e4tg
WEbXRKegxSCizMW8zAcw14TmmZCZ0q3jTWI1Y8nU2+oJDu8aqjXGvrsNdHRg94j7
FxW7m5aDZcva2Z7p4oORKqWKKXQB0pdl9hfDEVYQ7mLz/KohKTjvnpdZFbQKRDMT
6PLa8Rr88WchgN+CJ+ahnKWSUGc0VmY7IG0mYQd0X+2KotO16/pxM5Nn+wAfIT+A
C1NovkSL44W92cUA2T8fTBk20K/mKAQAQjp5CP3sNoDKZR5EjA4V24hA2Rrhhl6K
vVXs7aX1f0hidz80qH60dwEb8T5gJIyw3FiKbx67RtJoNL1No0PJTs24/37uhI87
SRV4donEi4AjfAYWob5e8yKo3/DMN1EPEf570cYES9nP5Keo2bZKWvFirOw/4js+
vAt4jOlDOWpMS15VJFouGIuZVxyuktQOp1JrBgYsg+3ZdL03T67T1WX24JdoH42w
uZmRiaN9yS2uIGb9FNh9DejSECUsatlqJEJHDtgWCZKDGhdURqbQ/g4/2Wznnt9G
nkZGrQZm9zAQHMnQV65iJWAtZFWSqzPL5yAlKPu2zGVV4HG/8TcHQzMpi5V08Wci
GotDgNPpSJgSQZJkrtzj0POBGANysq/wcdUputdd3TidOYH5LmPfq1kbhA+e7Mni
wImj9XlffdHwNeTJAN8I2FHAqtm/mDLeGtjxcQH0LFqqBfaH+C4ZI8tQURdNJgZY
gf8Hy5ZijL0iM2h+euTGsCS/jpMlIyxHKid3yz4AjGw72GaINvKh2TYC3N6JD7sC
SvygCtp5PqX/BdghD8STeihOUR+en1jFvvq/yK+851p8NdngBNLt+kpeT9KekZKv
oBHHOD7jBWjxC8SjKqXRc2xOg29q1+n71WscaClbLqle5HWfAIvZqfJumZR7aYcw
sPzqzFM2PdIOxyZXC4NiOkkSH35mRZPjbyRwf3cmo7iwXKN9819YKkwYo1moImOe
MNm79qJTpdR/PUxiP1V9OGQ5WuY0kf9svurlUxGC/eOOg0v/O9GvVG7Q9rsVbD1b
BUKAETn/5GTJgrF/LYrghQS9OmQxzPNdvIEFxrAvWgZRFgd87eKK5KO18UuIP8ch
9p6hB3PyqZJJ1M0IFqAgnKJhntT5K/TDhO7Jg4zuWGzfAJIvacSjgbvWw3WPf2NA
eRIJtDU9V5ejnSb6llV56NF/lvNIA/xXdfPng0RbJRskK85VDZzK078C7qEVYGvw
6nQfg1Mj9L1DOupv2GTwUOLwnlN8g4KgP5k11HFuKJ/7E3ifOKk27USHy94C8gBW
pRVGifO5MDI7oRKPteMD9R3q/RoYkZj5Ebk+I9BkyUeAnmsp7x9OOuuBTmfeRQpz
+zQNuLyMh0hOHGO052bM4XUai9Hr3twbX7hLyMFF8IP6wd0aBzohT2mo1H6sDv0W
/VgrZk3MdimbzYGEEYwawJYXkHKKqn5P2jKpK3WNMnDanQ9lES6iwlAh3zTAxRzU
mj11LhCGdMjGHVqET34ylVPOQRpqItZNdJN/jpe+b+IH0IfocSS1gO+Ag0G7L0aq
+xGUABMU5Pxla31lgf9soGARCDFGc3RkODT/ZcIr3plvnjfTXdOdvIRvCMRFApgU
Nu28/e5z1HozvaRKAFUgwQHjtQE5YDMkzEk1sX1VcMlauBV148K+TIglM42374U4
wGJKovTaxgW0SEbKuma0wj1b/tQA8yOPlj1RrMkqYQgpr3nubohh9BYuq0ywDWRf
5NVwQQKuvqgNCul6sd2OdxTkLx+JJIFLHRx7KDWE8goRh5S0co4GiKznwR3mf92P
6IrBvadQnuucnn+p4GmWaSSQUkQEejWW0pci2GlpbNRDnADHzOZ75NZxGtwO9hs1
b+CRpxrslmBc4dc4fa1MFAgPKCYYVH/ODmg+7eAA5YvEswtUVG9cYDL62FOjeuAl
kRtpFHCsdAjBljB+jh61hSeZg5L6BjCXZBvNjEtHmszOPlYkmVvmOqd/ZOZmXjqi
tcT8NZ4YKSsEdFBZilrNfKyjqbWZ8Sq+FNIzU701roB2CA6JuB9ULu1AaDFX4LT1
7TdoDh86/1V5/zvkGfzfQz9fJICyFntPEFlpI7Vv0bTY7ikJo3w3BeFEScj66wOA
eHllravcL5lfT7IFROdCRgMpPlxNBSMWBTTF+CR1cEdqbvHMk0ZDDx/ozZuF9u/L
0XpBcCvJZNwfwjg2ENeE9N3JHtUPJVl5aoD9w13tc4IGa4vpzlFmkaVwRkYUriNg
PmzJ6xraLSDpSaXREA+1tkwrHtpIpEwyNKTxAW1RPiIyPdWTmHdDnT6vDf9UXisA
7lH14IHbHk8pC9XLpKrknFZvdd589ZgQj+/sSqlzs5rOez3wEeaYJvx0ZgIdNSFA
KD+jV1b4PIDeZ7wFza48rQ74j5k9eCpED+7TGZftkoiAWYoyEf3rz1Eemkj/jo9K
DThE49ZbjIOjCKL3ZkXymObNAmrSFpRp8vj0qEknRHQGfo15wIt+dV2omk/Yjjus
/uvSkeJEvlVje9DnU7cOV7SBNZhsW65df9ckIbzuGifCA6Ga/g4u6Xoi5TJWulbe
BmNpZGK4SOOvaN4OeWdtenQ70p9rX9cHzdKjTJkdNlw+k1N/HrD3OWKi1PLlOFzT
ZYw1iTuPZaUfKsDior+CkZ0YrS3EHLJe40wIGiISTZxUu0QgyuXzCYC7WKpuLMKX
0wRuONE/BQvl47cexxOqmwp+beqaF5UkkaOrUiwgh5qfMU2X3r1PJoJZ7qJGkI5D
PN+gZwnU2Trwaa15DJ5n/Wspo3qWixZCuDbec87HYolyWZvU6Oh+GU0FvbtfArDu
jI7SsQBBRZTE663kYmdfwYXrruCaZIVw2HGgLnwmjXKMKbcF7cOmDchReH634y+9
4NRlmq9ZrMBwmGg6nLdsU4YEpjI5eXie05SwX3yA1SmWDybBalYG9YC4D7n+V1ON
0HbTjPy27bg0yvfckw0G1St090cb/IrDLZlq5YRo+Aah25T7s7pJ9PecyHN2Knjw
qTZQvJOsX4OwZFodA79DijejMRn74svmdhg33PnWYM4IGrUqJ3MIXMEauxQCxhKU
dYujXtj5Qn7hf69Bd5ogKXP39VkkFFuaGlANHfVQV/F3+CCHELRhLcXZobmQkmDP
K2yzArdzx2TFHpl4D1ZKLOEpWfCny3+gjkyXK9XFPaLbH3hFMJy3J3xS8MaJrqFM
ZcHs6h+yKoGtxmxPMyPeRDlAI2Azgvo/LWn82eNrtailL4nwYOH6P4vdn1oAVTwB
ODlJ/6FM7AqXFy/5Cj2VP56w2WdLVL19wW1AraDS2DtPI6g5huQbQZra/drhSnCK
7/SiJILsVyta6mQuQFURuwuFJK41m04dhsFD1f8O9CKTqySwRWb2FRu/dDMJ3rG5
k/zWMgBEzMAY/D0+Fe9t2OR9zJJUsg3Wn7k19+bnLSwlspr3EKpgMsSplY4iAZYE
c0OtFFv+k5+SC4RNnRKETxZrr84AFmna/ODgzTOITVjWYPYP+QViQG2AbPNvgl29
44eJ3X21p8i/2K/clECz54+a/2xhuCvOx53iAdNoiCBtKWkv7WX2sLzGdERXOtZe
nmkJaKWDUoMU0RtiHpXDHUUrGdR1FnGAdChmobwBKMVKrvy1gshPaFbKIiF60ix7
31DR3tkTnV0WPJ+AVHcXnOfLGEl5EG3yxaM96g+YWEkHs5T/366VG4luSg5Wc+VC
LJt1RyhsSbCjANfsvGpIF2bSfl9wc6Yb4G29iHXBs4lbzT7pku+E383O9yyfHLZ4
wVoquWEx/HEP3yFvNZQuoAq5MAhuorKVt7MihmlFSlZ//Ye8+X4Rb6kK2dEekk8K
j0kStCUNcConblds3Pn9SMXox4kcVRZjZcZQGLu/awq/bgjGDoTK+DvWAbx8k+dp
k2JvLcB3vpOSez1L2kWs2OU7D4lVxFadR4uT4hwVa+BKibq4KyYK0SSPHMnyuEvJ
NycMcIxHihcMLHkj3mwgIxseCzxdgmAtxIydmCealWt/yNuHoxG0Su07LgLHEZwQ
hqJg3axDZI35wi26oNR/Zgti8yGo7ZjojV8bq160O8iZ8OYcueuAqUw670Kh6TSw
dWA80BAIKwovinu8XSVYwFJEM3yRlMPd3tMP5/QgOTOBa2J9Mr9bOjngxt7z0aT6
wfXHRbLr6CDjNofmKuD3+JkBN4gz3qWJ1AJ8FHWRxSaaCaI3QA3LPRKmE2wOI8Yr
PRzT5aobfXsfKYoGBsutI3eO338T3Yyphky7JH+33JMcLuoJ4T1uZCzyF88Ts474
jslh11zZSlFy70/zYWj+qP36f1Nan+u2KnE6FKyLva1g0mnFf2MhUhP7SWBRTfTk
yCqBcw+s/r6tTgJvMTPjZZVjukF9v/O80FAAc25nz2FHX8jS5DSapH0EKca7yyKs
VFbMv91x7LXMPq62sRNX4wU/rdhF8eo3paQJWoRtDuhCzKVmcQezN4sKh6px7Q91
1Ip78VdaNwhqlSPEgA5Zcq3q5spKQzo6qaH8Wi1ij4cFF3AGqYyFaubcu9v8kkUi
8Aa/KudqFdTSCPHsFudJzIaZRcLHVnWqpRdkHU8nKKrVbX5G0PEEXEj+M4JwENe8
wculyK1eB0xY4meaYWf4iElBTD2r/5NlA4RPGcLkyJJIGbxiPr+FB8rBy2TylV7j
MS4yAdFIBq816tKeEYQejj5LSXFMk8RVFRojSVN1D7gtzBMvmdJmWouxN7L/2b1O
L+8GfTwmhUMhEyaBZQ9tNnW5Q91zyql78tjEKtGxRKobNB1uV7G29+11VdC2y0ya
7d3CyYsbMno2gg5A7jAulqAxQ5pinonXhkS7ws5uW3rqIfa2gIFprPEKpbsU7bxP
gN+L/7NVuIIkfaNk3ORuMyuM+5Lc2WQm3Dgrn54CHoqTVKvAVZgUJrBvWXtLZrKS
dBVNj+UzebryZBkKBMMM5GClbqn9tW/5iOi0jUvL9VdNCU4Wq5a8uJYlMnjZbAdu
dX0WS54F5DnLJVQh9hJqeQNIjvmkB7asgw5yM0AKhG2OuAF+01hLtxBom7JcDVzd
d3jxB9wjQ75joeVEB/pULJJ94BgKWMQgdEwp5L3yyWYqjD7XEkp5kIfZuk7Vv2Td
wqAQqzty6UUGBNPs40MwYjkrNRwWfMhlIYGX+akQr6lvxpxRN+4zhlbq7I/oZksz
WzEuVDh4x7dqceSegDB7Ixb6g7hwInju7BWs1+LPf0tf7r6C2BNdjbLjy1weBt0N
mTWE71q6jQ3wMgv46cpGRum7dZncDRqpWEYWMG2R7zgupSn56lwniyCaW1znl6Wn
HbHCYcYjQ5CFfwyFtE/Y7Fr+b5tb+284BTHQGW+xFunAvmCmGgrGIJJusL01V13v
/sP9rCJAGnYthyA6BUDUFQp824lP+cj73CFHq0olreMSyo/+1Yu+vxCfdkTGhcVr
7eG62KvJWbZZ0ZyGvkUZyd5/BpSRXHSR4sa4vlq80HXH4fVC0Gi5JdWDyVj8tJaD
078aqyUq83SDrJzxwrNgTL58R8rrD3b6qcTrIoph7Ezfaie4otZNNlrTXEFcjVb1
W6bbMgk6bZNLH4z2cKlfLGyY03FX9HBqmGkATd7kHSeq/n/vj65BW07b026BM/YH
qN4DpRNa5l7V+oRYQkBLR75ieDtLr0/MZqreohmtK8ZZtkNUJx38v/cSATQi+3Uv
3gKKCNx/d0LyN4NKIHVbxMV21Tg5u/+TGjZd6QLJ7TcBC3hxcg+6h/oF37TBo+e/
CRdLOfOoURfXzCsPULPYEl3Eu9ReUo11oD5AjnqQ+sHe5wf77SuAupnV7qBt9jI/
h6iLGoGMUNAKMxgVsJsCmBuSSVZ7uL5KhB75bRVjH8miBtjB7LnJVEbICk74qmhn
gzyybRrRk4gAMFLaEvqzOdIyWoTAOn+D3LRI/bVDyDMe/GxIRTZLLCFq/sfJ/F4w
fI8vybv/6xjc+l31EJ0/mN4elEqAsgj4jqsCTEltsphARDTxnmxVhNV4L0su1fRM
6vgigW2fyBamMac5VpoKB94jDo2R76rpAxweQuPwkEiIkPIY1wOzw+Ymn2PuTcWV
KUuWBMu5HXCm+G0proxafH2RrrQ2ZexJ2O2QmMomtW36AbA9os86WAgEORIz0AAz
avIiSPx4pg3HzF/h4pUikZ61Ty92rCJw0RTXjKL3zHnv2tdqZEXz2UTwK3FQkNZL
6MFV4SoAM4DL5jyqmTr2O7THBJXYIE4W6lFZqBb7hNRAm6j5F2np29MkWUWPXYXc
d7nl4DTiM1OnSZ3S2DBALyZCnsLqMWe0aAADdkWlqMn4nlZjKeZy3sdYH1n7OSFx
fsniPsGYgSTGSFz+rJgWOeoCL/mV4E6SkbBxN433w04vLSjlDYNH1U364tQHLg5Z
CwUg9Mj2lECoROQ/MG1mXjdw7muu7E1Lsd+/f6Iiqmqez7yvxBUDECFX7AGjtKtQ
pqHzEy/T37Vn6HmToOySZ5Ca3F2HTN+dp+HKjhUQMi5D8+e8vMrgfOqDvsqIhMcA
hZYsCdvWIWk62qmGRCgG21a2Ub7FAn4P+r2hq/JWb9AsothJRf6EffhH7KorntM3
XVMtJhNbwKU5ROURC1ipZBaKYoF7l2aKyCc7bqQtZ8VFXOz5sjan0Ly5f5IUP1gJ
R7yiB8EJx0wwdT1RvuTfWf1rRtSKma2EyAIOGphTJZrJst0AvJmAqeJH1eDj1sss
EN+mAjqZA0PTKxXVCBKqj3XUfab0y6A0nxds+f94uZvBtaKC6Xj5sFmzp3x5kLqW
+uuKqxBOlziwKGPPA6L8BOCVaW+jUJgGCTIf7rwv/mF1jHvrnWVMwTKKWD6cKOoz
/fjubpZCmOE5/YUSsnnwH/f38g3K0y3mxKJRRAFKmEQ37bhgrqFuAEv40TZhrACn
PGvdxVtNhnMzagCvM5qYsmqG2ppKqHdXfmpLJrAUUhBe2fdePbwuDJ4mD+rXjp98
OA6nKL5lJLWgCGXQQbrPYGtTlcKpML0qYaOIC6EtzVUszJOirDJK46cbsjkzAf1U
nslU0Uvoy0KQEXo3snALRSBpHjk3MqF+ymOXX/zPlEcZzRpJ8B9Jf4ziZMjmVJhF
flAgxtOLjOEAZqbRFgIqNIvb06wu5Q1AL7VZ/YrsDZ1ZBKMWe5ksqhpdUmCpdkk3
HwyUWsPomSpE8mjtnVfhLoKxIdyZ9jYcIqVML4FMNlcO7xT84PSodADcxFnXH4Mj
aU4xcloOZ4SHIVPk4C/HmvHGUo13Q1FRmNrwV5y0KiZeQZtulUoYS8y77f0o52aM
5cVwDHw+7qgFSDXHM0kEgAfPo12nfM/kjs1oGoHE68BnAl11b/nqh1rZpFG5cxAf
YL07jqmE9757Pt5KSE/H3yKqO/nkRC4Gy26o0zHbcoXhc9s6J0eGwV6yUUt3aCxI
JHKpYq2Bydf8y3g5lLsHMoIB6CcgChxWhVZn3gLA6IuIjBj3oJB5S+GSqY2cWJsx
JjDMdCP8Q5+TEHWudx4oVXkt8Yof0m7FYj64jbrsibZGbCC0Ux0tP/F0dLdspNYv
ZM/T/J5MkHEdkD91x1IjQH/mYOk2MMNyFiRnpmzM3k//bZMWMr24PIS5UV+AchXg
tjuzcvAWjAwxTkt/BfR4FlxYfAJ25qlx5PSft7onTKkqfqjz3I+9vDLkqlciWMz0
QblZ3AkdCT+KbO6U0Bxu8Nug2Kk08n52w2VUPPE68eBWzdW3LbaoVCC+3r4ycRQF
da0Tzj/sG9bCKLPoDMwyvcvBM0hMmJx8rKkfOGajrIhsDCcL8h2ztmf+xx9UJHDA
9t728Ugk22sYvfOFmulc+nfOFaHrZuFbtecc0B27wBBBFbiuAMcXIOx/l4CkOrhC
uDhoA02AJz62KLfS/539XxKK+Gq+iEauq+aU7SEPsJIUKjDBzDPxkckxtqENFRJd
tdTqKAxvSx1ssP3D5G7OEqh/2D4NSODjDUuT0j9N3s3ztI9cag49KYnk/8Fy/xAm
c7In8pi4v779nB3HhaUIhcrYqP/9ijwt0AnDTnsuxtiTlrfrxVpTWJYl5R8veLMP
GnxFtc3YwsMhEAq6CRuoOWnej+XTLzyauBRvRaP6+E8UAN88wkMAElnCbwb/hykT
8sG/P7A9EOfIFd8lL+odll0u9aBd3lxozREAc1oxKdS2eeuBwvz4l4IobL6+vDBe
glUIrjaIEs2I8gDhCeM3uNk46NMydOjkm577QZK96Mx3Pk6uudjn64diD0PQQ/+W
Y3ychnNqWRm09vNIOVyFbocusba6dJcudIS2KoCoboQpFmzkhinUmIOj9A3LuaaR
5dHsCZSNBd1yYsEQfh2SB/dHy0K9weBd3Jj9VIiOvC3tkAKxL4qZdc2xDMnE9Ncr
cwTyV+MnXcrrXIHoMmgyp0dHy6lYlZFT1NVb3Xzi8UzpDAe/+dOXGo4h6xwwAUn/
JrF39gfLQJvPFg5hzU4TTYr3ltclusEf6cfuPONyOkB3M6x1+IYicCMMXTEwqWUt
tKRhYn3Rl5xWtTcjf0gwZJNMZ3oL6xSP/xCXaLk2Tbve/Ho3D3GN213efudfsFzC
9OwFgCon2+lMHcu8KMUeLJ0bSe+dcza7xz57ZnCo85ZxeOBBjDERsFD+DmCIe+td
RJmRHAoc0S96co3UwffnT/sIzZnz1JxBthyukzJnmoQONDmOEp5gAdCXW7URK26O
QbQbQum6Yn9GNuIwl5tp43tQV5KAI0bJj7QTkHqEq0m5hyZpkTuAP2A3Qgvz9HCx
ttocYstrD4nInB2+WbE4n0F8pFOsYXsunA6647hgocKrW9jtLnvrlfiAwNUfZ0eO
rayJIip4ef1b0BsvI0rEUMkGbT9fMcH1/Jm8sxuaCME+KWhcvjPDV3mOueqClVW/
27dVuCCrwysaKIkpKVRusFJXQzPBi8kwoqtIZumEQV+GditEMiwnBuKc/gVH8GcP
gc/iWkWT5Qk7Qhf2SLRlek+QDdraVcqwVGT/Jnoh7TXd8WuK0GL3kr5x6ZlMTIEP
WQ0RqwJ4GTZV2GkRBo0G1SNl5dZiRjZpmS4MNDjr8XoHq7RJT6zf/OFXElDukxay
xCDRzFvjVdhcwPnRx5reG88uuBt+Lu/GrUChmUOVCotbBuVE/Pi+VVL1Lwc87Rp4
lazbFV5qx95PYVbol8cSMuUSDvdSyOEKFIbqwNJeqPnGvXlLmEzpeRmkkE68SSnT
P1Jn+4anGm1AEt4vfFa6ZCa+5vDJM8dCQCSZ/QUjeuVyAZLwkyYvy06fm2V4qTy4
UYVy7ruMMgXrISPKKW6iXKKnttdkQpH1ohO+N12g/u2cqt/U8zs1cUbk7ZMaQ2C3
fFHf9hGVPjEtfa2VVqI9HLwRmvwB7mKQzMpRtPmbLsNJ+Evvj7xj5N/Q6x7v2rQj
ThqaM1m3bnz4hkH9LEGcLX37ibZaAQy3P2eHukMrRfVGr8TGByjWEY6M1ZJi0Q9L
TyARWLZa0vqwPfVIogRlfQoEiE5xHeKeLmc3RY0eyEAkQSCgtsZBhcOcg5Z5uKwY
gbvM+QRiUTIhDQfLZdbGRvCOA4G7t7IMQChO27jYwZ5j9EMc4Jc0eg2XC9vj2XwH
zbASI9P/SN9BXj7Q35i0uIMz2SA0knV+3OL7F/4zYEaBMLmkLa3EpJ3PEf228kXK
R3jK05D4kDFt6SE4UCYx0zYYcWJBthMyczvdBdz1tW9be8UIGrpnwb8+cn0TANSx
HM1FS/z38BTGV7jjDhhiLvmY8jWCnUBIOmozg3TYY1utC2dTBA8ix7YRYzXU55Nx
Qf4fl3Srnj58BDiZoYBSoEPioCF995y1enFTC7B/Gh/5ABuUiZORHEfCS6TRlLcF
niCPRDJA0AFVytpt9+ze4cc403l8o7++4Kcv7xClRZlwxYDMGeImRcOOFkVPfgWo
vmnQdHtbRcOLcKHRT/vxY987i4ifEJ9OFgEsWQ+MwvbmaNh7miLasmLgYnL+mrS2
OIaBY3mCgWDp6Ib7UAEcyzKmBSiDnQenFy3sg6ZVRsTanZg0bST7rGMAXqkunt9G
BPePCVP6spq5ceKpJDdbGvP484N2zDSPW/QwJTtopAbqFHC3YVxeB7ubmCtLiXzM
12TE9GsnIRgOxTRXD2QRWBoqe/MqU/L2lB9eRyqp4o+R9QcFMcP3Xkqr1zilzJdw
00RKXy/OqyDiRMjEGtE2lp3JaOfNhoY+WOSLJmXZyHMcRoqLBf1a1Ld5ri1slQTg
sRLAaQ2kGWCNyixAQ6L5BDTKRJFTtHlQme+wvsM9dFGESMrHygUBfD711thvaTsB
2WZQvLIs3K/6AptBmoAC7HhwlFZ/Vw8+s8R0yF7URE4XJKku9EjBjuJGLaA56j1+
/Korv3Y3zexcMW2IRBHVCy78mT+gpn4rAcDPRs9uzufiZyRPPcoEvplKZCPqvVPN
u4llpEQM403xTXvaUR9aEbO8Q8A/+IQ0YgyBusXuaKy8KLPvzcsqJ42xQhg7nma6
UgWUgcGZ9SAn1mJuajfirMV+FEUTiMOGnQ35OSbItPDvxzwSU0xJpG+XKby3zDPk
ZlX3DvvUQb2+KtzMtfzN79RHGVjpV83ViE3NpTS7LGbLZ9B+yabNF/CBO6yqdOBa
uddGtE0yI2sj58bqFNay3Qmcd/3UPexGL8ac4zqzOk1RdqdLQ0RRBT7NVn+GtF/l
j1PfY7yUSPx+hzOK4syxndqjPARCWNOrf4d83DrjfF7QwH7HNLyIGG+XwMbLPVpz
4g4a4Ggsgh3vWkaNj+2ZDpmBie5IlmwTXp7P3r6JbMGRArqZZa1tcA8a3Fvu9VT5
A1Ue78sBBJpqUjwoc/jAwIcMJr1mH3edeflDue3Cr351NNA5A9ZLUpe7Te7YTazt
XlGwzPHtvJ5+eDvjYW5YCQAL8E04+1nsanszq72FaraLQTJCIWdwnKT76VN+8++Q
9brUqGfDrOcZ4NWIONNKLEXf9g9TCpANqNGJ6U39hG23swjJgM+D1SHlAQOEkPqn
MCtq+d51KUA81S3RWhej1t79JBUd/jzb8pcF6XPvO9ua9r2srJmrW/AKXxrO+YGk
c+7nsdkH9kbWY1ISmTJBHVjRTJELkqd1vUJR2psR7s3/OFO8NVkmJj47zi8CAyEn
EZzy8zC6ZCL5EyzwqGiG+1zEVY5S+RUfYAZHQMCQfeteLJV9TBLtxNfDnY6JZi3a
YUUYypAWQmTQbWYxvzvQKtpaVmDN4kpBDwUT/Z/3XUTKTXmcalnYv4WkvHxD4lG7
f3haPrk0EjoaVG2tMX25aF4cPNUiJfzZI0l6eckhXEaMj5rgsXJm+iIBvWjelel/
XklvS53AYO36DGdbztakm9PT9Bf+UlzK+1GrRVNEpiNO98Q9x+rtXLZhbRlGj2z4
XAIZS7o/gjXBhapNgAw0E+6XO5emjB5J6Cwh2eJ++gSrgYSM4Y81UE+wSr12PakD
c10XAOUqtd+VrccxllI2kxl3NKsni5kZIHVlTXfHHDzXN6A++QAFXhnaFT6MgWze
uRDzVlfHS2+RvSQwhBUjPTmJyH5qvlxQUHdjBaXeYS8fAFoGzcrMOMbFKZKSB7iv
IuAV6wjptlUkeSr+z/tdwtSO987K5uE/HSMBmWZi1Vs3McXwx5M2W74KuWXVjsAN
TzUKj7jm3g0qdgpZAUIMULn2nqyMrQZS94frIcpu68o3mL9dtNTc/KPdMLGpmQVw
XiFBmZHEC9a43Z0KPsBylEWch8lraAElKOGQvZcRsQ8A57Y7PaCV7N7mIpPr4AVF
UPD9xOB22Vq8WrCvN0EqZ9vCxtAFcVTsfPZGz1CXxOBkyMYS4AGoGjeoCZMlN9OK
iFuVU2Ifx1uFIagid0IrihwCQz4E/uF+oHoy3M9GNU9lVd66aHSk1LYxjxwWBBER
Mn3VPSQT301eelOtIdV+ZXBOaXSFu7dXizCirQjwjpD0ZObhDN18yrcbgNzynNpK
YSYVI3Cdub0szdNAZ/Qm+zh1vWFC68OTcbq86ns3IC0SqFQXgsL2CjMZ8gam0AXN
b7IlTe8buaL39l5pZZjqCPTMGLK3fM4UT4VDsHDPmPrixLPw6JIMCqAW6wyxKPsF
vq4fvvchUzUHZAvk1gFOCILy6859aVM1MrfmB34L3D4Qq8gPfMBuQFJOOTtDSpLJ
H7bkSKxoK3C1tEypzhTChOJqCrvdhJqChyYC5q6Qs6dBjOSeOFQNrqQfI2AIpX0C
RJgQKbUiNuHb86S56Wk6Ik56pY44Dd98EzWWb+9A5mFi0vtj6MKaVrtBuHKISTWi
CRNxqUlbAKzhQMWh2zSDrUc+Bo3ODo8x8DmqUT2hRzEpB6+WqJMC5+IEvF0OQ5nd
1wjqYEHLCi6gg+Gp9mbXt+wEqblRwiHRAQ1Zrr6DcXaUNBGgqIG84qd/QWW3i8YO
zsfhajdJhiMycfRd0Mo5GDLg+QuwxKu0THxwt+Mgig0BPiQOal8dzDizhiishaAo
bqsaWDJPVjhSur4lUO5Jw3sXeQto4DO6ntFWKlMnsitnGKqixldU1nSqpLUmlaws
38kEPm3GT2iv8rFPNqCkLkjE4XGi7MMeSve9LJ2dg9LmcBr0IipnhfI6P8VjRI5a
slYsT5M7OJw9xYr95/NTtEabIjEGWA8T/FPaGPqmWL0I0UTSNb6d11+YLia+0/sB
lKi7sN8l/PWNo2WvlI7JYhqRwWo0nOvulzy7Wj+21Wjq74/zVOJ2/tuzA46Nmm9k
ylJD3OLPnZRpkmWwGvaxOf5n3daoTMZSmlr6bBvFPQugme/Fo66GdpI93scJZ2zb
tbZ2kByWrzi9ePR8QSXVEln+C7mMr4uNo7cMa70HQyalGQfcvbyKFl0ocPF0vVrR
lcWjtJrQiOyUs+cBEVrS5NNSVO9/ljrAqgwrn6Z2zDNoOsRw0s1MQOijn56Ebac1
WdoVqJY04Ie1fQk5f/tlj6SQcNYyjpE6Bw92FyR/QsaYQiFeRRVEt/6p6PtNimBN
0yD5YThlG4fNA/Gco5Yd4um81v8TivszKwqCd2XrPsNq6Zb7x6C9M8qhgLq6lhT/
zqOrFw2NTNwgfoI5/ufB8sDSaprMfYLFJLFq2aQRyg1JA9DGHxWOT3/CPB6C1vd1
bBK42VcyY4gSkzzHv3x3+C0ybA8B5Yar64jpIRBhYwxUkJATdEZwGQ4BQXW/J8Fz
6yqrIMSRCRlPcsdYokyIbuthPFYlEGJUd9XHUgo+tbgsLbJ4VClsSyOUe2rYcwBW
1iS9D+LFCTqcCyWF5jqZ0891k3UbJLoItKFyPgPO10zgtZzBx9WbKYpQxJ4DCWPw
3fPE6zHvU4Yf3q59N11ggXtVntYVXQ8U84Ilcukck/rHdudAyvm+sWY3JRQGVQxa
Q+/+waea5lbVtdCrLV4Cq8DEPdxHpwMXd2IljThbswxm5EY5CtSTWMfEC8JByeiV
MS05QbqXEmhue+MyBavWfhOWekepXEo+7QdLN8KVIEPSEt3QJ8oLm9Kpiqtu8rZ8
tJjnELvhLt/V1bESoED8afSXCvOuGqdQckKwngGFoASVP0FW52WZM0ngcQzAWJJ0
IIZkfRZyjjgHcT/awZdX9hmVq18/EZbmyXAsDljknGsZwV4MzyfsTC69nYbjt8Sv
Dpj6ob3Nlzx5KkT6F0GQO6odNqXt4D+W88yc3InTxSvRyzqHvVvNvBS1amXMwylS
5KooKGwzCTwG0750cySj3eKXGxN70rp/UDbG/+nhc5g8zn1N2AARaqjFTfuDarJI
9DipB/SMx7k8hrWjDlmWxVYIVhydfUmfgi3VGJfQncZI3r5pAMSA7ifFjq8ASN5b
KhreE3CJUljO8kL7ipwqUrFBBVE/9zkyw+urVsISrBndxBaPa14bZ+6OY+UNeT2W
Qo/2+GlDDyeQ+IBfBES1DRSWSS/XIOuaWeIU9IzUuA6M/GHq5KtIViqNdCCfYmbb
51XdEaxZuGOfPK7uJVAmjhhFCJjZ2hhtq0pEZhOnAilU7EUvJbpFYJDfVh+75qD1
7blSEvHF9NGMP7w8Kn64GonSWK8bw60jbe0yLGgRfVS1nIBwBfy65isCKKMMNWrB
8GxTBruwp84YZpg9NX7zNYW3znbUuziNnbJe2zQR7Qs/IM8s5GUbCeEUj72tMOYF
4lX3cUzGQEUqVhBUcDf+8NFIEf7bQxcBjkGeC6/TYbvBXLA9eN1VaHfvnDg+PRgC
skJBcxvtA50JWwzqm+GTyHx/32iGU6yZOkZEstTu2ORITUmwRk/VM40wr2F1lB5C
35GD6pQ9B2gA09cRdNUdAcDTubh4ZrTMx2xtM/zNazcQDx6Ey7gZO/sMe8wxL9jV
HY+pltOMdCb5nYixxpNbGjwWPlZT0Hb41Cg8Iscoqf3KxxafILiJWUCYKUxcGVj+
nylc/70axGWDlaNfnkWlTPDmHgrgwi5b8ruadtEFElNxALCH6SJZgUWgs6/+yiey
poPQS/fawSEzT63zRRZhhEcaip7jAiYijL5p99lvhHC+ph9Y7xq4s9zq/QtPK3T1
R5lKD8G00NOSTYIlOY/Tyq60uBQiuzYLcVstUOX372b3Qjim+bWOjXR0hfKfhdWX
QAVuWomKU9HKrYJfVjzOBFOAjGvvRLWzyE3YGkOnnEHuy+VJABYIJtyVs1zLKJix
LCAliTIBzBBpy2vqiiImvZm/A/uz5EMMAlQ+RT+C+AkSKHuCe87Mis5Wv4D8DzEy
M650we3OP3KajOiEKHsfaf+lPZfKOxFVkkG5OzObkUOVddS9emgUmMg31RBZL0Pj
coH/RmYX+sul6a5Dq3jSJUlDrxjOXdxOiXveyOO0NTdRkxO9CtJMbXukMapa9qDw
8oPZ8d/DNIkxHbwu91NnjotHOE9TvxpDla/BXUsIkeXMf51DXgZemfiykUFu7SwN
b6CMRZCIkRCv3ebzBiqa+l/IiLdm5ptM6djrFfegTslniP7MaxRrWTrbLFU4M7xX
J5sVBz1rI11s97cls088Ni8TcOkPhDRQ91h+847t08LwB6cFy8k97GYMQzAhu3Y8
pGum/r5Rg5ETfKIYmHTAg81WsyFOGpQZiHeIVQ8rdIN3GTwdEMp+ZYtJ0fsywamw
b1IL0WzFaaefcCeks7eXOOu1tfD+2fqtGJ1fO7dWf467ZZsjM8Jz5tujvTvQUCZS
HNcmNOk1FW0FwcdWrh9MGr6oEkHZK2OaboFA+W3/GufPDcOuYpeESajnSIAoeHFm
ZJeAoN/aSm/U/8SeXuNSQrAn+kHm/Uq2sm0nzobzuBUB0G680GeAHUfX/3JD8BtF
7iopzB2XD/46zFX4sapks8RlkSKG3xfcFJUGvXuGJqKP7KyVn1xxXgjEyH0R6jKT
Ui0NItGQDjUaNApGpPU8mQBhgfjOd8C8vP+90AyawtS4Z4k0JBd+5ul069JHeC50
nRP4ZmY+mwU9pWSRdPEO/D0xGt7YAO0O1owzMuIt6lbFj3guLLMmorPIX8GpWle/
8nnfg9NHbuMlG4y20tjIE3f0sTvEh34vprxiKucJQ91x21ErysH2yomiIjUQmKXO
IGcLiVK4PmtVSr4FQhjfr5GECn/QDrQ4CfHlP2qnQTfqcgRGhfviNxi0u6qZ4s8v
uSKmQZ6ZuoZgF8Mq4i1RfRkkl21cwqmPO44+nhXlB+/bYmRwphm34h2LVkR3xRZu
Q9g/ig/5ljGsxvPBjz4umy+2VUuH5R4AThFLJB9ROmUbuuqb/WrQaheEaaDUB19k
HD+MrPCKCYlQu26Qov1Nbdksf9EtuLon2lfCCS8fBd2hS0BNdiYSIDnfPvnkIqee
0yddqavTnPlWxIV8bQbDV8YbmUjifyCFRbuAPDs1L/dwt3WvB/LWpakuRJhlyYvx
GCMfoaVIE7Jsz5Pbuw9xzMIBvXBwrAewkRQDodsPGtYe//7CCKEjBSeA6u8spKhp
wd345bJyZFAQ2u2wVECGlxbDa7BIQNdWC/fucbQjonR21iYHX/Has2byZenxJzNJ
ocYOvQj89zcQuD9VdXDmUeqcN/ZN4p1OvsX1wpAMHd7zQSpotKiUNg9adL8Sn0P9
DNmowwTmnS0rSH6NyIT2RDClXa5+mkhub+iBJGRMLyeBhPBQ5K3VsZ+HqAaP+CkI
Xr3u5eCxMUc/7XcyUGChnhQLgkw1v04gWkvvBD41o1thz9N1vnICBABy8qeTuAaG
yOkluI/t3IwAevZQpgkyhEsq9neqR0yZu02yEEDKDhEvtuyS50D5+lGnTB7FAwSC
TuvTdD/meWe5rjNyNtz8oPUO3LdE8ecEVka/1GoLUWRfHHAGAX6Ej+bFUHBSA8bb
uWLP+IqfLUzLOJgEOzeUK/MwF8DCvdoL4IjVof4mQQD/hpnLj3EG76kvjCZXnBRu
HtD3eSeZ2RM38KWRtBoTUgmgHqNd2hSKUoos3mymUjzeZFhrURvWD7ZBvA3InVyn
eQSmOM0qvqwXIW5gzmZylZSK1X4HnUf/T92MbFkjIgmedUbcPuAwgndR0yryzaOh
QftBs/dSZQTruTguizs+3dBH2opQtbt+h2aBdpCfwZGqaBnMPhd+wNWNXfgMO5sO
iF/UKuAk6Kh9c+tRCiPbs8AY9gEMtZKWbMIYzFSZpYCyujpNRcA8mAb/LfVHgY/S
BLpNbY5F+p45ZtRU0L+9RcNUwjgBdFam6nVFTUncmaYmbDKKtVwmTw0fJ0/rUzJg
+LRcXAoL/nBOh0ZHS81ogZjrM5ebIxgPsKDFM4RgieP2xDNWWiw0LBn4BaBKMUA4
WKCJ+zaSeY9n5uXNDz9iH3WCjLuo35cwkcucQxDbXAgZXn0sk0IBLuuE2BdtlV9F
wCPdmFg5XGjjVuIachibjvUMjSJASzDD26tTl+uTCvibYs6Qcz9SIL2kn0aha4/Q
pv927kT3bx3mCqu1Gp8U65V0K4jkgeOR3YcQvIC9a9uxuXnZwYCEZg1zE6/ekd3W
VMRIC+7Xwabqcp4azMFniIn+PAEzVpzCsi94tlCm0jvnr2OBS+LLyukATZfICinD
1O3oJAIbKoVyYhEC1KEfn4b4WGxhZSIT0cy6w3KpXSlT4MO777QHBLCrlfzrmKFI
rL+OTML6HYgdrNHZY8J0qXmHoB3c48xR6AagWBHrsJFGzbYzhp4wcrJbWYS2pKLs
v2UZbJdx1TQDrVp64GyJP2akv3On2GjsG8Vt/QFbvGxABBcdAEQTCrcOULVsEvj2
2SPtBbH9jZqfo2FcUn6YCSxJWoJsQ3E4MTsnGYMfXEmZ/pjYUDSXAED0Wzufz9wn
I4b3iXHVeBS0XPFG3dRhM0yV6hlcz9VagyBkf+KCoZuMWuMek/YXVS3Cr5HLf7m7
1FbCYGKXJ8wpsnfTtUbXhur3N4QDdgnV/zkIcQAR+htxHHWQ0ktRCfATo95Rozud
Ts8qlg3+rS+nDAkwp7gYM+luCpeve8LYMRhzGHTgXlR/0AsEpQApnks46RYM/s9e
6c9AePiao+myf52s8nEjVDHbSwSFAi+odqli949/kQM7HgsW93s7n2QMWjVPFF3x
zCJQje6KtgeBSkvkwbR8HMOu9lnIG8e9E8K5gEOHSKIv2xuKaYD+rQPG3OQE5oYQ
8lMR0cbV9CbjJde8LkIdNrK2MVO/Zfex9M/2xb6AYRvaETnR/POTD5WALmsXGm0r
nxCZfytg26fIKA7g0UEEFWgkfDPRw6lPiWIb8aL2jMiwrRyyBnJ1/ezYLvGFyuD2
WyNHjudHldr0sHhxCIETvUWyhqAE90jZfxlPm1V7gOSo/pJewa1Ki+MpvABcJawR
sUHJTLWGfL6sqJpqxB+CLqlN+U05LDjo+wj5IkQK/r6A6dnNjCfmcP8WUu3c6Wgh
1bGlUJ2dJDxj0McKrwADdAApLeqOLw9rEfuBz2izUN8sF5n3Dvu/WNjHB3vP7/rb
RDraDjznheQMcPtktwZFaelQ+jrFJ9Q7A1N0/tbuxBvzAIg1RcVvzboVIW6dLt8Y
+yWJX8Iq2ekL/AqKo/eWsNLWy/wx6nlOtHCQnUzT8rjd8rKYUuJT/l0fngI1c6Bc
5VLCNBGM8Eb8xlAH9omfiCnGvszIy9VTLyXWHlkTgtkEZcsNxqvety5eqj02XLiO
Km7oUOHkYuWQrTcXla3QbKGoNAHb8A7VEDPryH0NZps1QAoUoRLy4SGMOCfOPsGx
0l8nDFryjvGIQpji+aPyz9ifdqAW+Inwo1lcsOVCGPO84xS2d3hjM3Wcwl2ohuNM
WQEKt6u+xxRBvi7RSkQz4EH3n83YnXhQWMPMkR6BNtnLTL7l3YcnQaxhXAJoJF3A
qd0i+4c501I7aQMdgkl8mIIu8WfG3EeaGvmXVER2niA7os+1qF233Cyi0RCfjTCP
RelXWpHVpFokVznd/ZQZPNiaFq/yozeZtDplGKdRVn/i1NPKOhJEn88weOHUB7gm
ic1RyPqaKBvJFoe5c0VnO/3b/338osrtD8oUeViN73Fn0mFNtyaJUd+gWRCmQQP4
KCPWhlm7mX2AY5ZkPXofeYeuIgSMQd8+wtU12RJessHRScNnwTYcVW9LZMNTSzha
1wz0Y2JGY9XBTpsaOhFyKN8EJkeLSIlDubS77o3aJesF7DAVj+DfmEcpCZCiUCxm
DZPViIVxoC9wj0xjG1MqDrelHpuySM3Cg1e+ncfufyONDuAftrKuBUMGwPl2Wcyp
odmN4W5agG2s4+6VDS4hCemLlVSYwuoKIQ4XGbQF5BVAuw016j6NLTSin4VdqL96
xpJHZ3/ESD30o34k0J9MdcOCCzeTNuDDoqN8FSet1GHPnZydhNaoC0b9ruMGPT6q
+sMzoMPbHzpYsDvuOWkIWcILqUpL0oRlzmw+g8KWRQweg3vgSvQF5K9H1pCcwWeW
Tils9O0o5Q5PQsHvk0aZhQFYxrGByKWOqEPNq9bkVGYCoot2p0El6vfmBtN8HjWk
4/+q5iG+zfqwlK2zKYxHz2aCjsBOH3qlmRpuLh2zVIj4LTzJ/OsZLx7KzTXAGxFQ
cD9vRcMflHJhN9ughR1Hv6Ta1dbQ3YwOj9Is3SBr6Jiheid6as32WSTOv+AIGTvK
PKNetvrbS91X9ZCJMMkP2SqAeeBXnyto9L2VFBfe7XP+9bwk6K/Hmxp/1FyPp2eZ
hp/dsGD71/tmxAMIlws93RWA7KHDsnDbYLWtj1T5Mx+NNdZy4NH3JH8kuvs6l4Zt
UyFmdTgIEIcLxNVeScf4YTL7Mr8mTaA2l+CE0tjkYbUKvTiBWy/4jT0/+gMg6L5o
43jmeqi13bqUtv0wPJWb6VtlRqi6vEN8vJ3nY8+B32DEKJGo5gQ3A3SrBDRSa/Zv
4A6yZypp8PoKdTo+XNL8cD3bGOR3PYn/QjeX/pNj6v3NjSecaKqamTZ1WNPH5CoK
g4yhm0p1f1Y6whWpx8PMT33oUMsuNfl1r7TiojkuJ5JWR5EXDQM52O6RmHyfthcy
xTMjfbjmaI7F4MecELmDDsn2cIv7P40uTSXDXkpRZnASi0AwREtjzVR1y7/1bXic
bKOR4Bnz2PFMCksVxTxRE42+qGhF61gJIehEdl/vsFHrbgEWoWeZR7w36B4I55ee
BBuK4CFEq74nsQDli+7ddvkUCVV6dM/kiyvIQQzFtKTnMtjKKxXfyGQoX1peqOlf
r22rZHxgXWnkJi/SoWQTMVXvzoqB/kqtXhFMSE6TB+P9XcJLrgIBYPidF0L4ZBDX
vds2IRatWgdC0BpMN+v97X41S/qwqxMLftq2Jzj6DpCDgJdr1WZP54kuLFMQGMMF
pn0wS+T0T6Fsym3H+ZXVeU2Hsxmg3z4C49iGFNncGobV7/EV0PHau6hnLPLg0ybq
Art1ED7bUCLoeQhIBt72+1+rphJJIVNpzjG9MViPlOktJQ/6u8DrYLFoJOrRFpQn
rj6qu2QD+Uk/YLKiLd6XLIScb4v4qENTPqs/5EaxSb2on2OQurJMklelIngcUrQU
8V2PJWdO7Er+zydfZBj0zmqKw/NRpPi7k5Ky4pMElyANX46VO9DzUlup1Kn8F31L
EzCroZj/2cHWBTAigWvF1nuGEW3bUoxy493QxSFUsQwcFWsBNZwXJ1xF4q7R4+3Y
U24x7eURgEXtGRuxfSwpxgH5uvuDMdgqTO2UbMCsQ3P2KnjZ3AcqtaSqi4c6u2b8
D4IJKYbnjRj7DiHaNvlXQQU49VYwF8kSZa+6zzt5K0/7S/Et0cNkSYJwZqD8IdeY
eXIN3rHfdM9wX8veaiWxA15Z3ggP/xFJMZDM0ZsQWT9QNb8Bsc4c/l1OYPyyFT2z
+wAnWYRurJU4HHT3sFFV/Bwn2yIMCPuxQ17DO+qSPEPoe+zwaAznZ2PnDJSmqWhv
v7lGo01p0setVzGiRbO2m3tFWvdMRylEzoF1XyKN/l6XbSIfrgAHZ1AMie/UAO0L
FB7R+OIQBt+SNtHETmekmJiXqM4kgNodLjtSJBgqjo+/a0O/3BIVlBos0PA5esBm
eHfU0DgKSwNpNVf2AuK6sVtzf0wav381qWJqkBNpWKLYE7MsrIaNZ8W0PToyg3n2
BSXH0nYJ5qTViGQbPPWAR+NZyna37121aAkJXXutuxQHbGSFYe9XRh8KCYOJYa/I
zU1b6udZ6Q30gepGrI2+N4W63WzbXcG8xclue2ZW1Jx6OgWrbiHjYA5fdMsB3B3p
dgYBqUJ6/pzCa4OAHo5avYkUsI1BdBKlu9FTjsqF2dZ/DyEoVVOk9BcZ9E17emnr
ggWf5VrTnYERETV1R0mrmxp7vjI1Qt9x5smtO2aysPIeka2sUc0kbrCPe1WyPnyi
c0ldpzIrxJInoyTEjYT7XBBFdm4E/P/d+ALgCy4YPkvceqotWnV1U8RVWHHgkYvZ
n7Yajy8DV/TK2ZLYp3oNq1EzEYCYT2T9m+KfRHJ132WJ2jGH52ElHFvm+NWB1kHQ
wneKuOS4NCoXb1Zb4xTq9J0oKZBoftCDuSFpmAzwT9vzjkvBJA6i6uA5TE5paaGc
xNmbz0Id/rMxVqPrgNZuV0CYm808bqSOwLhpNqiAqu90LRtTsOM/K5mrZV5sTvuU
yDPwfQw6b64Q4U4fyjJVq+nQJ1DIP7vDZ4NsoPqptbiz+4YFYZGFhVdwa1SYs7VB
WPuCXsxk4RtlQia292fpIAVS7TPPugbbN9J8TJ7hIs2/NNtoqTsAFYynCRTurpAi
mexoVJoYkQgpNSIfRz6YWPedIajteY2enUPdII6xQWX+0mTpsUBbNEqHuN2WLrLC
xZJ8ry3xYClbSgRGj8BB/YCnPkL3mBGoWoahUKAXzm6PkQYRj9K+MxQLgjJZNnHc
Eh0pPxMdb7+lSX37HexmSt9K/LCQA5NMzDGrK9zbf6sVi5JiBEFMgQs8/Hr/Yp2t
BQR0xqBtaQm+7EfVWhIl7294+dT7pedQZ7ea+HoQrcOaxNi1tx+V5CEYn/ZYsiHp
TzDGWY4gBWxpwT4YvOInlNHZhtY3hgWso2tSeGXykpL7thm8KJAsoXaJGFkbKVuT
yQoZx13wahqgUE1sP/rruO8/o7nqUtRMadLBoixjWCBeCH9G7YqskD5r85w9HzmE
PCy9mdp+uzJ5RjKiAgfI6KlM/VMvsM1EHlR1+2ydAyGJK/76PfL0LtkZx/FMhtvT
nYKJKtSoLXS6nnFX5IfUAX2y5YhAxThC1Dj2kYoBiCztAZzhBwzbFLSKcHe7S7oy
+v2fyzFJL2RX9PTlqgNbzv2G2a8YXxQJpCdOV2ri0a9gGc2WHSWPTTSQc4o0lm6x
shzeIFWd6Njr52t9Toy3NEdQTJF1JzFxqtrWp8Vx5trfbx8hTwLuqwcMA8l+pH85
uZxEaOwu3h0UcoeTZCV1w5F94kC8hhPGmTIqTD5mGlwTfFAt65cqYWMEOZvB555m
AxH7d7Bq2lp1dGjA6VlIZCb55LMWc+23yyjPF3wAYgc64vhPYyqsewJyZhx3d09A
4GTh9gP70Lr7KE8vXHpHwBDCAvcGV2sqUEGJ5p89tz1vy57Q+U1F8SnfS8qvIlGU
1Ekuz5eZ3Bur3R94MYKI2LO6aNYhAlEZV1gsWCelFwnPosH53urd36VywpRfHA8L
mvG/LJ7rHfVG124iF7QVQYHh+vy3e45GSPtBto/81ib8phcX7xe6QGcwyhdOHKdw
bDongn0tOK8fWx/Rb0FKdM8crJR4RNP8xVFpdWtbrF8zZdnZp7Gkcii/u/CCHcFr
UcH5MCAZyFe+Nu/dQXbLWxIYnYfT8bKVWha4s1QnqJQgRbCb31oiTkB25S8AUH1V
dL+eV7NF9adntHAn1mKb/JjdxysFiv6vqNqXQbunCUYz0i6mFc1OGBHtRf/QEHCy
/4t/eZE4TGeYgfLenE7ZO0ZUFwW61N5klmgg7ADA/mOrO979re/29JXEsa3LACTn
8wdajhPbXad4O/wfMmUGqXPgvlIAZEjouAtDOfr/WvSb4/ghKua8yytZHwCuNmPk
PyC0yIM44uGEBIwfQmw2a6N0264bOVI9vuVoiBVOZeW3TEJNonExPIVXTJy8FgL/
DXw9qcEoPJFwkt28fQZQLMJGmsBR/ZcoFMs7ol+NXUx1cHbPS/L7Fmmtce/+MrCO
0zj3gjH5wQIlYK9yb3Kp+Xkti/iuU14UKyL+UMcSMRK8Aabc0kXXjP7QmbRnIlhe
WZkvBZqggNfW94D1llS98ICCxWnzjMhgpD3QypSfBli06/o2bJ3Ay9APZvQfUEWQ
qnlVON+2A1cx6uWezTKiobOrLBU7zDgs+PZwHBEKdTkLd9yilH3D8Lis/TdcHtVK
0bmZhAThcpCf5seotpNnCT8hv28NqnrJywg1RcSOTYK9UnD0yAYMI1VwPwUEjCRp
1w+05MhiCjTnJRaFjcDkgUq/u2Fk8jEclL/jlAgp4nID8QdnTgrw5AlsA15MMOxx
amvmV6J28tBHBUDt2BX1Hhju1TSxYkm4Gn/sfedvz2//NYtM16UgdbRuog3Hz9/T
lxmRwVYF74CFeCjJlN6yKkMKOGyCfR4GxlN67tHwWslpkd1Th47yDcLecy47rAyc
yxbtFnXCkpZZGJJ8zGPqr38mudapg2oY+Txw/R2K/IVQ3Ra1131HydRArm6gDCzl
duD84euXEdC1wMmTEnGFOMjA889efc6XhYTrZKCAE9M/xWIzZxhaz5ODsxGshzr5
po7KnhLlhj+YBdJQ3DcF75GyrT2wb7UEOvrbVuXd7IbH9Pck2IhoUrYuyFySzN2p
kRoYE6LKKLRwQamZZ7J+yxdQGgn1AuiKHdAIAwrjX4hiy5hI8EPJfLPnhKVF6K80
eJOQba6u4e6SswaLHb7odwPlyNIUjwwF7YpM/I3cg+rPecHxe7NTemUTVDhMQnWG
R3hnkbYxw1ZgV6Q8CYNfApgaewBxAJvlRW6rdgRF4eaLgnJEhq0atKybCbEhzDwZ
HlvsTYpH83Vz14Q4qblDPpZddysi8Jm349jz/J10YNP1hXlYEyA+vzQtoaHAUpgt
gRhzgYU7NxqyhxY++JkSPQonjvPWHKm+wO2ivcaB2qEOTeKgFlNBeui7Chv74Ntj
CSudGrkLVF7aQMEClrInKDpXPPWZS/rWvjLI9PKdLji2WZxJLq7U1WE5HVCQFsIF
iWCu9eTYGdokRy0DPmBSAL6b9QbtLOQl/DglCO5QYAToDfrYYbQlWNKSkxfuuESI
S1c1F9ZDA8NWseVTv3FTPIvAot7Zy5kv1lBECxKhfX10d0eg8bszLlb+ErgyfIoC
J8n8EXiXoyq4jn0ObkJRT2hDMpQ1nmSATmSWq8z3BHYJIBIrSlYLFGRkJqTuQs7j
9wLV1eCOvN3cvadZ9rwgwab/8wuhr+QLXoBs8tsL/GDal0LD9LxBZSPPdPM9U+Al
wZXbPcJSsPA9oKNO2nCra6+yM6TXTEjIcXZlbl4tz283Ok6msSl0Kt7Rg7jRf98i
lJldq/z/jcl0qXCm0b10/LMvKHmth+WeceMzQspONQCgeGTRoCpRWG3VptXoEKZN
qDXKyhxZmviD6ik2fBZll753rpzLrRrs7mQGYrJLrMD5Bf1X8cRknPljt1RkJ0Tc
hptgCNmYuW4XKJ5IRAMH9naVa9+ZDo5c4JZm4P5xTJUSttgdmzDHsbySg10st1wa
DPzaeOVMYAU9UqgzupaLlDf+Sw67nDg94x+i+JTK8qKO7i2YCuz85k56Oq/oEjN4
5uCE2AFLizQ6AtgTiyR5YqGtbq7upSQMpNR1wI34c5PfHhJn1oek0CN8h48KkxDX
yZtQzjFpw4J4IKtQTOKAExQ9/OGOlBN3HGwhinJhmAGPltS9W6k4iv1N9o+YnjF4
LYeNnEm1m9rpxFSW2w77wLu1cvmnOCACb3TFEKJH+EzlkHI/hChwpvuuSyRjIhOS
9eI/vU25jI+aLmzTMrVVD4ZWhO2bJ8s76VV2tabSyJ5uomtg03fxWGMJBY5tSAT0
sMVM/+qqYpn5I3iqBoC2gHmcp15Xg/edordf2n6QXjHdMtxyxDcva/K8e1HaFnra
eYTtJ5cEUg30M1ksLBX4Q29pEZq2cRwWMFBjUYxAcwxfdgvDhzPn0BOnO5ZA2SZ8
wQ6Fp5oB73PdnutM87u6wx4j9AcssYS0bE/6tkzc5pk/2rv3p7or/a6u0GVDvL0f
S7USqKbkC0e683L4zh2S+N4H7EFAGyLWBXh6a7J3FNi47WzwrIWjpg4C3/jO7Jo4
0g1ubfbExbVi9iHt8ddy5w9tgqqOFy65nCQYQVlhXn6Tg5eBj1Bp0jaIrtTL8iOI
Wet94q9V7EgCXOkH3iuDchnrIAMF2qkY7ZccSp+W+accEAosD6f6MwV70T+pkBgK
hs6ArmewSCf71OvRcJ3oNA+W0PL9wWNosXvDzq6NVLBPHpAFnCMapF8AbMITuV/O
n07iHxHREm7dmIpAlW6gG87fjfRuqfhCG9S/zvH3q2t+1GczfoUhO8qBDFo8FfUu
ouNAPMhp49olixcaqR5LX0Z4tA/pDk5NOFddJxZU0iG0jMcwITxa7gRKIsYOUwfd
xAgaavSS8yyk6Hex4qcvoSVPhJRK10Ovra1gZbgHymvkAVVPCNJ8PM4ol0f5lvir
YLiGoaWb4WwGVp/qqheKT2zHWktS4za2Mg1OsKX+WlmUw+roOiEuoCm4oNIJqXLP
rzsHn/0pACAWagg20ey46yq8n4p0UjKyrpQvys1mcAeBu4nLqKd64mOJ43upm2Yj
rGr10dN8pdbnm+OQaIT4SJ0g7cjT5yR5zsttFud7O8LebuG3qODNNt93eZsr974s
zR5ftu39SW0bBCrAoPupbmcMNmKCgdiH+S4t9EULq/BS/FvTAJdpqEcNNXzTCB+Q
LrE3wGkA6dbilC/B2Y4LhQYmqHPrGtu6p919D4p/hYg7sWl5/20s+PghGYTPyp8L
yQHyAgk7gIbcYIjTvbG//vQ/X9OQhmiRjzX1c9r+pLQECQp1dOZJDrPLqOfl4cye
XxdJQIU/YyKN20/7XJM4F7hnRhRG8elLZ4QcLvYJmhWP9Z0pOC31hVIThpGjnqEN
zNQg2D1ITxzebMEybX4RAuoUKrKSpDwAtSAAm6jvPoBJ1Pr8JC9TdDKcWQQ6kMOn
DjEjFQvBR1YHevRFECw8UsfD3Prm/yBxF+0sedR6tWRvFuV6+dShVP7EUagPOX6U
4luXPHnrh0O0IMcSQqJCO5z2DYVctdepQKj2gTz9JUb/IB2WKA3GKvktbtawjB99
qYiiqW6qKnUUvIfMYzwJmZjz2UE/fVYnh9CP1bQx1DJZjurNuyauHXa4QHlglITp
ksmKIemaSVapFwYPAloLGboz2254eox6MWJuZjd4hVh7qCK7tcJ5Ktn22dpcz7jU
MBDgd9CniB2fB6AppEf0Nd/+Gi2LwBU5hdbCfhFr0Rnx2bN/2Oif3C07B2kG59r/
SqWjcrMJbObY3EbjHNZFMTIHQLRI9qNwv5QqtrfR3jkdklFlmhGPndDdpjZGyKXC
VpqoSZryWhArWvDpDtbsZ+Oda4OAmc8sNOPCAGBiE7silTohxSjdnkHR/bU7ZxpP
+ORtuEaxggpf1QMyjuPN2l5E4Eyf6svPHJO0BMm6GHCdHawfZMtQyIG+aRHGvArr
zRemWCnBpSloRtluax6lXpsTEy6aIW4ZzyBT/QK8AYfAPAUo2rWl+5C0l4F8vo60
RZwMdGu2OJqh2lj4EC0CkgNKBbKwAS9wD7RbMDmfhB9qCSQKMj+Ty9eYIOfOhIjf
16BtQneBP/MzJzEgt2eK7yph9A+Drl2Fw/NjjZ/QnbUT0C+znngsy1Tv6m8CGYby
36S+/FJfNfHVszuAruI37XCcy3z9VLF8jZkQSvLhVhLHoiSB8/MwoNha182uOaIt
7rL0NkJP0La+mpjLr4jAeQ4xeiCxiYT3xE1CGcs1OYEyIAHu3jf3i7uAgkFtBx0r
VhdK5Gu4kwITR3QyW6QEFt2b0hUQR0mW0hia/GSzKEftOgxDBKYCoJhU6tJDKGaZ
rtS9tjEfBuQCy8LYx9Nlm7WZSKU+3JCXh6RPWHQcSf5D+GigiKreoVHJuzy2b0BJ
jB8+8QU6Xf9LSGfru1Ggj/0DBCe7mBQNmSHf8+FDlFEh50ohe8/enTpdH6Bg5hXY
2cHS9F5ZLANx+fzucgcUb05r0MeTnyV8qtbWgvwJK46Gnoa0Ox1cnlayAFGyZQ/3
7l23M/StUcVDqfMJOPKbzRCfbT6ccdJ0qrkv+uSH4jtQuWOvoVl/LOqvr6Rz6Qnx
X6Aost9cRfjtdRNdCKt3bCEVMCRCSWD0SBomaX9BRoYLTL8n+eNvsriKeB+KpKbY
R59L7+3D5zgTEF1cAtBBF2x1LXttTWk9gbZRbQvCYjNJzIybEk7VJxKIP0/DkEOP
uGCTGNa9OFKCiB8ZO4og/Eb82nSu4QybXLPFMa+gZqbVNzv6jBWmp5BVBMSJMDUf
H+pJSm3n0hiCviU8Q4XEcUwsicvkrvIzJO/xuPAzvNvEadimQjKsaLRnZMGKRLJx
sdRa/Y+zB20Jn5Rc0aKPG4TJKb7dVzAp76Grw3sxsRkwkmyN2SC2xXJUopp7jxlU
muGdMfS10xuuYenLcmQrbSW9R/IQ2Lzhv4VIMRlod0mn5YbCbd2NzblORFF2+LGu
poewqciVZXkQQnxkigG9Z9lqI5Q177IkGa5YrSqm9YhdCCvdV8RcbB3/eCZRU4Pd
IId5OwNSQuuomTYlf9KPUvSE+jEAj2cpMJLvWzkm2fWfmGmkshpw+JhC4xM8e1Ww
1zsU0Bfu7YiboebFkauA2OsHtlSBgJSLnjjLKobrJgGbWnUs4voSd7WNdKtkXqEF
5hStBDXTD4r6qSaKdaHuXmSM1Ir9FIvfUr+WMhaDVcM7Ig9PH4J+mymrBHO3aI0/
uzSzO7uOsscSYSl9mz5K9nzJtZ3trL6awQCMp31z8SoNzL+CdXrQzuiP1FEJp7t/
A+mqJ/iUn3TP84a4d5WOMw9dh5HSIbwcqQ3ox2LTmmwQCPR69VeuyT9rEcZ4qvV5
v9Li4rxJEPeG3WukFvWlAbSNHkDYrPT1xyBnnXByor/Egqp9LfmPh4NHBfYWKV3t
ALXYIG7+0dAPjV+ofZC9dhGjNEjrF6WCRtGkqN+2d2OBLW1bvzavkjh3/cQzGgo3
N802T8F43tvA8Ab58vynpTVohdmEskpkno/7wAFSIs1wwDrmdsaoeyfsW2MJ7Quu
WHXByd3iTrmeDeG1TQTl50SdsSrKBt9c59pp5P154Hc+yVAet/tSvf3erwrsaFWR
NNuRx1Fb1DLdchVttv5ph03IEhyNhdua+6vtdIR+ilPUvQbOJPOvOXgyHRMcV5/H
Pbh1ApgShjcU4HGAswDietwib2sMASBmkfBKRP1opK/ECztmF8uibqJZ/GcwoFSU
C4aPl3A68nLWH/b4GEvArtICtIfaNA70P3hyvEpOolRMoT7ggCVeqFcj8H4D/dQ6
VR9I9t8naGgNqK6yzQ04Cg5vDCeLZdt2k4ba0+PGIEtI2p9mFPT7CeFltRiWRKoi
+3jRhquUzrkHowVAvFZW99adc3Nc29u+wc4BQxdsqu7QrSSsE2X1OWspmSxR1A/N
KvRH11eElKRr/LBx6YMQxk2pbiokgTr2mtdGwSv5ZLfrpasPC/ugCoI3zapfzLGB
oZXkt4AZQ6dFkm+d/NQ1I2P1MhW/gwCUDLXvdydpTRcM5oeB234VSb1qTXpuIj1K
Jd14DIx8azn95sHuPdaWFGGZBmUj39liEFdqPNoXeQkAr8kP+jvaMdsSvMQ84UA/
E51QQFZHl1GNaMld4S1s1uj5m3bg4szRsm4xja2qw7do4RydlWPlAja/HVu3322t
m2FssbAz0EqZS/9JdrEuOkbSvsVu7/VvX4/6HhOGbBkK/WDJ2h+yz0SSyYjJ42vH
yKXi+EpxA8xvrh7prHZ3OrIwy4p8OKkamTTpiRSTelvjqjYNMqpf5mG4xqC0lpG3
IjdMxFSaAwSKXE5x+vjrBc4NcBo4wgEBlWIv5WoebSlRIsAljNHJWYPFrQeGNz2v
fxMUAXrpDgi73ygDmxfAYJ3TidoN8kiWW8L4VkjLisnScz5sy3hVlh++n4euLMqr
ZwFenQAs53E51F8K0qlZgHCszXg9DMsvKUp2fgXqaGRcanknrx/X+KnkXzV/VilC
2GS+9rMnxETAQrvv5h7aSkMZWeRGiKuy/QO0Gm9AoBJUNcW6hnMdkDORVTGku6RP
N4P15RV9khJysK4+ZBTsEhC1STgUOz/4NeoJzo51FsH8zLtELwtPy7bJoZ5twhnw
KD/c/dkenW5mwcayoZ1Qhg8hs9Ut0VjAJG5mOYjRlTa4tu4pI92dKJU2f8Cq9svy
Wes6e61BPEDuQzSZgu16Vkt7Y9549YSxoBC0yvA869+AXeOYK6iRMhpEqgZWdJOU
vq/y51uDt4a9uhydDphX/L451Nr6APXewxG7ci1S2h9nwONR9dpchYQ2dB3KrWGk
AzuVOgEyk7tGGLOKvgbyVGbHdgQpHwK0HQl0Jxc4+Tbl21yM1/KEb4OyIDNSo7Nq
u7Ft7g79/urrNdf9iPYN+uNyYwF6ecxb1YdtgS//xAt6x7+OF6RhGwjNphKNsAHq
JpMA+JBkEtzNMC0d/H+N04y281ZRjDtVIUomjD3dF9Oi4g8a17/IbjI/1rDcKn3F
pmTTvto7bemtO42dAVt6xr1Q/oga5Hm0vvJPUSFs/uDAMYLyc6qCZSeaGSyrQ+Z4
+0QfPOJD611lfeQJlVLiVueusIyoN5eVJ0AF2NL3LwD7W1t9u27i2Umo+VMdW1gG
qnkPdrZlBH8aD08Bzg7/KJmwRwFyw5vsyoC0o/3s/bFousJ2RWimaacD/hNp8d+N
2aHHBhZlfPNznoxlvFGWgUJwWo1zqyMMzRmBZbxllH81GXzhi6kaVCDEhzea2578
o4vef8sa888MaM0UhEzQuLAO2OHZAMVC+3V5+h/y87mj+M9aFH0AsS16ZaFmTqYA
6D4jLut5mk3MFx4ftGMtF9d3uQjAAhsL00O3wHh95bvULU3suiGv0E0V12Xy8nPN
c568mJkQ7i26lMvXd2YtN2HcPHxvB9PCYxjLzq/NDT+7ylesvdnAfWxB78sJZM4Q
CQm+Lr5hVr+O5cXqGC++XlZICuOg57QSvudvuSZI7BNPKL78hcBQxS1VOdlJFUNT
X+Jj0UF2l9sSMADmrw/TT2lPlz4mRXzXXtezie1UGqu7zWYGXT/qtnR8CeWyh5jn
Wf6zjUIcLoJA/cN4LcosflhJ90mW0bOKsxBaaf5Is6QPe3LWbPNjyf3Oq4RwPAF3
G0nIYZseotHw6jB9/aiN4SRxNHyKaeWdDxWGK3hVQmoQpQE+QpIeyC4UzOJyrpTo
9llJnsPI20gO/zatLOLXCSx3/+2wVTbUFgobRqtAA9LYxZAeEdM3yGIJ4B1r1nf1
iR1hsdR4xjTbuwhn+CQTwPa1sILsySJbKaW8BFJbh9UiH1KspeF8IjXmmgqLc7kI
oRqbNWja/rZU2q/ZFSdYK3lvCYUA2pYgS23jEpcHPLqTyVa0KAC3CRtiBc404e2Z
NtC3nswR5aaGCzy3LbsKRlcTltMZo+q2nFsQvC6/gAIJGuckHtGjtQa5NY2asadK
lWJwkpWOtwxuG/qF7aHRshSV6BErBTaWLwGRcvvUe1gGSwQWejzWz7n38aGb4Le+
COt4bSkG9Gm+kmGk8oqIHa6SfdLW3SOJ2jW372eFlmzwVyb6lJY1TuPuS0+KZmyw
2hx+5Hj2owgLWd2JjYGlWmE36t3dSeRl7F/vwajHP9SNc790itBMDpuHlK79SbeW
z9e15vYJ7Fvko0TRice7sTFmhweYNvLcn+J4soqT/CidXukPVYOGoBdGydCfAS52
x9tczpzcoE9+3nEzUvYeKF8lST4k3/In8NH3XoAzLeIU6RI0Op7jVcdmCXQadtcp
gbBoCZRHd9I4iT1aO+rqxwKwP0DeYgMeeJGuSy4k24p2mSkGuRSC59fpa5crsgOX
G8UIZqmZOzn8ALZnElP1T1Yt4STSINV8UQb+Xj0yr4NFjuTIma/LTrIE0y/iviTX
qID69mWalsbp0ho2d1iDiD4FRUmUu8J9hWm2Av+327qjYq51dKgBOLsATQDvVbC1
hSD86de08VVoYZ6G8GCqcikzlIADuQ+tsxceHy41RlzhXUSXxQDHFZeC4ICvMo9J
EbABR/GsadWb6ujmmSvbdQRRIgBk++DqugWPWOZakOBB26BPC5qzdBJ7kRnVHiSZ
KVtBCMx7PRPFdGsFTaMrOLXqwZ0TBcB6w1OD30FL/u4l4J57QD//k/yMdKOBM/R2
YXUuJcL0mdYiWxzGQEQbc8HfqIX6mqlBFKtWqip4pUnmn3llFZSlQ++bNDtvukgy
pdIqI5kQKKXkYW7yyAvjMdTA8PqvB97dQBvGS8oJJ3INauqNUaMD29B33u85eErD
xCvCjn5lFQfdVlHpoG296We1uh0hUmzc4zzQZoM+4uks22ypxU+XXuFRRtrXQ3tw
rnDpp9LkeZnfJqF1BhiqbdH5HQ6mhKR0UPyZA4L6XcNHrjui/dtBDVsdM/sRUDGu
3yP2QlDpMXyfUoak1rOXvvMBT0t31XaGYJB9cYvF4nfpOq0tQy3rowF0NcS3pzrR
CUKXstocvbv4PNOUpuBZrdKhnb75BUemVKUWisPx/11JqgoEHlGrbToYgsEb1X3P
GT9T+j7wQW+LIIcQl1DtMcqvVgPeVFkQfmLeGueBGPkk3rPM/f8MJzMcJa7+9aOe
VBCYlcOYjM3Ng/GMHrVHswWPGUSMa4Taxj2PEfdvsFT+NxoQk4ZwvJn7gWy3PAhw
VD2WKqaClE4WGfZpMoUbbZNtrO64a1j7g3gG6fubS3ao45tIcHMhxBKIdjLQnZGs
yAK9pukPO8294JDsUwcRzMgv2jd8sHsyyFEi4HdcAQHH2OMQF73weVxRrQktOjPX
mIoRzL2M393+j0fDXduqW6ARbOj8QjNTcBlp1XVU/JfBtYegU+m3qwkLop2lmzTw
B20sN+iFiEM75oTR1JSl56B4tZGEZBNWS2F/BXsPk/s+Wp+wJ66keq/KT1O757P3
PduhgCI7Xl4hbU0maKHIKXonl82U1X2RmB+GAVkXKPEM0bZMXj4iMpnr1EhGeRrI
ppIZH7Wwl/eyGBTBXHETkYQKl88Nj3okLOkalh1FyLtXIJ8sgIGP2l/hndJnQf34
Z/KZ4XmpSoGxXtMLE4bsBhJ8lzoPpMxL1GFKslcv7NAMVRYXv0ZCFUO9Tv7Zht7B
fvEMHr+cv/xVcuvnp0zZbfWaEW3P7u9dHYwGmCmGvYvvRmdTAxueWvoxliFSpMir
qrvYWmXzA5jkWcCvQLSwsr28/YHTCMY1RuLWTbGXvCyeNKlCm9pLRHVqnk/kGO8D
cn1lPxnGKDadpYRs4KR6/DwEsd7USh+Pa+GUAHqR3rrJ1Gr8wbDZbAI4Sg9/1foc
kDUOhWKCfsINM2aqtJCWXimtzAGa7ydigCpH5MM0FXlL9Haz84VEEpdTicEQj56d
VjESIL/hjDqRk6urxmk8uSLlGwtMwMcNYtqyGgkR3+SJ9S6G5WPNYPEZEca+nc34
qqIK4fbjYc+1wCU/a85zuLjjwGROTmaNIZ1g6M79402cY3pYlB8ZQWZz9UIefZEh
VWmp/XWQ/7Pol7Wiyvn/kYLQuIJmgUKMg8mQX472EQU6nc3dzQupW+CFWgf942VD
U43hyWgA/fg2nx62y3h6uaq9ru2SNP/3y80VoeA5btazKPBflY1kQ7MLNWDb5scM
grWdfGm6OCiaTZmdV+jUQhMO+fEPbrkMVMnyaA4/b3CVncxJ6tqoQgkyEiAdlqIc
smQV9InKOyRMgJCfk5ezsTV7spT/IVrixmIXRiVld6h+DyLSyUihgXCo5bwgGSvd
ZqXcZ/AyKqO7IpwVXW0LugV0ABVkw+pIvBkn/diz/P6WIf+bUnqvdX6izRwUSG6J
euq1xvcFd8StjUiATdgwGtrry1rDBl7hxPfx0PaMPbnDpWHmwTtLwOuD4clJ4MbA
u05W3y8PWj0F5jZ+O8/CdyTtAhAuewPPBafw/8Kl7YMEV2o72nU09NifPnS4Pc7a
n3VRZUr67/HrQr758SgW+FOP5fHRXRnGupfNHWGiXIXjsz5JN+NQ3xPYFpf0DwZT
/SfefKklt3p+0Rz4Z9jGOmAom7EBEXZi6CGGHl3PkNsOAeOmVDmePv1fiIFo1nyF
oY9IznDvQSkIJAJ5r5dOwaKg+URVNpIulgCZTPMegtyDLrtH7paiSzQ1BaS2CdPm
yxIxERydhfO34ui+iXLnKdff8GlTLJlPs9CdUCtrD5Iiy45QZQTtSOXUtobUmLkL
T8MdMbOXV1WKIP6piU7m7g9fE4Gc+qRJ/ZTYdYYWVIFPzIoD015Mn7K5kE370Xjp
Pi5ZTfV7g1N3mXCoBZjOBa5pmzAEyHoJgHnBM7a6aNAS3177Qj+Yo3Q/r7cVAEZR
dSXzW6NCIh+oGQXRgojkiycZP5De2OPRTLXQ+Yv0Bj/reBJQFdlRUb43tHf7Wy7O
19qtUQ/Ri4MzF5esG5NL+wsxT7I0UrF4bdGSiyjF90uzsBGLYHG4jmDoa23O4Qcv
xuLe3c8L1IVXdGk3/szsfipVJnmeJlkGX56PffhrWt2/5ynUeT+6Lp9HzkQDMjbT
yGbU5z0tkQ5WKot5dGODLlvxHixzimUAFLUa4Hs3UO4EUh5JXTBlqQEKuLa01ZTc
hR+kHjqM3paRU7t+kyHdfx92pdKjGFEJ8OglIvLMkeVHgRionopss/480vJ+0CAu
ncHa69L0bWpqEwSZNIu7kxFKQgK/CBtQmHaJf04ll6tv7onUgyBrXZL/bpCHNqdB
Ip5g3hUhiZbBGcG+Kr0W8dROhOI1HFB09Ebk+tzxyGNwUXylxDOKsCtaUW6OmmyW
Xmfvj4dS2KZP2bltCswLAjEZL7GtFsu4D8qmojH/mUK5qYLluBHN0lYzZfIEvgfx
o91K1XZN43C+MVICsNenIUDgVlJTFx1mPDQhn1CPM9u9Syt7iJc9No2z2T7l/XN5
lmc3aSgn+zMyU4b3uIfAnnXogm0JrxoVr1eifLcnNGvUNyb6KoXztoSpOqw+8c7n
mfbj1A/oxNFj5d9v8TIuZaoCid2WtSKMdcVJoFPHfzq8QWf7BGfgm9dF1GqmP5jM
2vhGGQp2mpFDyo6p8PhPaGZVVN3lsvELIdIYUI0ZeAHWRdTOhk+9t4tHp+RNvAtx
HwSqsHxEl3QZtVag52A6GsbSSpsxPmEr3sV0nEAR65vV6iIcbi+qxPLpdcJ2FzQn
MQREOMxVJF0KFUI5X1OryyyFS5zweGhGrlM+jP79GxztVXm0WnoLZh116yuFSlhg
50+asbDNH16392lWxRMRorwHihZFl+wZ60sVYfQ4amxdpR1tWTEkpun6qSwfuSSi
vPeetnKVNxTuY8MVwJa2Pfc0SPG47D/m6ctb4PynQsaytV12G/xGZqAzBXKQ8DwD
xrctP6RtEoK8lxZUoyiH5/Qi9ni+Rwjxg28vHkZSo9bNEbre9ZXe/TTFLeEh/JVq
K1YRqoeNV81VwBgRwKL/7GkVYT1aKEzOaFq137mSn4+ujKiNxczy4eeqiqPVCETw
mbBcmoVju6zJXSnLZX71nVPD7rlOEwS9Z+u1bi3HzlYhhDJDWOwbWSFkS1irv+vE
pytk1dC1Wi40SaDZtZlwSuyFZSvNdyUFcr8t8mRNIvuRHJRCY8AD0apGeJt/XsW6
70TcfT80UX1ZyEe0tFeHmyWV67KuxLC1/Tld6bMyuDVuGOJ8svF6ijMIt23ghGjb
KoT6MF3hzeE912sbNRyaH2atxSfkYa5V+LqMqM/8gBQVu3PYAroB9hJADeQbJl89
V696XwLo3Zdrz1VquDit17PbimiJEL4oa7Fkwde+M2fNQHssWSee0DOeJZ5tih7f
VTp+yu3d25SB0+1jn0cjIlUwzw8fQhyO4KZntSODJOVEjwXlrdviTCUeOy9HVPe3
kqsKaUYD56+jDhdYZ85G5djWQjc7ewefVgCt14321YCCPuVbb06bjp/Ot20D4kAC
detCbNQbanJZyfmEr7V31kZ/0RhjJFoydXB0Cd4JnXTeyYVKhGwD/EMmDhtUBbpq
eBoNUtQijXo7ob8QeWeuOGf49l5XcV1waWWjTONWGhFMeg4Fh7/yn2w4dIOSq5Jo
T51N5VJqLj383sT/hk5zN9k9D2HdufZha3HitcWxmwlpove+DB7Oa60/jR3JkV3b
aUryZd2eJdhwbTfuMHxxZMk1sqF9T0l9ReDKjEEb5Ws8m+JO2+eGoda+lPy75uE7
xhFwz2VfFVlSTW/uM/K/GN+U8WlTZT9RDBqedKt7o0QaBVVTCja4gmyurFgaQmJi
JfJMkSaM59qyExhbrwXVCYFkCci2NxBB30zuppbUC1UevCFrjA4zNfUWKU7MMvOY
LJE47Qxk3JYJQm+NRp3EGVa0RQpVyQa1JcshpJhBxslxHY1NvVZn4ok3J2LL4xlw
bwH0ciHcUjnuaLqM0hqSmOtvSF6hzuo/1+mLY/99wDE/9gwE/lsCC0mmgBRN/RBE
oOv6egQnrWcevgCybJv93DJuSrDFCWjgIMTTMJTy4Qs3EDjb/bqljI7oZyj0kD4d
VOcN43Xz7A0Sjgmj050VDNvFtlzJs26PBJWYWCbQf89u8w2sWKWpOtJIwWuqpLyd
6jCs8qk2/77LkDeZd1wJRAGCMZNktAv8cGVknNZ7DDsxgJM3Lk36/8tr7Vhg0sd/
x+iuUdrFtvi2IehyMJciMZzKE1MysNfunOYUeI0oieVb8Rwz8ikBFc3/6IrBk9OW
KMjFS+1y8oE4pfm9ApzsPFW7xfohZMcxqPO/6VmpJY27wmGvOAJiOvyHHqjT1ox0
G6zft8ESugTJQywHrVofAuOF7TFzKYr48PKwP2ndOMe9bMwAs4J9gZ0IqXWQpkQG
A0TSkhe+A/+Xhk59GglwiPWQitCkHLdP6OKSbNA6yACeRJA8097a4D/OTtD0pAYI
E7pgIRjpUtaKa/SQhh0HdCEwPHzWYvV4OlNbrHMnycMJABb9Wyk9E4txeqWHxkNC
AnGuOxCsOenap2jJXQW6bR9soautLlzupZo+8EybcDv2TJxBvzH/dQ+cNkxzN8tp
TdRE8UE8AMQJCqVVOe7KXP9NvIadqZQE49j0YHg5OrHnwJrf0wwxbnPa1h5ktuUV
YhXXcin4/1BcbIeBtyO8H8mtQZYyl+GJTwKIcr7KgqQeGu6rkwUA0GyiO/a+DC9O
tZplShI5lLv9IsbHTR6NoHzgsz9XTISCr20WLM2mJoet3p8v12fMzqYl+9+Kzsfy
rKQOGHB0sKsw65UPTPz2qJW3bnyV+z1vC/lU9jzUFJf805yLTdfV95AnzuYdaHFQ
o+2GDCOUH0AKv++ptS3P6VwejE1/BEXLfheGZqUYGEQWJotIuT8LvqtFwWaFIJBr
ZUM9EyMPIAnWPviTSH5GLa5n9mMp/khPsxxhrw3zkeJ7W+KO2a7cL0lAjsE72I/5
sOR0Vf7MPCD/yvWWV9mswIasSQyIKeZYpzx60ABsR+eUYby2Kwk9IUQ4Nm3fmlNi
96UCIRL1OERpyWIJp9As3ltiXjN0cYpasR6WwSoOuIA+5eeOJHdmXYYH1cmbUAan
8UxyfBEt15XUbZSKQNx1bdZ+L0zhmrZsYTQ3rlbx/DbUe62W9Stb4gyIzCOC60N0
ocLgWRUXbQXeidkN9agmzr6HXOG/H5k8OqJ6g/vUO+y9lrk9NYw85AB0QnHM2n0Y
crpnvvieiRU3N6WCMlVYb2giyto8OyMy+yg5peRVoumzvxAAgUFNQXCWy3rTXAKb
+EZ/I/1I/WoGIHi2YNawsZHSlcF1yfH9jXxh0gBPjtISNDJ416W6brfXTgP63FES
uCcBHUTTywCTzmb8sZifjsEu9cDZur5dn6qi9VNY/LFXQJJgaY2Kmc+d4sJ6tm4g
JzRmVxpxnarS/YKjHVFb4tnf92exYoTtI32NOdIiHRGChF7FaWtWE/DiHb/VdZI/
E4cwCiVm2dyZw0FTLwWzc5VK5CR8sKcFD2o2RmHeEJrTKEHK8ARUR9/wPgfG4Ogn
CRnjZmBJFNQY/Gvx03bhfSHllCqkoR2o+7U62o1/r88Dk7l0mlvOMVnsIiItkPOo
BD4JkapcnPgUv6SsTW7WhM4QHACHs6flmkcorj2mWyKtkrNyve//1GlWJ6eZqPxL
EQ03dXVlaRSzb6Kf7Qy0Zq1mPGklnGNS0LTesanFwjupeZAqofp57E6Dyl0plUcx
n6TbZz69Z9bFQNl6auqJAeTlI6FRuss0qHrJoNeoA/goDuChpJ8P81RWQHc+msRZ
UXBXkBrUQSEAPMesT/m71Z7eHtad9o7TiJUlVCynyQx8urCGf6ZNk8XovzpnK8Hv
XpkURYGvdxQ9g89fkacKef1RXdYHdPRUgMABLUwyEJji+TWydSouTw1O5agwGM8a
3qWj7Dk8MSR5U/HyMfKTNcmc5IpcbY4vDPPd1qStenwWz0neluPEghKtyZNdqm3c
g9L8vAAafRM6P89usjeF0G2DpGhLQxL1TthWUB09g6m6o9O3l4c+/pP1yyXNJY4E
+6Z664gLzB1MXirjUZG0ELsfbL9oKaTN5lL6Bk1H9kSy738f66kARA0H4HHYns4X
HO3kmAmYEvCkMq2pOjRaykDwZ/99ugteUaZ+vtuBgMbvhDDluM4GZmWWve2t0WeZ
YaQP9g3MdO5J+5kp1IfUSM5/hBb7RJB33+FRpA4zCmOGB6EbkQUVND6n9VdAjCej
43LIiIvo6Dw5MVkx9XVjslGNO75jMNlHneuLRV8KqNHfsRZdgGXdX0PYgosrJC58
hYWSIeIcnKw5SLF9jvD8nbkDwPvbr1x9LH7e5Ey2wjj06xEZOrtZZDDNah4oQ1yz
mmBt4kyYgj3Bo8M0pl4OblftWvB99A5j9+YZT4+bDkW82X5jRT99Qn1rv/0CyOHe
Q894BCP7j7bvg6g4CtKlbIf9W5B5B1zVK9thnSZR/PjzOSQTE0+OsRP0Ujk6q/3g
jJoQpiGtYFUQ5/Bitlglub6xF9VDXUBjUZu7X4Sndmov/YaUEFB1vKPndVP3igKr
ZSnD23o1Z88LvQi0Qt3lh6RNQd1JoyTKP4LNujQlosznW7VSTgxE13IVWCsNqOy6
H4EKhLMZTjRsb8ElvHk+cJEqpnQ9TQPyh9Uk5lTFA8m8Kfl8pkgUfZ+lJrfAlVg6
32cqlnVnsIQONrtOHsiK1xhulIo5AFUxyhwvxlvl6zXQPpnc4GeMwHUZc3TObJyc
2k64gIvUq6DnMBTHWig236XngpiVIgh3ShaD0aJaB0NzsOqaC6PGUFpdYpCbwPH5
hIjX7CZyS8LYQ/r5VBEwfXbWioN7nLkOfcCp5AV6+JzId6DWn2Ekz63hAfFT8vrZ
LTHcas1oCU3aitkB/WD6wbpr9y2y+49jx3AeI7AQgd697QoTT1CKoCe4ObWExmi5
YVpCW/tcP4ZSRBB7+h2BDy/DoL09n88PmzMvkWXDq0kDJExlE3ClRg+4Js2vnfFW
hFy8dtce0ZTSjGnkBKaBM+fGRXk/nUGkxIUCcpThFkj9czZ9FTW1PVsEZiQytWJT
jbqbGZzvdiMl4OTi/lASu3GmerseUopePCxaXF4wkIRBgnixVzPJf5V7hMEGCuv8
lsHqBcb8/71TlXfpUoOE5MGB5q93TwL5Wq1k5jtdnttpPaSbquYo040VAwnaQq7e
y3/W59gs6sibnbwIRZq4RjwT3KaD2Qe4Q0SqlKuajD0z9njq0r9B4bd71G99bo+V
CxA4syc6dyL5zJB8ZSEIEmTnsA6AMjfrulsq9Y5NP31euF49OcIrubIvFZWMZ1+R
gmu9d8vGHrmKUAbB/txz4Yj8a2ZOi6pPXcBhA3KkiaCVD/mfSnrCfoYQCk4DhG0k
cKsZ5Oc5OATkOOSTClB65pv4LFXyF9RXOO4wAoUGEXLbLUkcPyvRGzjsAZQB43DJ
p2yQ7sszVUMJH5wJT+wmhcnyM4BV0zkhYIQOyd81E/M+zQMZ9cv0TSsORSNYuf+X
7Lev6HGde9lSFsLgoF0aNTAZKq4mbYYEGHlCxZgLZpggy4qIsBH/Hs1ZATWlqIPh
y9d8nepfJ869GAvDj1Llw6kcLIFpEKJQcxjJLCxwoOAR2vnEO6HgTEvDpSnqK2p5
0+TCHboIT+dYOp2PxQE5jKH6aFVfD1Jmm3FmIcd7NNvBR9JtaCBVo+ckMJP6YxjN
rGR03U+A30pNsxNKWCwH5a7J9iL6ytQ1sT5eArbOUGUGFMVlbD+h0O7VUTVnsoFy
TyIxRzj+vC50waMOncFB+YB9oIkSjYuM9LbIFlMg8Ur2vOJhaxLnj2TDe3OU9kTj
tztiKtk193XZStWolMBcuHAER3vXkUmAmVc9xMg3Y61wFPn+m0HKsJapuMZ9Fq06
Fjh9Z0AybVLyyzFfbcbgg+hAavygj7mkQ2MehETumiec5No7WdoBPuY2AtSwDl+A
+QBgxge/ZRz/hudYiFxVFv+D+25CAbpjq8zSrCx0YwmJSQvzut83HkexcUsu/asH
ZzbBn/qDvs7DFxvuvBYP3cl5hoobScIb6YXx3T+kbBystNk2CX3v7e7y8XloCt6c
8+fDQhbnAchEe5gxHJsVkWKPUIwwF7FCAgKFf5vMCzMnIFIkqXvSN8OpfpotQGot
bweqRO/hxKdOLPzxBWvIYKGEfMRdO2jFFiQkuS5lBjL8C09zdx1suBNPS8pHiE7G
mEXUMZEXYWtazEV+szGl/zu/G6VbnqeNmFzaYsmsGxQNLqIMt0Dryy06u53Z4Szr
qVDnxnOrFG06AWWh+l5tzmwSNY2nkiSmV9KNjVGTnLnnuxCZlXMnhO/Ssex61KnZ
g1/2V0Ol8/DysRezJHUuqNIfmoZlH+VQ3S6Den79E11CAd1G76dg84cHk+phnzCR
oA/uzxzd4u54hEI1oxx1OkJWF2e5tl78ruhUHrwe+TD+B3iR5bv4PWoLdrGKPcFt
PTNEQGfmzdELOanI9/2lo5tEvBzp7eTzgOgoyL/c1B72ZxLvSQ6kMlZuYfWgvcfD
Z+lmfdj59CqHZ33dVy8+ymHKIKQRDyKo3nxmrUcOPW78Ty6+ZTijB9p83TslchO2
y/rxxM94CxHF/zrEaUvKZZiVxzuTaX22HV/OkZLwl4ph6dTVguSJIZ/UEI8pVqw6
5PgYN2VK97jc9QevOAI57P5TjhosEaH68GSPNMjiTtBU4ZGb/dOhf3D5AWzYJ83A
dGN13wxPaEShGscSUsb/z4TmQOBSHLl5BmGcK4/YjjWTXaYHVPkc5cxc6XweobIe
q/Ia6ToJwjoWVskMpDoqJCP11GLotR8nfgVsUPgna1qJIOEOmklOClXJjLMFInlY
nGMv/5XYEuLqTAZFYqvBBiO+B4Ok5pwqhAhL1yWsYnfgwydIyhL3IR6wtVzVUjKW
z9Nf84l50XXtHlr4NFLWMWI9s5AgXEPZSf+yg90AQhGzfWtdZZXkdnL1PAbYbQm4
qddU1UmLReR7UfGu3KGz1uBr619CUNv/B9de6koumuz6qE2HNGexV8ohOKwOqH2t
3nGnaanLlwYM0uaCasFJvdKICqXRdHI4p1EcN3shRct2lXaw4q2oF+obD/KC7gEp
PJzCxQxOHoXBfDsCmflEEpsgbGdeO8jkQ+LkwDgYTQlOWhJ4p/LbDpJ+F2wAanaE
dynm1EnaLER+D/3I7ZkRkmzC5KAr0hqw23hcUsYp7ImvSxpbFfeTy1HDOtOGY7q2
JyElba8I8zH0lbwUq+9eGqVTHE8h4erDPvIeXXpK0Tg03M4ELFpfIZGkMHVKUToP
ZIeGwn8U4QkqCZpLriUt7TakI7r2ZM7zt9iavbVuVWGTzAJTyOd4z2aHKyOs8Op6
7HhxnmJOPpXxn8pn37+22Qka+qotUNFa2Dgnnm+RYZKDW/hnGdavX+cKa0nX9aUR
tf0iPjIuT2GrZleeFaekb3o57gDVkQps/az8oFr0j77OvsvKMH7C/5cDxU1THJEQ
c8X8aS+Olo4UMOw3xDfuDNKqe4VdIjIsJSJMYHjk65HqIMCZVlzB2g3opKApHRJ3
hgVjnET5+m9lTBCjVJok5XFEFjcNvKfz7lucuksoVn1UuBG97RgEdqBOeyzuTRqM
dJRQ/g/OFNH4BGt2p8Rue4ZnKteqBemIHmrCDe3xXhbVemk+L5W1VfeGo/Xduh20
eus9Aju9/r4zNnjtCNnd9JKe0HCcISbUK13/pjxJhGRwLzbY7J6N8TMDmm0aaEs8
x+I8eQSmULmjvTz3oiACnuHmTXYRXkmKf6J6t8eSpRE8cfqFfqzrHLH2uZmMloBt
c7OBxamBskc6ImXuYEJNmJLy4RM1qWVoKHd8wnuXiuWi9K0fJGFa6XXlW0zKnKU4
tMIyA257iCLiOZ4YVlepZ2fv58WhDIsJaSUFq58sg0DxlK7wfRtZ5qFs7lbDDP8l
QexdbgrO89RtZkJzduccvQVDQjiw/l25ah693rWQ7onlGM/DXn04HDiFsLUGK5FH
zLk5JF4jNYBBPwfI6bJ1gtP8mNqU2GoW0fj4J4iWBzhKVcBG6w2BvKKqQNJpHnmB
ISpngo0gio7EG4pSHSUTDE4CnZMXz8QKxF1AQUf6bLRBjB/uCdGiXUW4rL0BaV6G
A4cqJTuOoNk6GlP2Y/PUl/Reh8VsvQU3856MzrTLrgAOQ53+F16cOc9Ro+DIzeZQ
kTuhc0FGnIewTuKIzvyzk71pee7sY5EervBoEUwz9g8TS8d8egtir7MwFs9mrm0Q
uvonI98j7NB4PXfScjO417S7Mc1SxA/QNsHOgau9fJ5JDC8lb4iXLWrez2WDdZks
qSxAryVmQ44KLQzPm8GKq05dVzuaRoKQrq0WflRief0yrIiwoHZQbBljfEY03qAn
Xjc/Y+QKXXHq/T82Uz7oGQeT89VfG+W3GjN4P4dpV6EezZq3JNZh76whYeuCOlRo
Z6AQgS6bb+1lb0+rbnBGud3qYmlPm4tOXQg0MmjVeLwaMZvTqS1GkRRCI+Z6H1ib
rapIsBln6vAqgqH3TeYVvRzO3IBc9iaGdlQ8hEkmlL4lLteJidk3HTx5amdcvSgC
H9fJumU91pFPh4bwxlmTWOqyLoT66daCJ5aDApzbZc3A3XySHkQ7tjoW/Mi7IeXS
A2tR8PIhW9lBjthwPC3LuhYue+WDmB6ppk8/rPfSDvIukX4atxdC7jRfnz5DBtxC
Dr3TE2+igeiz9KlVuL+Ng0sHQM8I0iM3+Bp3+moCHnKtTmMobpSCE838oYB1Mynf
4Cz4tgzQRJmI0DlKY+ieWPAIWYsI66DKUb28ISGSobBms0fW050xpMEDdX5misma
h2in6HM/DB9mLvJg9SnEm4ALqAZ/Sk4PBev+I+5PFMtiXu9a4DWgh4di80GqkWdc
T1peYZW7UwF3CDyC+Osj50n9w5d3ThH39Jld2rJ7ZN092Jm5FTDzyRi6ZZ5JExw0
lai9J7ALuryYzhpDfrQOL07mxIGh0L12B40gOWWpkvzrzPhsss9d/+jZi19Oq3PX
1mlGM09v28mv9eqsVIChT/9miziZm7724XosRsV+1MBZNzDiH/5Tc7a3HRxGw3+l
87npcowvmISTUTOzyPRjjQ+JAsIuNGfQmKTYCRpqhiHSGD+ja8Mk43Af6USbjzoL
osPakVJ4o3QqtbryWjN8Fw/n234mJmpQLxAzBteloKTnmnORvmdP7t13tmmgCmwC
srqzS8CAjtkOmJUsxttMTUPigom0l4ILtKwze5b5+DwgYoBBYcB2dwNjYRn58IEa
9sBBE2tWtdUA37zdoit/S1G+zU6gEzjHLGnG1DMM8uJcby/8zCQaWr/mdK0yMrmk
NjWqSQyi6+AV9FQyYX9CTLQCL6lbH16QvBmCrUEOWbPGxbTnsUUz5NTlhqfYi3hw
jyVHCLO5xlbCQ9VQ3aC8B4lWNjaL6U1udWiMskn08YiJjyfxWA7wUyLHuCMN1xDg
zZ7nWAEWqhb77fqRLz00RZwMNTGfySjlI9FV+bZsID1cXRXmSpgGlSVJuJXzvEa3
Hti23L3+UPkbA8nBmd8HucNY49PHLFv3vIR9TsPSHtJ/5ZNcgtZCzqdXRA4gTD9l
2sXl4muqElCRKB+9HPhMaZIAJuajbtmAXh6zjcaKq7QQVg7V+mbhXHP/7vTa07LJ
/X3zspCqyJT1ppN+Re/cSIOw2kn3MfeLb54Zi8f3g+lBCDKMNnQf41RqXN9Up4Zn
OEVWZyZEUr/TLQCIENVWqALNlv+jtHxss4FT5Q0zmQTr9GC1NCmZxmYvHKRbJ+6W
SOw/WnwioPSo6PtP2Thwb8DbHmjqCnBQtP1Djb/MKXw9vaWAjLNuEA2REU1VwesS
XWFu5+nypxropWfT0zcWiv9iX3OxcROZFK5oVzx+QR5hz8qv08StpBowzbCTB73C
Q+XBDrqabi6QrM2YmFTDvo5HzWGqDyR0nQXNixc+eyXgngDXbbutFkUBvuBlz7sK
1rxv3RbwYyMrte9GjVhRp8xOkbMhWm5eWj7ImtyWGp7kgevVMsn9U6iBgOnqw5CI
k6n97ckbZDRAcu2/mTjC1ycX8sftgEH/usaS+DMp79BxAAaT1/TMjXV4Mfv/EqhF
SVgKHAY3DbJgQa0al3PUKg55Uos9KAyEXZq7ec2WL860ZECo2otF8Kd8p4drmctS
tzswTgklXroBAlk/9eNQNkPU258XKMuPtgxUCxBUY517cD03WJE0f7mtZ5XAzhld
LNZoqZ6KERhWOLtJ+SRhkU64lH2xm9WEfm2BynKjcOZZKR7MwEF4JI44xxenCrsj
IImSCcOPSp0UQnOSZWTcIbDdvvtXTdTp52+gd5vc/MeJrNSE+HahFper04xIyNHz
Y4UaV3I7qYTgglwjZQZuoGBHLbqsNvTasb2evdqV6OhNJLqFtjDE2SE1k/kRcFUM
cSLzzN6VggmpOCMnIL6m3VuDd6QlwOA+2wQ2DpJ2ltTyK7jEhInnqL9i0k4VIJj1
Iqeoj+E7hTk9SDHna7/BlSgvNwN5tPIEuJebhbeGIIZ/hTYnRiBeIzT39Jm0nDV2
sJ+ySHWhMwXwp4IssHxQ1lEKiene4P7Vh+SuAaoK50IkLLSsEvkV9Z7uUyiQqS8C
/Gmw+S3Abyt8lwF1BitDNKBOya2/qIvAb1CvFe2l/+cJyx8Ajj8PLQ7k6KboMtv6
5mrOT3bJCvLWLYKgTpimPFK3hAfi2hzBHHK37S5drKAZk6lvw3nG3ruaG8vNZASJ
41hYbDiEHbRSQMB/aroTaewzBEsllkE0zbXiJGbfDIB8zQ7rksj8beqRJ+3JXAIW
+gsuvFcxE2E/IGteJYYfczrqr2hIk7ZCBVUo1MPk+gpPtxUwzetvYhEx9Zw4Xyi2
I+HO9wylkHmc2aAX76XuUPFQ+gj0kXkjIt40UGcmyAeFU1grAohjmJHBcOcEkLK2
9imTOVQRhK38PqbbwSj0bavnZsQfYKSzx6wbaiTRrTu/M30x5knMGgjCCIxnk2JN
YYQtLgPh3h5P6+SYsc3t2X7g8N1up6W2vALhOQUKVho7cWEsbG27Jz+/7CGNqqp1
tXv5zWaog1mLjdzFcalbAmA5GqrwdYe1uxQdlHu3whA0Nnetp/wZalZgjnJAz6u4
2+MXdIe/pcYMCF4erAQfELU59E9HP34j3wpFEiKqlrpvRbFKslbl999M4qqwVT3d
YwJg0JlRq4qdR5/CfgaWCzXjXdIaSDCHDW9yIg+CcJUSXz+BDkTS8SFkYK7ldfiB
IB5jP4HlCSluWiGjcjyLtsn8uZ0d8xsNZLrodexBqn4520uxLbjukup/VnAPhKMX
dCw1eVpMDClChzuVn67U0Tb4i8MFX828ePKSKmMIe7k2ZPJhMkVRy7X4r+Rht6Gc
QPThkaGy0vmMJBcXU/5W1B26NeQu619Optq/TY6cWoIdJDHosURGNIEgjQUxYBSK
E4Fcg9Ste5Si+dJ0n5P1n/Y4GhHPvkt4K2/e2bKFr9TPCM3eRxfer+fhglqq9Onw
jUqqw099bB3zbRj2ICF/kxt3ZWMZlcVL7/Tec/VIeLTfx8OQVaCNXW6q41Yt6k+h
iKVmxhd7cEqZxq7taBspdHztnqaNowdGoDyybwCgJi5v0X0pFREsOHm6TYO53phz
n5m020clUXoUEK0PfU5dRDqZPKMVOkk+4hyb33H7JFOjTfhZNPIFkDz0qykSNvGK
6UQFN7QfAZagRqrJrfAjPp+t9sbzKGVUn7DE7VbRdoVyKnT8p2IncrUXFbp5bzsZ
D/TdrOYSHwT0kDk98tFA0k5LmPmCb/u6OOqt3fgMb9L4MF1RfqtHIJDazAwAZGb8
0iLwutYQpmxDcdWHFm98XZNeRSAY2KUmm+n/BMDlg1bEHdLNg6/OaqApggyAZV3e
3fdKhZfPJChi2926sjdc8YoYykYLRmNZISd3Tfq3t2fdBIxB2SFhSnKnYPfW17Hw
hA4nXwnww8sce6IVy3n3Gf/sw82OcS21KVP4nWPJ52tWqKE1L3ObQ6j4DE6tMO6o
zhZ/0rR4fe3e6vy52O3FgsOJb9MUPDqIIX6if9UTsNsinoY7olyJBvPVDfPtQPLo
jyIXU5tadsBm/CZ+s7GPG9+SpvVhRbZJvnYxlSmRTAvx1mNS3xFunFLO/GauDufH
iOSccj2lBUjscWIvZ0M+7S5miAiC8tvfY2Y6aXUPrIV6ovZ0s3O6D/lBsjgCXJ2U
BUCbuicHEX7xvkyBL2kJFpKLBuusPTRST8cNPCKzt/bqkLEr1EwnahIjPLZYtVmN
uR4pGI402rZ+0p0mIvAbEp9Ykq3Uekxj9No4F0iUeyVZ26Di8UnO8wKbRHMoYU15
kNugUHpukUZrJYMn5DEJEqGv83dylLxa8meSeKCWtLwAKG1j2Qtu7jFfMaGEDsDb
gQwh7K2bBsI4mMGQsmKWbCEt9cAkgEtBOyLvdby1bEXf7VJF/mFF7gnrlwaugk//
zmUI+Fs0q4TP3yx+o7jUk5bW8xg8QEM/zP7BDFsCgtp4VYlM7r4pbopxskmFrVZb
fHVDU5HdpemF2ndioc6ek2njZt8hbRANSIeGZDdaJ2dMlSMC8Ou2jixjOuJFj4wv
AJBRYh5KjJGFcDU+7be0WiExQXgF/oFaEtxgmYTg/kbNOxHWOCp0Fxu+QIzroQLY
KpVF1CffYhkDoe021hgtUK1Aco5+JFWAC8ZJovstdenLtwp03d5MeJP76gNskmM6
n88eghX/5/rBQK3ei09wDlGot1JRfrMgG/IueOTL5XIg87pEuKEEMcI+gM7mrIfm
YSWDEDN3Z0qmUEmZs39HbRw2UCAlMLR6uDkyEkEwiYhOqnp0Qnf4+jUwdnjpt4U6
1ZWpTRAymeWjFIzA5iD1SJ9MninFVAue2aobyKNZv6RVmYsYiVCWIxDyDilSHo+m
CaiHSA/18jDf/H1OZTTJUD1rNZAEtwhUSTd/ArAIdlS+cfJPeM2ZcD59VKkTHqAX
KZEZI22OOO8qvNYVhY+pZxrUyQu6o6u/ZarwtE4treOuPYJdSdhS+axhv/bpeOv4
2Ng26AEjUUZ8BvSTP+ZYRUrmxb0mWCLGYBA6Sp6vhqWf4zjGWZCeyTWimSbNwVqa
JpPEYhlMwSeyoP6Fx15JfPjXpCvK+DxdHguB/LHRR44hRNUce3mjuNQrmwaQYKiA
eEPYESeXMLH2FaeIVx2u34vXGHpRkyLinda9iRJQC+HNh9dBhvosA02txAdmB32j
U+e6lHwfOovqsf8M9AMjkSpOIgiaaTWpQrKRJDT7bjPTXiNZyYRqUvP2e6yPSL3d
v4ynNHygem5510fJykYVlovcREILyBWBJxeCeTHU5fNRanOuZ6ycY7C6+pyQ6c/D
kaRSKgLKcgfQZpn/wtH9pl3/24H6YTy5+ApchnzImcF0sToV7Y3otQN0RuvKKTil
7EWgHBk597JaQoxl0iM1ZJ9ZZJSrdMXvAql4VOc2S6tmp80i7Obd7dIvWli/eEz/
zXLAScrVI68YD+BLjItqUsDGzmjTelarp9rih0Cle2njYRy/ZyhzfyOlKZ46ALHr
ynWkCt+r4We7Yh2dSycepaiaZGGQuB9OhFKJVdekthwndtiJtLicdxXChM6w2wQ8
jGVubiMTT6XSmqqn1XEVX38+r8Jn5pe0DUyA+z1Zk+gIOyHITc6iPieB8wB1yYID
Xj+sioB915HhJehTsJnfOvfaOzvvupv9UfgpEgy2wxyXqEG4mAsLED/L+KzeSRYA
EcgPKVKwbX7c8G2wDch3z3+ix1QOCimzkbR4rh11/VmglOvIfj8TeMUgW4uexXo/
yAsP1qaakYdWBIapZxZj1ncIz5yURDJbTPQBk7G7YRVScW3S/AuPaIn5ib8fPvbn
VCb0e7ybafwiTYK5ogpG0uYRM8w6SXhi3gYJOEGripGucUbbBRIx52IPD0V7sNTu
HfSUOozu0bcQdnDP88XlCT/RYqurNukgPoN90YBH1WmSx54MgaOwor5R72uzVzNi
PYNT3re46AYmYGyh/Sfp00/7nuPRoxQKcl7KNb8PBSHe/K/CAVyLozKNWcbOhzJW
jwlWeqcINFGF3RxHejX8sASy8y2LblaQBi8TN5k3z+RQadWZytbUns2KZE4/xfXy
v5jV59icofEhEoler+NEmWdymRaqTVEqD5B++mg3hJzOyzq7fqiJV5Hu64Y3nMls
ZTj8jjxr5/07y0qY9s561M4/ahbbo3c5woKl8msqrOQM7+W9wq4RkNYnQIktdfVy
zMqhjq0aIzJ+oF0a5EMfgv3digEsif7OuBVeUcZhXf9q5IlI4rW4tH6sx4ebJ+2L
mo6x/0LGFuGhg/aafvOW4CMkXUnptQG9YSBHhktjt7PuNDMGb/hik0sbVMwgYWVD
/LE2TEhVTti/9+3zHvmCvXJSk6otztf+tuQfh07nqGS4MubtlP+CF2gCBuUF8DIh
C5HUx3RE7EtxWirTKH09UpJzcfUEdqILS4Jmbsoz0R7qQnbClG31J9+y0/CC1Vdh
xwSa0nFLPJR4nwLi3YDrZtsXPu/kKaRuhKOaKH9/CRHb2depBPEcXqHcfYmZQ4wq
h4dK52jLfOqaC1a2d42LVb7yG3nG8Hme7HM9nRoSbLf/+VpGNszUYgUcPlG+ljNZ
+lrCEsYEPNpovWT4GgL5oG3XHIxjvak9J5SHzknWogtSe9WETBl8jQoTSGUU3f7q
lMoE96XKpeqwpOSqlucpm7/4y4aHbr+e9vwnJe3Z7CL9NKJaOuiuQi8XCnpnf09o
mhc3GuTF4W83EGb13BLrjApXv8hulvpMIrFtyg2Cw1YY/4xRWJRVE4XNhEwc3laS
/4EQXu2VyzvbZxSQf8iP6HHy8ayeL/zjyh7dT5QMUZhsmxzUUyVmPiM2QQHu5nkC
Xm0qYHQNsnlWgVyiotpa9bHv8KwmFrX/IzgHeSk/1aryr6fNFBgHFMQfaIfu7tmm
0/Gc4B5XS6kkiw+GslRrRwJDkV7f4YvO1fLJoq9r9sEAXVZTCjPgdYOAFSq0YFxO
o9iWZUoeXiF/D00fdU/gBWDxnlLfQ1xZx7v/QNzA9BpdEUSRuZuGfEedBVdc2FA0
UWZ9tgDKFoI0QpMS93dIjn/07J/ASVn95C9+YdMXeFZwdHjgRa5bkOZqL8fKpcYz
Ne78a5YYk23QFbbOsovpskVZuzFjlvW7kJRSdJDrfei8m16A4DZAckIw1K7RpGYF
3CkJGjn/canNYLKn14a+ol1pi0QJyt8P2RV00piI5OCmTq4fFK8LMmLMCHGZN+IK
biu5sJYdCpH6rmaV2LOGqb2bSzRtsuxPxcVpWXwOJBGc8LvWNeG5USpRjJ+6+Cel
73VVHbZZuWVEeXhyhIMrN2ksXR+rt9YW7riKsOvYcGduMQUUIeX+KajsQc7UnroJ
x41c34fA7vTcFWhcf+nDG8sNFPQ6qvR/N0ahYlwZX5DJReyL7CQ4F1wyPxMj78KR
yHk7aYu/ubvVJQCGSiECSe3L356k6c9mfaJH1lKJs/ckqKk//giol/y1dNLFr1cr
lFNYUCVIPyazPXEAuDpWa9tY2r60ogXMxqFPx7ubgnulIujFwNudUCo6iGs/wcsx
3FBr4gSO8MxRTKl+f5bpE4EOsPZfgKLAsxrAr/TqnznJQNedPhpqD360ebPeUdOO
JpJ3CnXyJswO3MW5drYDRYtMOlJvxOUW9pbdt/vq/1/6c919hQDikEwFKwN+RfQX
aKCWrYJqSgbjI6/NvNp10B97yRpQg2W4G/E/1ldvag1sZQGCepEyPEHcMJUCzka0
0R1HB1kBbNXN7mUoLkXQHubetjtthLauj0WKteLqBJDeuHOS1tRq4vx0zDRLLR2H
eWjNyqWQ6IuBYkq7w+5u9U1NG9iJVwhx7rwk/eN76cdRhYp1AA4YUsaSij3yATJy
hCbkkIrnxKAQs9Aeyrk40367YX4PS+e/7YlhpgjPoi3m/3WTjR3MIkqZBaGSJnv8
hgEM+DuMIvl0WbPH0NFRB1z1gwu+LGWz8H3o6f4BdbEu+UWkEJzywyHvypiNgQoH
ne7CO7y2Andf6271qDVag6TwdQU3FFY+5MXEic7dQZUZii4oTJzh47ygYUinvtg7
+K7TftKnIM9mt/ka1idb43NuSpb+1ky2V8PGfBz4D4nEA2edvItEEwQX6XwIJy1x
Vb5d9PrlWZM5IlOfp4r4Su96cjM+fqrimHKrm3Y7oxRTCGQhpj9s5CKr8eRy1xjt
23eoB45uCTVkmrkr+DO8Cr6R4knc48kanxhF9NOO5Pj4UU5X8tQ2MXeJVRJLkuuh
onn9j81krdqoghpOlll11KiBha1Ruz5B48XIkAlZ1eA0CJ1XuA9Z0s/ntYjbEwPG
ppqeUY9h8DyCpVGb4vEz/HK+DqeCZX54C2cxYTQT2Inxe3aQ3gvgUlQKyYqaFIu9
bizfG7dWC60qyUN3z5dBsoPxXnjc2+VcHhlFeatqgCHHvjFTZLS7hq9DtPP0cyqQ
W/K3MkeEfAnxhZt6yiZaz6eFprQ4KAZ9/RVlEzSZ/BAn99WQWhGTVZN21oHt7nE/
q5OVEJJoffYRfAIpPn+W34NKHVJLd5D20vR9b1VoRvM3ITgUz8TSMbS4vD2LQ9Vi
RULyGEbPIhXwo35hbyABHnCTiowoyG6kID2gXbSSyUtPJ3TU9QUJCO/7L5E+6+aF
0496S5ZFj3hhZ9JhkRGD9IHsIfCwSC9i+bjkP+aZ9GqJ0UaXjUaozikpu2xf5t1X
4FBxpG2fBHBPNkAMvQJasO5+QfmDmtu4tMwwWq3xuSfHLvsIafGDh8kXOBD2GOBk
6XSwUGztUbt8IA7aWukEL4AmOjjyILZDH6EIYtWuNjKtQ3LyfKH0mdI9Ip+zivPB
MxiKFeNdSJEQ8B3dg1h5hoEjHqK64j7Y+rNBL4RYm/Oko+yS6xsUnC+cLx/O3DxR
+SJvnzJFxZT07Gz/V3pE6OyZMN7NZNqdfwQbB62mR7uezpboFDGq5WDHdmcWJGyT
koRSftj7aHGt3fAmHDwk6gDZ9DAlkUuCm59wh3U3jCaivvwfIIW+ENNxzqAl/AGg
pk3YEmL5U0X7qD9QIY1XbKZ57COXf5ZSU893bYixwdEyFo6qPBs7U3dl1Yxfynmi
HuU4VuZk4Ab5oanEPXfpy6x86RmuxIawMdQbQT2TsKj2FeUwXu5ASacEX8gZjg6s
LIjJ8reNoI1scTl0NY1RCEoDY+q6sHEK+NlYCh0UoKJJSriSg4YvvEPjw3CdIGMj
v1rppV5+KFFc7eWp1wLBChux1NSYTlbc0s8lvTA3/XRWjnRWQpG3VLzcqbD6HOEa
MXtw7vTeQK7Z1BYYIn3+hRozO/c5XYRDEGdastBSbju2fNgGLQpiqIRcLEgYFNWD
xXRH7MCYzLRHGVjvPsMNtzkCEPcF3UP099KnxxCiY5A1m+cYHFBwAj9iC3kGe4RH
msg5ZVXA721U/+bCjQi05EiT6qouqlJz4rpBXeH35O/i3ZQ9PCOyFkmwVplChATm
SqNsJPWkDl1JCqKzTpAu9YVH+2Q/kbS4gbJkCxURVWWYIqEAWccYk2NJBdG9KgVv
GO1EOSJvKu3eDOeK6aATWwXdCdcI3RCys+BnAKcRo8XbaMLuXp/XCgW93WFZkuwV
4XmHyKK+izgQntRFYVgTXJXeNN8fRV0zToKBwCdnem7afrZRrb9GM7mY/3DDrmsH
+y6E8BMfEK47W+K31OSBF0mMSAV8/tmV7v/rG/L7+q09XgSKix4XlXUG+iY8lPHt
XOPZEVbDz0opp24UqloQNCXGWttsnN9wGk4sLlXEsLVgfs/RDiT0ZxDaaB2dsXZN
TCCfPpgiel0ofHRz63HzAFp1bsbGQKuPFIfxIgewcniqw+T7Qs2g948MsUqZvwgb
C7tDAKzIECgHyeZwzEiA6GIv6GuKNaWbbpcAvw9jxuzDyVleLdMnCJZrym5IdT34
Us4VoihvUE49+N6ZOg2EUbKewENjf83MJqrWBMobbkOGIapwJW3lVskJWnkjAFdF
gCVWwQzi8N7WvFvV3ZT3389PUtErHJuwn6FKBde+r9sHL9lbb3AywIESn4Y7I0cD
RarmNVyOhV8AaS12wO3PZne45Nn7YqKvjki/7Vj4R0uacQcWPi2Pwdzx8cvZi/qC
5URuiLMUkTRxXV1T98HYm37WZWKHqa/Y8J1w9zRFaqs28KgFySdviJTOOSBqAphX
9661pOOXuuOTpVNZdN2RuxkQCA+qb1f3b4O+VkyNe/Z56aAAMn9M14bjtE9k73Ix
d4dCG59VxNmkKnW7f9ZXbFvnyn8YaFwyltzEZ126doimkCHHYYQuzEeWFTVqIFxc
jK1Y7WqywTjazXXkzQY6VEoWzOk+YdJ98eBomK9Tgmmri2R20TxsOrBaUCLHF45r
6fnR4WsIyLGBUSdnUd29oxFBcB6Cj800qLIJEbcJIeVjG0gBaJuAP8df3h3Fr28M
x0X0zVZirM+VUk4YiRIwiBNDSrb62w1podQMHP6hTwzWFOGG4Ohp1WipJdTeihcp
WbmIqjKQu0+N0hvZgWBBmHEKGjDTJgzMk19+p63q8JOhUzBF0bX5Z/VRREfFCrfw
VxogLX9ARzSIIFwwGoaNareGkGJ9oWsm+HG6+Rl6SEiC4L9kySzmdPD0ScYJmsgj
G76xCVEO8+ltAA0/QtDoCN4Zite9D5kc6t2R7kqfC3i9I4SXVWKBEGl1A0z9Iqx9
nuwEsgvxRa+YAU9KocvjZ9lgGekUOM8RLbaD1M5MYLf59vXSaEEEMO/rmN3FqJfN
ur+QgYn6a6QBSYWYHRhKpZEyBA7Do+5JYDea2aVVyg6EtMv3hTMpajMQJFIvAsl+
OczCO5C2gvsLQHZ36OnzpKidP0xpeIu+67HMRnvZAiMaQ1sqksH02/lJM5u46fUC
b96Nejo6fH0OZ0LU27nGVKUZK+VA1fxFzx0vr0HCU22gT/eTRoYAVyNVa6IbofA2
5HuQxjpcuUQoJFevCYCPy/vW4dt83RJKSZlLGjEhcST3QWLFsCI7OWAHPSg0TLjy
FEGJK69F5sGr2mPqC/kZ8vBPchPnewj29WhRURxEfrSHpqgBxwRq4mOegWqcZjFx
GEMqUnZ7MebcZhX+R44nkf7ZsxRAKdPeAv8dINtFcidOeb0RKjVuEjYdYZelbYZg
+JuOuylCXhZWXIP9Ra6P6rkvD3Jx7cIqlGxW/LbfchdSIbiEy0qbDBH0B94A8kLD
s8M47RshpxOdHaOXV5qlqBj5nWqEnyobZuLB31sO7NU7MTMUPTqH9gQBASsQhlkY
atCj0ax2My9Mmr1xJrSHrWSwE7lYHGLUDfibVQ9UvXXzBvOVghsBN+aagKtGjluT
0eNl9EJZ1o7RlO+1+Cq4+Tna5KztQM3y16qqCof3Vs3xD5oI8rgAhVrsTL3SG0Xf
40ihTjlVlurPxDuWW+XU4slmn6GEWDhYgTQGw55YiFMkNz8hbuQPC/dbL547R9IZ
SeUPn/XydyifeLY4rXJpj+zlKrJbG5PwPX3LAfD4x7KBsbZv6g+Mkp4vB3LAtDWz
joPEzQCdkBAfIbBoRg87kRANfEeWSW6eQgc6rg2FKsW4h7UQBysb7prO+UFeTjKr
fcj43OOle3NE5ibEu4IEDuc8KNRU581DDh/jo3v1nPhrMQxIx1wiGOnHlCWigCv+
28GHwyT4y0aAaWitblyifgsOuo9oKGB+8uNrggagBLlC3yFNRYyz1XiCKkdfqThS
n0PXI6KBl2Z6uhas7Jkoe7VSSN9Zr4RdGocZEJh9tt9X3S3t1fn0RuEUhCgVYpq2
HWfwo/+09Qf9HlsdtTMlyokCq9bKWqIBHkRp4uMgDqS9JdO5TLVDkOqZSoD/xVOb
uitaoy8nnPMBUWGhP8rQnLLpttpjxemg6boGgkSnL3DEwG9lQo7tLQ9AnKjadAis
p2ewauj/1NG7wtcqB9XJfMNZx8Yewv7OxHVnuT00zBrgCfrdIOL/K9S5UJhUsZLz
0GGMvkW7UoqaWjN+2g6cmM4LxusNP1OksLbYrdljNk+8C2rnPbeizFjreq7JGs54
F1MIFKgSNuxuIhLClm+AtCRSRWMCtW/609PeDqaUnHqAnMp4LP+QqNyrSFClmT4U
w39Xak6hJ0/kz+nGlPrHMhs+MS2FDcHkKEA0Mw9Kr8+edwTtzn+G5IpM/68lXt6s
E+sWlXbyqEMW56yX1MDbHBclegvklRbLhmjOB/fRlbDVGZuFgA0+1E6ixX12Oa66
Dw0RI4V9He7gloYzXYEfitWdwwxZoe4GU/s4hOHfJhl6uepyMfX0th90HKQda5ju
xotBc7FqpMIUmXTz/pNSEUAqR+xGHKyET8PHqrj2P77Qo8i9GY40f7Jf4JGzTtT6
/ASnXZR6YySYLcVtudb9Dlj1pO3BZjFtHa8H+ZOpfFyAJNYrv3hOaq5vrnLx3xhX
VtFOdpW+Ot9D3S3CQCTP8Odzd7+VxTVikWYW6rjZI1MHvzVgpCtKB+u0sFhmkVKg
MUmT/9lD/zUB28KKpLMn/nIR6DjnGy4Pg5zfykvdnqByh/PYgwYbkRsD3N9ohkyX
XYh5soJbZDPlI0WaeYWP9LubAq98TkLAFq4fAQbWAyDqh1W436vjZQQh4tcD4iaH
DfzQ3E9901A3s2jy0cEb/yheT0sRpaHUqNC6Ij4tpP/kiIKp5J3T8vR+AVmnqjxz
z639PMk78w5zVxTOY30jY1+MLMorBaRNKNWmXl6hRnlMnQPGtSv5xzchb3tkzPY6
7q0ZhLgMmCCFLqgzSoFbrr0yoDwM6SotfdOiD6X/ydjrob870RrfDRaxy1PcCbaB
dFufphgWeNlSFwH0Dek/AC2O1f1yIsg2B2wnuSmoidyMRZ9ijP3xc2lwPYeGE08K
jheEWY+RCW3SQ3pVQPPMD2lckyPB82qQz9fkdj8nkXQxSdwgSGuNMhzhM9vLEOxy
cWXKH863osYJsbQHC1C2dgwJ6xvtv0yGogvHvGHXP0qPIWsEQm9pz4i44k7TveG7
TARAAcc+bgkBvD6SU+DbQ3pcakyRmwYqY7OqI1A+IY2ijxeP3b9B8UDqV9+ZmUHP
NuZfualM+9uIrseu9dP2TkmAr8CzqEBRUx80Xhum5oXXm+xzjlE0dvQ3NXDUxLU7
Zw4iBt8CNp4pYmPOT2j9VmUY/hn3u0VuBJ+DdfMHpjE964KCDPzVAdkBdAG41ha7
SVuObTMPdy8uuIef9voPbcq+JXfIZM703r5dKeViGgUl1VFfSZLhdS68TQDgobeu
6Mqn7PORxSvtMPYPv2hJV92Bl/Hu9jUAYUCpi1E8lm6TZ4X0zBvmHkdT28R4FylZ
0McMu5ub7k28b+6qRyLCZvFdt+JAY2VR2TCs8Blw+irOKUPe5+NH7SOUico0WuEW
ATMLUDFCzpIUjt6M/gBFTM4T+CAO8O8JiZC0lTbL7FHgebIWzGii7XOe1uvfcWXX
2mMnKd6rIo9eeZJoxjPkqgr0JGVR9jPPMZpsgIZcA6/PoHHThl543L2CyoIe/v4Q
s5k/YjcoQpqptb3Cx8jfWeTeQjpS28RbanUWPACcVyjmTThSR9lQi304G1H7sFaT
oVJKO1EZkQ9Faip4uZu1NlaHeJgyu20lb/RLmHpQHUlDRf3EfK2nY05IPhZLJ13O
Lupz0HVTMQaFNYgw+aoWczOgsYOMAAq+9HV0fNDXVocoPCq3H5Pq/jbIPWsgzKq8
HPBnjPIfph1JUiXROJBJez9ansIpvz7Ncucyf5m4o809MJF0CwATcKVeCj52CXhq
fVqmDf/rx2t5Mh5fKxqueRTWnPDhMxs2m5SeI7IH+jtF1Nm65FxSaKCxuMq9SjE9
Wu7LIaGYm46zLmPF9fl4eSj2WOvB/9DnHIhRlBtqfornHuyGlviSzqksnQwVDcmk
iPtnj4HBa3J5qjTZCA4bUsWAvfrotHGV4bK5mYxfYuTNMe9SzIONbUGRlBT3uzlh
LVDv09nMpq3o5AJLGfajB1BJp2i40ppPAa5Xyqi6otGl67vgFfcpPOWIQVwyBQo0
6L5nTxjfX+Zd0824AGxv5pKRr1GLOOuo5W68wZOwNc93bA9NtDk86Jg45R0N1HSd
8qDFFuoged0uCYbphdhyLAAaGdljyw/A8IZ9i+PPaIMxxT0Y5tZtc192hGjdamyo
P9bsPOVX/wq/FNc3SUJsoRnFCJv0NoTFjQlZRFzOx1wCUtlFg7rug3Bzoxebfx5I
TGiDWJViaOOhERmvDYqcoRVSoZKTHRiPj6IK0MaYFApq0Kuu1XnARPxPFI+6bTNp
sQcWhXi2c0PiJUBdAgiwjt+ylfYbyNlwt6ViO8LonRA/4RyHg/JtL4eLt1ESjfAE
wj6OkEqxXVqxRrc95STJD0SdoTb99sNiHTjqBkefxacANROgV/Q3hfXWAMhGewzY
+JUcVDI3FQZwkJKhE+xBFl9OtGuafYRkJ5OZZI9x5OJSL9AWM0wC/eWlLSNg4DGB
WyT9xLQCWee/tu2nocUn2X6wNr9hWONmz0qmdP+YqDJy2pbb7jRnnq+RxsW1aw7L
zIGtH+27QmAa2r1jrhnKFgMGNcQQmrOiXEFZvnbioIWQQGIoz6QkKLj5+P7hCGBt
cveFzdeLpEN/Hl/wJwVNM7CWoggWaJ9m293E9mqkfnMP64UXYSDbW2EyFaldNXF1
YMqRJk5FcDHHPF2/bXTzDU4IcNzRxE3b/cUdfsNYYUQeBL60Z+/CTMlbw+mTF6X5
mG/WEm3CQvKfiRFcetlnAl6xFlJgMVjpH6LvyKuLqCRspAHXHLeJOdpnTtUyRgnm
rOZfxDH4E/g0ikBKPwT4eSNtNxENmX+L48B09S+2aTlOb8eTppX7S4d9uKKJlvg/
Gqy7V8pjqJlwB/MkfUQkj8QB9ALAl0MjyIXki6c6PvBMljUFNxvRcm1ChauWpxMg
z/0JTnYzGqO25TJ2s/ZqDm6n0VQ4G2RXDLoB/im5p0Ldpi+Bz/ocUfjt3FtyFkB5
v5IJXPGv2kTJY9YBBMJ144cvL0VfqNvcCUdqmurUWdcHNmwu8S8AHT5S7wWhg0wW
++EI2onkI5H93c9xD9oln4yM7E3XB8P/GBrOLG69BY7p2kI9yC7CYZoelmCdPDq1
mquPp5djuowhuoaRRqzSV173B9CR+tZc9+8XPoeZ6OeUn8CQ8Fl4tzJIiNCF7Lp3
0HoBhSl14InxXNWYjIDiHPZOZsOAgnLV0oTuDC3MdVmknLodbuRlZMU4qRkYcj+0
Z0/sxN2YsI3L72ghWa99dHcI+jHDxaYw8ZpFz3/jWw+NWTRhGUueXI/Uon4SptdJ
m2vcVCveenhIdsP/rFMdMuJO352doZRBf38sWf0S3+NQtz83y2N3BY0gowMTme/R
mxGwPtMdtKvz/nUbhqannZSU5IqVjFDmecwfBblLiP1efYxKrzYblEV3Rz1h6dtK
R7mEZI0M8AFWAd4tYGRywSXKh/T1lwYv9fvJzCyBO/6vjg4Us/oDJl/3y9Fv6SPf
Xw1rGeq4ZqzZr2VJ+wpgxXVjRB0+QTR+MxKMAGgPB9IV6/zKUPL5qAocdTKjvQsD
DbXQJUARq6Xe8ZfqqJ8L5XTWlICgCU6LBKC4UR0btLdJMqPLaB450jhqx4vRtWq6
Rv3zNxP4QGx1OuzZm80jNP+Qw671KOl9zo1Ds0H9J8gug12YVNj0yxngC6yxvL5n
r1ewD5gb9wPoWPA6XXvX+2nJneVaRZKxUbTDvXR/IbVlljOE0pel6hCBlFqvwtsm
0lz7aY3G6fPCnumAhJ0LpkD2l/5b+p8Gmr8b2YHJ2PBMCwpIUxRxOQJjziGR53ov
UBSboid4NsTd3/VegFZqGlAbKykb9UT95aDXa8Wwk/fOhZAqsHbpoDOpj4+EEBuR
4aVMFd3oegWzqybKDv6ATrYHMnVNGHZhcynW5NIWWLnDiR1drO6vp37RkycRye6i
q+9g4xeLVNy1GpFOr+9DTtcdJ+qdsxOLjOOjLkcTRqbXkVhbPGmOR9xnGO2Z3xKe
cWyfh8WyovzcKEFgb7PN59FROoclrW2zb1faB+EFAhy8K4LEoE2y+x59IAErRRRT
3CkJoChDRI3DIg2uV2IvHXUhNhotcLe0O8b76hGbau6mtIpEHO9Rf1AXZyZdbXjj
bbM9sS7JUZf2TDwd6pteSuPLP3grd9UO/qTjnKI6Jbw2VTkS7vKT/maWcrfPO+2u
3GcGqnx6BVC+tmoiN3YnvlI5Y4S7rVoJdibw/mEZRd5gvCJHCtj7kC089EMKG2Fc
lTNU7zZhxSr0SG0knxUxdHJYcoFhpR7nqxXuhzNy08i9oms5fW2ZjEmZsAMLOPYE
opDFGq8PEPN7YyHjW6B8BlUPjaWTrUlhR/7sad0ID5LgDohR1TxIlCnH50OrjK02
LnbvS6mb56GiNrt1FfSWG8O/U9yFi2X9rm8bhoHKS09SVricUGlmp6RXlKdN5quL
qK8oDO9S+yefpZERXswchFb7CWMrWfeK06ncdJlEmg0+wLxLXN74PSoh3oOiRVUd
iezeuHcqNKQLY8ZGlpvMp+c4yUNn65kXdTmeLmfyAM0SbSBCDFiCGe3/7Rmbd3Z7
lmWCr3LqniPOoZlcGGyWK8imOOOPX5PHC/Z5so4d5oFe+dGKtI9UK+eKEVSXXAQR
7azHBHicmiaiyiUTKdnWXLF1ueyjW4P+Xt+K5e9+GqhpvAsQi8yWvJ9rTnVKnr4E
v3T38HgN6ECc1YM0YmHkYqfoQDrvTJOruaNLBZZWxsMMDSaQC52Ww8EOpwxRrI7w
xBjOmr9wEIwijjPoDNTbPyOq/qhtbVNekVvCRahIh+EYqAjp/xORIcTBCK8/UwzZ
CSanC/Z1L/s72zwBvzSZRYR3zrJbShMSCU1LpyeCVry66+WizYEOjSg+GddwxDUS
yAEBw4thC3BONU4bEvdKEhKDLV/+HdNihm+BlMEZZiZIrN14TuwaZYuRC97nwB+d
RxIsThPPwLQQBPqNH7EazLHeqyknmBLBy99xf08ShylanF+JGFO62jkWQAQddhCG
DXYwCkseZHsO7K4TIER+WXtQsZNIJ7R3wRKoaesgUIS03UkMHwAYAo93ZtR+16cB
hrkAMG55L2lEBuaXkgs8eRNTWxrQpXMnocYk+37YZKjzZyxOyVmDSt35V7I7NASD
dCAwqTzMTT/brNfpK4LfKrkWE6Vj4VNIfKJ2KpSFB/SHOwdNiUY5NoqdtGJoW82H
T8nQ0Dx/jLJL8FD/qwlXxBXZhaQDMhKK4LQsUx8Q87ubLr9q7j4h6DW0ifNue9KK
sEBC+K314ecxQmPaiMQqGcD5pQYiWNORuabvaKsIdkrh02ss6XU4NqhkSmxFEpLF
DDqIyP9MXB3CHwEtAqq5C5hJeabhJ8Wh/jGuyb9GR3XImC3JRGjWz1t210Fszzyp
dEL+gzK31hsXnrQkjY7lmwtkVIaMt4r1CEgxXAUsAOxEyd8jr98Nw+BMvLdNRATM
Xc8KUjj4GSpjbgSjRyOXgV5qxRifVY7KU67ZDnamEejJLfdp7TywXiVgwrkVhWB/
gp/EbqgkCWl9AOMs5OIVDDx9jnqJE/BjdtVHG3pTIAT+mXrlMuPBboiJzxtXomoB
lYOF9ZgtM0ysrjWW0Ipds3wIwCwEqFsTd9T+iJPtMdjcQTuvqMj9Zi8GE72mPpLh
eJm3Z9a/6hWZqTeiPuWj6MijP2hDiOPeKds+/2mj22F33Imo+WHuo6u4SVAxogYX
XIHilUXjwfGXioUNUURlCjFPk5oCjWXSpHfotniV+va3FVCEPe94D8dyxU9o5VsU
HY3yKZYcBiLRsk5hikpQ7NgNo9+x3M3IhVPQTZuwiBx1s40VG6meiXKdQKQ+Fjho
1zIdhFn8sLZ1ddvRrbvZigBo294Z6O2njlL1PVljYo6RCK7tNmOB7X9e/bG3ARkF
pIK+hD9kqkC5DsNVcbrCj1SGwXnTRlZoYy/jKai6pc52ha2+pbnMSKZOglPTNpX+
2i7VGcf08rVHi8UdT1j/9LxgCJUGmkFe/njMv7/79t7IcwD8KdMuCbFXds+h/vWu
9wDCZD4qVtVsNct/G2eefDy3SC28wrEpyBfAmi38LDJwkAWssHYHEUVnOK5dj8Kn
AAW+zZG0gfRV/vlYQTQtiJT2OPlsgeLlxzZt2JazkpI09vkwsHmeqU2XoXUz9rkD
l51SosVmwG4rWjSveBQI8h6U+uRcPrkFTDGFjOktOCA5byuXnkhta8fcp8CwiGP7
OimkAjJUYtEN+wa3ZDU16bonq7Me26ktOLHjDhjNWV5r1x8PGtEs+b5LYpijSf/i
YrvZkiggNgLDHmiqnlw+Dos/8BN+sAWAgvUfJ/8Qdm6RbEnYWBtwC3kEm1IE+9xT
HGLhkFOnq/9X8zjw6jKC5LM0AzrJ31DEPXd2DywZplHB5LzjzN2+Dxn0++BizmQi
toudKdoHUxuXJlMq1wCpbhxF5u37Wojxn8kQScOeYYBSQA67rFcmhjHT44m2TitZ
EW/ZJW2dJ1k8NjI3bpwe6Cbn78EY+iK1/TUNp2RR7rAvbjua19QHSXbduIdxahWl
jTgMlkdpR4H1XMq8YPKC45340ei/wui5aQDEGsM8yQHwH1/O7ZOabynmubAI1SHh
6pHQ0fHOUS7o+XldzjKXNGGEF5FBPp1eWfsNUFgRkqrMIVW9A2JDrpbzkP09kzQp
DCPIsO/Afw4MFk9ZMutRUiQgp4LZZwZXrz4OBSO6rn+8nFV+AJq93Zd6KcxLSDVL
5qxID40vpZazmqcIulw/U8jt7TI8UU4H2J5Xg4vBcxjosZY8Kvn/Rue1P7DgsyYH
bDN24BIm6xEBTcvtez6GpcAyYGzsM1Ug+p2Vz1b1+hXrAY0/MdDMOOz7HGvtB+8Y
L04tiVZwaYEEW+tyHQy0eEocfc3SVKThrliX3xZXWAvB8MVEixaDAExsGYNyLczR
S8qkzjEO/1J/myAbQedFPgLqBDr7g6NqFcWiPkzyyjtkgqtxAxxjP7jjbjUu6jD8
Lb1GIStu39dw2Ex9Xe4Ih+zwbWrFbQqDWfvvZAfYm9f3kFM4vc51TTv19poxcLmC
bqFKVblcScwohkS23pF9zoG/ncyE5LnbFVTHelZ8r0SmBeXIed8uLk9wSi1TgsXE
qGIVvWGu+scKsGIPqIaXl0nFdK2mmuspPWz1r8o8VEu46+yQuyd3QoekgKTu8UPE
/hCl6Vk7AMxbqqkEL364q5heOT6+3l2v2qaE8DRvdyxW4wqPyFhkPGMb/jMOr6hc
9f/A6s8OW1w0hgKUXl0/FRRddiSsRfGW355OVanhVY43N8ZXiVgaXDkyJmtpoep6
vgsgbZHh4IQpkn3Gy/BhNgDgkR0TGpErF1bzYXUoARRBIDkEDAZpG+TCsYoB/vCy
kKOnA6bIaqNARTOosWoQcXNLgNAdn+RqM9X/IacYknaemKzOqMfbi+wLKpmDMGQ9
FsDXVzHePXx7KFGfJmcbZne/cO8PbcfRXcKTgG7JXVNe0IdudinUsdxnXQoemqsF
FatBcSgWPzzyuBKUJxwQ7F9OOXkPZXOAgy7Lu2uJYeYSCN7EmBUqePdOAGct1N93
eglHx89RZNEiKwM+34zMKsnSlNYbEndfJ2ZTmY+UgPBVmou3o8h7p8DNf585Wk6c
UIkizOnDVAfuzSP5Sk9GlfxHm5wG53tSML20LMv3lR/wawFFBFTx5aKEW1fhT6WY
tVbP9KtuEE0d96WZXfCSBO8E9aXqeQVtzOn9dxb9oQfpV8BsvDwTjz4FxQddPP/S
/vjHPq3Cv2tPtoMoVeT0bkvZ42IGFhLUeHQYak0zWie/9ip/m2U/TIFEerklCg2Y
qebLYR+QpXfM572rGN27FUTbu3z3rljzeCjNgjTqF7CQtsbZlZD1Anry/6dCPMif
M8LPf3SBNhDGkCGLWuuxvIkS/kuUbVbbW7wZr08wSt1pNqQZSv5KglYXv7UHlglF
DbKucw2SJZKOSNExS+IcKWQTrhiBIK+5R97OmuXv3HeYMd0asKVzB0vV5eIbtOjH
C4utVNXBylO1xl9lrX7F4s9gtG7jzKjrdA2m8YTa58/KVlPtgu6OLfDQChm0qsSa
6DTqd0sa+yrAm9SUsWRd+ecc6Z61Urp70sUbTBD8D4/nwlvUNDIoEJoI2PPp5hOi
4/YPEBeur0cd3/BQ7hRfekv2OzfWmtcvQTJ2a08zJ6Xl+MYXk1YQVd0bYiuhuxl+
RTqoEp9kL0rA38LbVKD6bdLVwgWeYdDvLEWp0YIaXfbrOaDQmOVjp6pwDQkL8e9h
jeZJyPuThXa4N9FWgwMPKmlrvoQzE1XHQ61KSpj4wzNHsoXbIKGik8jQW53c2JKS
lR5jj213gF4dK2AWqDUmK2pskCRYV6MgxjSUFCL2F8c+pYs5+ZDDjTqTDO87+Xpo
I6A2Zbo+VCue8BpmRf63OlWNc+uAmDUw6TB8EtWdxfG4e+cz0t3pL840tpijxOzA
fGwT+d2evTlla9zmuaoCe9XDd8Tb6nM43upWyQqf5rfY24yPtM39IVJ3XCCwMIyU
Rn/xBB0cqeyEDtaf2uf8RlowtEstqHK7L6oe9ItHWX6HS2yQpRHuCd8Q03oljab5
vt18fxfTGiCb0YZAn6rSq30f/+9nCsFQ7Qf/1MAPFpwSuo9RogCmvr3o83hoiB9a
jJ1Pt8a8X2fQUKJX8ipAj9S44NLgEkcCQ2/JDN6Zw1qOFepjQ4NkaK3q9VvncHwq
YC3e0fgEZX2RdZ/sPRh4sW9PlTS+x+CeDAPws/3mH8wVLc2DS3c0OYk9xeOJd48d
RvzTbcvQoN/h72LYWLJ7tlcALskagX4CoTsIggXQ52vHZexyfXPHGyxN4eST91h8
4VmtJqnrIpOQ6G7pb5djl7D4WNWdXVa27edKFjoSoXRiTeeIWWZWsvSQXzpSTrnU
T7NxZNsdrtOXiF6yEL1h8q6jxjuJKt3uTjOHwWwN4Q82slKlPa/Os25WMtAw2vU1
c5/CDchltLU1wZB0Pa3cs187lT19soI8n/t+xz20tnSUxC0lI6UuMlQuH4t/49DW
WAsAyTGuLGvKL27bgpO35ikUUJUb5gGdRK1rFCZBr482OyQaX1fS5wp96zYupX6M
W/4rSSYgma3ej0DhAGG4DkXaPINo5+ic3oAa+qTDIbZEKNePxhvCEvJMK/ValWWl
pA245Rk1sHrtwwxRaXn52MUafOGhQIycvRJUIv3QwVtC601Lv4FWyTZWep3m2TvN
3fsqQ6DtMcsxdHLJtof+9UtVsUdRlyhGHTF+PE4vrxyRIpOWRShBiGBI3ZzbhIyb
BxJuIJ2F1OuN8FX3rLcfIfPdcd7s5TOluUjQIaf8c4+18H/jVHnCme1BBgZ9E2R3
4C3/RD1u2Yk4aRpf6SKz3CnU+lRO4xo9R8mA57feGFZGjNYuF7LQl1lv18xOka1H
PstFRl73Wr2F1tuCaXGbJ8U+EAm4MYHwoerqYZYjj/zS9LZL68Ki0Gv3J/SQTGLa
J05+NFgj9BTEtb0k/VqQqSozguanjJs4eNPrE4kguMkuttP4fOEEJrXFfXXK15HF
5xQQ95w2VjTbXBvUg66siBwdF/C4/mKxVsYYCqdSYjynZGCQz6V3Ut9XvVxu4B0Q
e7SBG2Oao8BmhksjexAk51H6pDNcSBTsVdfIWM8Pp2Xf7JWXBI+UNqMp0khy/g2d
ZyztCOb0uBhiOdq7hilMkqrtGSpjcdoh6Owa0Sto/p5POwvB4c44K3vxgl9U+oW5
oDTIoDyNyJ1hRQviJ8p8pOY790Y4fS8Sdby3XLDXRlns4PU9rFk1KxAGJWR+zVFa
uKFqOc620Z0eynKI250PKod+oWNA3bE1UW/E3S/52kwv/rv3vKQdhfOaKHL2XUDN
o79ImZGhrHbnC4so8tHymdPdENdYEJda2hCPWxhifZdZ938zUy33sG4SveDFjinU
3X6/A80NLhPMRwesrLaAn4pdu6A6UMpTSCzHUwY64HVQ62nkhpvV/3ZPJqinmbOo
0IMjJFh/rG6AFfvfWxQ9UPwD1DzkmHlvf1L83L3Vv0v9pa/GbqJC4aIFGFvFb49h
EGzpP6K9WjclD9gUv8YX8oyVmkHbFjuc/csMhuo6eRORGSWeOS2CngqUsZndruaz
rEvnK4coTQ95m8Hzr0j85bjqyhq97mCMCGfKvYxGiY39ZkezSrfVzILWRGjeSEm6
wDrIT+/tRgTmfQ1WRyKo+d4VE13de3BS8/vqBt4T/N0wkTIIDjxMegg3MepAoVW7
aTxGvmiRPcEAzGWgnxBHi5Oa+x3/Vh8xidrTcgBviRsMba4ng3JsaSPBCKMlGQjy
If7de+hrCB0GH6f6VbQ8XzNaNWl6qtBu8xbQM/MgKXwLtnWbTJEpaRcZ3VyIR1Iq
zC4W8vC/cu4fGYQ1FutaZD+Vkm0L9UyZCI/+RVxQvhrp48P7GAxVXh1XXPkY2kTK
J4mOFqu3+nm7CgxkprFTLm6PuhTXDeq/b/5XUegPbEh0Pn+8jEdXBqpFS97FEiS0
FVm3Pk7+axnaaLb2J2C780U8rkQ7uNJsCO0etiXxG7BKq/3Bi7ysqdVNs7Q4Nx3O
F7/au9NHxdBmCDe4FhrqLQOJ1Pra7dvhJH65+uMZq9IHV+dfnYBOMSviFlSSUYSe
suFOT/iVG128jcJAAq2dgL97ikAxtt38ZgCg0Ol17mWI7xlstQvURA52g4VX28jo
Y0YvZ/7YtuhcZMod2CleQCdQrkhlxAxlAxA7xA/NfviSLvtG/uZKMFFpEV9tIQVP
Fvhb+GOiYtEuBMYKbTgapjg6O5jf2JNZJ9OzDuSkfbRxA35qvm6/089XK5gx/irC
OWSYA/HlxaROHr+7OGKpq/8nHCib+CrcYOBFJzU05try1aekaNNayKdfhSkEcCwJ
tm8FogHuAze8S51NiRrDii24SGRhouMMEOUDeJNq6CT5iUoMJ2WFery7xoYuQxZo
/AIOZ9kpAqwAO78bYlWs4ntutJTNFpfmNry7wDH9Z6HnA7c4Q4x927gCjDA/vN1R
EHLmED8CyIlwI8VnZ07lLjco2+WjTYvEBUiuLQmQIu795+pkBDLpbw9ABQMYhDkD
A1dAAPqxTXd1LdF/QlohWKV3nTTfUg59nUak6/p/zbVTaMJnJHOZGOo4EUBVZWtV
a9bbzrFJrZ+FUFGnGMEcXeEKHnBIXJSPZJpPGhu/hDYX5tL2xdL23XpMLlYda3XD
L6HS7cXIRw1/JsvYeKAZA12pgTHtPEEroyvhAr9j66Yb4YaT6jza/YOxitBEBUI8
mFAt5/eI3goJAhnw8+4WvSVYeE8l2b4phU6aEAjrgTx9/K5BN6iMqaG+bkYbBMi0
RlHGgVx5hjEw7kLxI+dcEo06qOb2kOMe4/KCS2RvohHhbrdeRAYr2kABqLn4ASJx
i14XrOdxg2M5sLCeyTY5Z0TkQl1lf8/lJ6x7jC+GUf1UCmfVmm6CTfPDXUasUlpA
Bk+iVyN9EjGa3rpby3EnuZz8x7KuhB9Qpi955M250MVfy8Vp42NQXa/T43SJcPca
UfWqPGcFeullA/ZQNDEoLmUdhhWTTPdF8PS7VE9MOsyF4KQqkmmQPCyBIf8hiA6l
xi+ILG9n4jseJFB3ecdP2RLRMfiClnWOhrsXBvjHZNRaCIBWKT3csnCryZVpoPnu
44KzKhp/yaMqUjc3FSpId6/cHRUitSRCU4LYKzkcHocto5gs1XAA0WK5P0caVKz7
xyhnMZmfohatLOHjHpiMLOfE9xtPJuvZXvd9CmuLRoKiYEZ7sjAkwRULaOePmUZx
FZK/mW/NDMnIxQtoKYw2ESDPapgQ4RKLadbsRYqL9GFHEshZyWSUbi3Jy3BHiwAK
V8GRp9NtBm2OupUjBaMHC5jhWQ5lalmWvhLJdaeUwBD+CLr9pCXIuN1qX+o7lt3F
S4JHYHHcnq7kgddHpERf/aPk/EMpSak5+krdUUaG4hpEy5vJ4i8EYMdyT+KfXx4z
wIHPy3ToVAapmgQjieP06Y1sVc0UoDeZl11d2LSgifOQjJzOpQ6q27UxJzL9vrUI
5RGQnpCRV12H7aTb5oWK7OT0hUlJNLfs+IjkwbV5YK/koxFwWVZAp1UJ1yy863PB
jPPd+qkq/RSLIwiBsX7sCd6UxIqE7pu9SgQ5tpGFZe3k7dzoaedxA9Tn+KHACSSl
Y32gdoD8GqYu5CoxbQpkA/PMXfz3E7zxYGHYZDp61EBprK7lExh5X9+19WdSH+Fl
sxTuHo67vV4d5PXG/0qeKWkNei/VQe2xei1bq+qxE3hKKxRQe4Oj5vaJaKyeJueQ
aVBg+XFUcICrwr6VwPh/gLmXnu6gDhL94jM/dJeUpO7I3tN9bv2XVFdXSoQoenwL
TUl7tlEF4MkpXfTRqESLptqjIjKr9J1jQvjMDNebplJYBaa3bK70nAQU8mbcp2M+
PNvwXkQ1n7vHIqH3ahymqY97FyIRqqKnPSBB821gFLnb9wCKa5pvAUxF8/Z6VWSK
wFRljlGKb0+HJ68qLUMW4+A9qlB98WlP3qc2sixozCCCABKgq0WmHUA+JYr9uG0p
kRuBOKqLsd3HXq/rIaFcfDHuw3oGqOAFEOAc9WgY5LC6fzaAlF25e2OPHZ/JyttI
eJJ4/V+vwirR7rGzVmyucneTJwq7pZRBR4vNmM0qEFa8YX0SlzqAbRpwT/+UFhJj
ltWK6pN60tKRE0s1OQTonsXGypksCUA8u6hAeHaPoqkm/W4H0qUKZoeB1yR3LkXV
eiIrtXSLdxsc2r1Sf53oS9rqLTyKpInvjauiRNfvitTfJ9vyeRRG8lirI82dfp4+
3inUg+9t19JeL9+SyXt4R8/R5VZs1twhRwKCGtFdzM8x42qpLGRjYoM7XNNOj2+4
Y3S4q5JrXjfUFE7yx9FiT9PlsMu2cLHDSsZSOfeyi7DfeXMcgLqUe2CVJXIIVsEH
Y2/KdH2BwVwU1riVS8M2MXHl2+yQEqclg0hDqIiteNZ/LjkFRECxwzyprFoRUlh8
uNMywrVoHv7/nvAbNoBNRYkbciXZZrbqClNZDDqhpJTHza0pXcovljBCs+O64f35
48RqCqbHTp+k2IR7mzYazYKwr3AUWM662o9dCqzdk2qnFzPk3RQ5czbPyOwRO9ol
TSMAgNO5HPK+VBh6Tqxh4XG1Y+RrZT9gSClfA0tpwTVL82fFQVM5m/EhTHk49YCm
8TKOLXydN/kpxk7uSlA7kp+iNH3IlU8iLMjEkJ3vq4UsHA64RkwHyViqqIMtOHL8
u3fs6/tPVWzFIQdOm7XOZl7QK9TcZyH0gVwgN/Fko2HtcC6GKVyAQcJxq/UzQ43o
V4tlF7G8LNnz1b5A5B3Q1lgpcjEp9q+MHeI7Uz11wQ66OAwlbaOoqIhRPQArHEOU
W1Y8kM8VOuF0jGzFy0XBqi1/7XbjgGpa/b8fN4U6HzjJ37+DxSt1s0lt2dtB9w3Z
4ufiwAUOcLGODMn3b5L3kIuzoz4KyMU93mRI3ZphSAm3028SIa3UmH5PSkhKyA6N
y4vA0/9dRvoabakpuSlwF+UWssgpZMXpy7zHu8vYdVwDwiU/ZY8c6LlSzsXETTq3
TJ9pNT8zYd9HCZNcv4hB6grScTAqlbzPP3CrcwiHIDTXOY6+IhnhPbq6nEkU0soe
PeLMPxfJ2zJ8s8Flfz4JpDLqi6htd8PXxoAHopXlkZPHSIkeKQzuQlloj/qLbpUJ
XNW9+jzCEy10wfP34ha1uDlGKPpfw6NHG+sic+/pPX9YCaqIffawKqGTNGw9GBTI
oRTTdx5Wm5akuiVTlbBimcm86MNMMfdjE5e3jaOr433B17SubD9aoKZAzdyEpPz8
uJ8WgTctz9c5JZib4fcAyd7SDPiDV4DzMhC72IZQI96LkgRL5KfehBOSzNxXyKnf
iLExckGsPbW0GxaeK1iznJydcw8BD3btdBLaWiG+OrnS36EtnWmKfIYohk2aG0TU
tw7SNvyfQDVvkhMzyPHsYalyFbEk2hmrtuLZq1s9JCaikMzJu4YQ/OfwGgglLxjI
489UQIGXwU6lBaIaNoEIlgiNkc4TOJSX4/1LWhd3A2rKVE6XlNP8Ks+pWFOrHoov
/lRCMfboMMrfyt6mSkYm5XDdSL/Nr4CDbx+cwkhD8K2fmhvRqix5+HJjUxq1QlJK
NJBcmzp0nSeO0lswg9+ZTVs8r11rX5+NH1YTiAzFNezdWtXkO5/TnB4B4KIsR6Es
ixJE27ZST2BxkIU3fFmQjVZ+Jk9rZhlHRjr3OZvUMytAkv41NVUPwPmj3t6p2ieo
bLSyY50gEBd8GrR0DXnRgYkuKG5NM+buGtSpHNYgYE0V1jG+JZ+fbsgJF4EFy+8M
zl+Qlep7bqexdTfiaWIhFRrmOl8i4BOjprsk7B92CbTNbVUQ596HhIpqIpmyYmYt
lNh/K+1d/S13+yNKzI7YG8qxl3bXb4kqgQcWc4fib42fjh5LuJNeQWswgV37vKsZ
D2k/QH0/Qyigqjv5geCnl+tU+HzXwUee8NgkHV/Q08RFGSY0RaEbcUdAEqgxGZSt
0NdOuyjt0yHyzDcsOz8nNIMUV2Bp3eotuDNG+Yn6eEQJnMBQ1EoohizZcKfckpgT
XiC2naWnjSYC7vu1UysKw9lmF9WcUShDjPIXmrU2TZiCPT2kck+EJNxnUQApDSq6
JUT98/bIcDKsrov2rlQlQ38MhRJaU7TKpakNNKLnQxySNpwWrWUUvz/cccAQPgjd
HEn9X136SS+2kVgTh/shiEcFGf8mlJBYjF/KToXmoqH9Bc2nDt4xchtknrg/bvDS
ex/d/9/PVYFhPrrHL0LnRCRpST1bPfIG60Peb69HL4LTEzFOWagv6m2BE63uMio7
hlWLTAox4Vy2nv/aHoOHkqJAfA8Tsap43SfsTZd1ohmbqtYovv3csS8C8WX4jHJ1
yR3xAKabba6wS3tSdSU/6b/cq85ZvIBs5riewfxbF72fySVIc3jz5LxEhYa9G1ZE
A3S1ea+QzX4r2+h8K4nOYv32ipjpOsKG2BPs6+zDC0s3Ewf1SizAxAs7RJruw34Z
g2WxEgcBNZKgAg+yCMT+2QBRQtRe7HBFf/wGEP0X9kL4bn35rnLgtY3J4L4ujHUK
BGEmGAMp06ARditq7hMpkr1xbT4PyCYRJhgz8BYkdubbm17OIxb6GjkGYs7rfuQL
i2RQz0G+vjEiNJS2qWtm//oBPNTIvhvTFKdgYd8x1rHX1QKC/YOHpfuHWVOPli2Y
S97CIcnIN7OlQwpbVdpFFjrdjuWQxO6u39RsZ12/sV/ZnHNjS7CsZP9uW999FU7/
MPRpIFD3aN1UTHMiyAy+JoEwoI4508uGPoO6bB0VRiQaSDGb8/wDUe3D94yT3DqY
eEtW5SiHBaULL2agOgBQCFkA8gk0Kg/628KW5CpeaBCrMDrXv0ENAi2RqCfSEuvj
B99Trw+P7O/oVBtEyZ/RzpL+w+8mpKMBh+2bFYC0Z4+TQfQnKiEnbnkqtN/KqpTG
1tUxns7ZqtwDOSd8Tzvcvlr5xIDaGgUbSb1x/4MefWt4mlQzP7ZJaw56t9tieNfa
6YJRog/uQEuelNW7RqLES55a5HTDuLUZuYK0/FqsQyD3XX2oVuytABfLT+wt85Ew
YXeTod162/oyZvPx1fa5N8NtzMng/svTExe8J734uqwzqeZSdFQoBJuw2Yz4NFX5
DHQVDd78HtrOEj8t8xfLNcHv0l4/0v5zDfiKashC6fX/n+TRa1wrd0u/X6l+NZzW
ruk9P1Wu0TVtBCeB0UgnPiJ4QIC/LxSIAqrvCMVXEXTty4iqARI1PSsW2a4A5lpw
P6TF+19l9sLOnmh+ORanYNeVyVDD9QsIyAZ0o7j8XbR3Qu9+I9aP/ScVMpjv+SG1
OMJCd2Z3QD+XzrtC6/Gvhz+dXzt+p6f0BYgHfC1UUT+/pUtAtUHPCmdXE4RzTHAe
IEU6W169f9+WP0VJGW34cxB7A1HacBr93S1QZl4AZHGaEfs6GPBaKFRvW5gHZM9f
Mz09MBzlbNnreYzJMk4kmHQleKSUCky5lBs/35R2h0KeUxm1uSpcfXBPZTjFaLAd
6FTBntKpBRFHWQTbtgXa7AVj1nYetZlRIPyGJhz5T7OJQb/hETQo0znYmTN6cWKU
2IvlI4wYw3tmmjOTEjnFjRtqz5L6a14hAgaI/v1QB5jB24PlAczNJ7KtKIZlTbH2
0KZ19Ftq8JwiyN9Rf8A9kHgEDjfGfDHDRE52Ath4lPP7qD9p72rWDa8nawzwAXh3
rGWAi7dsZVbFN10nJZJ5uzJhp2GIcD5JovNBxqxpze7gKlOrWToXsyQUVdT+M1ru
w+7mP07aen46oPa0uXCpVGY09lkbx7SPAvZoS+Pnug8xxK21SA7A4TGYTJw67iVS
TRzRKcgysMbxCeD98BkqVT4dowxQv/nkAEZaaeQ+FiI36TVf/x1tbmLsC/gpwWr2
G4/AeydWFa1yrK2Rco6604+UlG0xwe6xyOKEt2OiuJTDWRO4lMYdCrVZsLFITY5L
vWd1DKQcHMgfw8bqdjt+nNW5R+4ci7doB+vr/9mdyHtIHPoTSEOIJyUfx/0Hb8H6
OJYnjgyY7KfVd0DbXdNKMOaQrOw+srdZ6HJgzIe+fef6pVkM7SbqNAHXbx2efpQI
AGOAKlqIhnPmoq8fskHpiPcyoAR1Ucd2PRn2WBcHniIJLwHDqbL6Cxti0WNsfXrs
R00qs9d/vdwGJxQ1p3FjxuwUDDVOIEH8zl+dJ1M3fzSSowku8lBhfLApePAwlHyC
9+Bb0hbI9QTOAVOQBCnURKgyjHzAkpCYyA17x1S6JBbu2REIMBQWmtiQ43FLM5n8
Ukh/kZsTto8YusTGpY5VHeSHkidAvDaJ1bxtAEk6slVZCYzKKkekcvl7jKqbm4hE
Gr4/nN9gXtSIWf3wfGzprI0OmfOf0L15qzXXcvRAqFVtOxToHPvdEiGXhL3ptAnR
Gh9LrF+503uL+oldPGhFol/mV9u1D+Rzcwp/gFnRmI5qG+81HXb1+Yqsu2YPPKeI
4n4tinSDVcPYIz1pmEui5SHmxJmkEx9lZt/GIQJ+Hrs4sYNWotX4dNUNrpF3uWeE
g7VD1kcgTpSI/p5ovLOoVsuGy8fqilO7nc+txi/V934Z+4SsYzN1DgLUrB/fsRy9
iBSoUN9l6/AmncZh1FSr+zLbrBos015jDWXb3jhrCtgcDU/yzdP2zPY3jKRmmKMo
BkD6ty75QcpgD85F/fa4O4/65s2PfNEP1ikJ7RuR5f5NH8yG/s7jjKCegzmJJBHg
od5ZDeBQ0YdvBkC2OHMf3jTLOjgSGGZh6p3jO3bAc2XEAxU9oOS+pCWQ8rVMHI+P
xj4eOtPjFe2RSlLtH1UuzsdCxcJeV+oMgL1w3l7R4WmHot0Wmg6fz4HtbiFKzSkk
hWYsS+y850fDTvJrNC4+C8YkwXRJWe77Wf/W0pCaIWSDTiezIT4s3BuSZRyQpXw/
Q7cubE2OqiH/15H3Juv0+cdrvHQ61K6QX36h80ucbENgpLjU9AuRGfvPBeMX4AXg
ZOqDM2/sCQ9pLziPmI7j1lEn9rEYM79/ulByNvPwAQ+GdTlrgJe3TqVU5XJR5MBC
czBWrdjbT0xZDd8lrrWOIkonaH6rYjLIVBpvCTN5aglFe0xDIr4x/IR/bVvSEOLW
/dIiq5CGgJSLd3Lt5T5e9j+25f5XpBwOBgW97hnS83OWlq3l5i9Z5gucZFMg7bsE
zvuWJS0EdIaN5uN6GckGGwNq09H7tnESvv4uaGm4cTaPXa+NxRzRqoDQUo8XyOAU
mZndSiNQ/i3uqqSoVwxRpPswMQtXp/Nu1YhoLt8vxNyI2Pheiks3vY7EYdy6z5yM
XG3AKv7HvBmV4CP0dtTh4V9DIj8NqAHh3Oay/EmT/xxLCEKz7hz2K5Lu9irNac2D
71fSMkaD2ELbLy4zyr4bYIKFzx6fAxe5w4A+KXiyJJ0eKjba7O7SLHvDzR9sD0Rs
KwdshxdLhO5Ue8BuK0mjQVSIGuWtqUVyJumUHybCh5oD4kxt6GEoYlJx1wroVAbQ
I4hEsk10MOqlPn6kwSUQyLKRyI4XntOr8m6ACLre57HOlC5FmcM0g8dSpf9KQYCf
bX7NUQ960BOKtm0NUSMpLpg4Xboig7HlosWkZ7Rb2cMUhO/S2czmfi6//MoUn0H8
hs5m6nmZgXyUVi9/zDb2JV2yXUoQRxdqmQb0oxfC/tn4HoBnFwD4cdTmcnQc1KmH
G9OpGjzYubkXtfY/bIAe/LovxVr5M9imvsUycecaBEkNYgFBS8H9OQ6+aLGkXmLt
hbF5oRaGJoEDCNJjm1Sms5yIdc/noNrOwUKfHXRY5T82ee9z3UCMTRl7uHEKJUva
avhIc1gCu3KuK5rZtbpHNjm70BHBcJnX6kMeXAqOV17Uu6DyCWY3eUHaGET5FjYf
VtYHh/7QB0ql7WGw8gfHwpVnA1r1kIK04vE7jnOOogJ/5iXeFu518hOboaDgczyc
tY/SW5k73qiYUVlt6vifpgkqeHwqnvwTIYuI/Gn0BR7E01GuNkqPhgkHNqbgYTbw
LC29jkG9OQL5aZd7C7saOlfinUEPgsblTh8c7BDxynPcVOED/cCTrRcpdDLkIAyV
+BEd/n665A0ivd4u6sma8M6UM5L8XUIfAU7x99H1BCJwHChtqdTxVpD6u0m2ThTI
7S9cQGeQMHB71xmjBsWzU7Y+Qu9BNceGya5OocnGvOND4Cbu90qDoFGrBtXxe0N1
CPIyzLhgqScEVmIc7MtyObzbiJ6DJbhR8MWeIe+hLIA6XSZQpZR+Mj6LO/kXwCd0
xdBIDBGRV3V+Oo4dO329fF7VdZ00JaqXFAIC1q9WoSgiwd+9rPICx4//Eq8gOhdN
jgWn2usO0aRQWASGlkXF98j0XfhsUlIxHdp1Ym9azsG0l4/fCma0qyPFwyVEGvEX
DOr/UTGGjynUmZOg0qoabArnsRc0YbGSvAg/AarrcKxbgqcqj/jF83YN4VJwz4w8
EZGZxI2rJ+2lFOaB1o1BkJoCn0HEa4d+7b0/vvpKgmE5hDFnlpxNKm8JVr/eRbgp
VBCLPonZjfr9a9Q0Y8ch8YDFhg+2hoGIoyEsQBIFFC42T+7kd5XkT2EAL8vFmqQA
MtJCKiWLitQvtbWvYYCYhIXhSgF9GABz1OXCUe6BW7mRTwHwC9NQrM4vrrGejNBN
tlAxGtKSQsbrchAXtQaBGUHL74bmuNgukurCcuJyGOKuOGVQS+LxuhrwzEBZDY8h
98wOaCBxfMPsiEftyVhqm3VL6gMZF0eiBvHRWEvBR37WnQFL51J7ewMDDuvZp3ju
Bofxy7NZw/FtS+aoFOdrjLkS7Rup3sD5WgQLRiYIenQquGCxvm7QNWgl8DaUQSAt
exZawFivvExErzPKxKTpiRQxR/dVLSGX1feN61+jZm6SU+oka627PAnQeKan6yBO
oxr4+A0Cs28vu9BPfCnwUEALat2UzK2nDkv9LQfgE0zFvnVDQSdvwrVKOV+lmELA
ReqRP9qpARnMTnW+9/Ylsrm8bhhv/IL55Qvn1zVgkrSt/COv0sYbpTuuNNP+BMzZ
pVIPwYzOnQ+V14qzXio42lAE6lFEka32vioCYTYDmisCUmDeGJ1KYIJmDNLxeO4O
Outn8J2fsrBwFfIwkCqSkIMKfy/QrgnklxKspZia1Oan5CtwmTuvnXOcRWVGalnn
rnIR+8aN1FDkLY+jNr2TuSqb4kp6LXgr6YMFGgtR1TMsVqnBpqCtdpyhyqwviieA
1vFin84+/wXRAdBTMWrVbo0dy157oh6SwNjZMk7X2IP8yrTA+cH0mwhDoi3fRCDC
7kbV8BggzW4ilYgOwuTwkpBpgeZd1Klq30smf8sBOv9qZq3ghqpZqC67wetSDJ/G
682uWGQHGsg9dMaqeNPF3IxrmE+/6bZzynIIHj+kKfl9xdk5vyy23LBnmEr88kfE
HNkFdtfICfkelFu+Dyq1y4ED2R4ec/HaePP+01Aj8tP7cjMUyr3SbWpw/PCSiT2D
QEt00lW5iBt8nFoAR7CvCWZHlzHf9edpPDxHfh2WEBQxBG12yYbgaORoVdh4zOmb
Cn5dz2bQ3wY8aMt+B58U/JexfASwOwRYYYpeSaQX/2Ay17wOGS+RmCWGg3zgC3rg
Z0NB0IU4Z/HRbBwQGiMQKGrR4jIqP1lvq6gZ5B+nGY/ckB31CHu278HOdGbuji4V
XLA4uihdevD9sJfHe2DCx1/jETnNdRCpjVuM3xo50+LGt27Qs//BRc5T8sB1LLMt
yusMOZPTCwJc9Bww5W9GAQDJMeq+VPSZucn9QX9fqQ6lCdaqZ5IZm+CSdHpI13lQ
denJcH7m+a1qk9IDR0es/G3J/AyZjlusoTniKu9Os+tRtgidKAVxcPe/xA3JQ1wx
A5HyfEORPkwGzCwgtkMLdA/UYqJNSlS/YyI0YqO+mKaKANs7cPfzRMxCV5jdNQsn
2udKMJuQTWNkQ75Djfz5KpiyZcLhsVt0nWQHpG49L802T2tncdqQqbc2Deu+WJ5Y
jXzkRavao2KcO2B8kUH5jwO74hxB4e9matMLtiG0fUSFUJs2kX4pOIiwxvPF5M3a
lfUT8sJk17JTRiMyTpl8CFYjBzuaao8AT9md3FlAglPUaJWvWL75L71MYm8eTknj
2S1zRDjFhbVv8jAOU/MalvPQECMpJZbNrmYfdM4v7V6PwqvPWIgTZ3u6Jp1G3ID+
U0hTauslhpuPMZRggMWtluJZobt/PPY7BYuE/v99QK8zmwd00LPehFDAnu3O9nyj
MlpFJFn7j9KiSCvYTWhHN9EAHdquCa9NRNocSqePYYVDgydsVWulXM2NFrcTKlrV
n+oH1Q0FHBhSEbYtphcvuVIEXcQlrnTLdzUhdaiXn3dPQx2HOHrltu/v8qi8YwkJ
OnHxoYaOjMKY3yxo2MH2/rq08DA7CWyGNRGSI2JR/BVNFTu00kSAGC6Q9pifqM4J
pV32UeTgqjRsdIpkFFifCnhIxUMWqi+xBNC/b2gM4LvPMykmlLG2jA8wPwXxTPyX
VLbhn9rnugyutjQdBMV4t1LCRz3klW4H8wbhZ39FXVcjZFHNKPbRjIVhRCBp/moa
p7ecaIsiaavxRrrF5eCqhkA4lQlmnnz/v7MABygKusx25ikDe0qPGRMRasOchV/8
4NKb3XaYDVSHgj3i+G0DKY44CmrHb4CshdysOH4XUmkUPuR5PrdmJm314/jXSlxE
DjNkWhC2X5nbiXTfafFFDZZUFl++uG3HKuAnHq/K+DuHq/Fj/d/y/ubdphAuFCso
NUvOHKhA6N0kEFqyhJKf2xHWUsMzzsxm893GaY3RKgv384eLK+Gbe9y7oCPeooEf
1JM69cjTucFYWn42AQD99SQdT294Nz1CEIqSTWhboZNSIYcsRY4RxJ01cgnZZCIT
R65J3fzWVatzFAU72SXCiFah2eRxjvmxHavm/2egjvnqervuA4i4QczewweIplf3
c47aeBtroBaclv/k8w96cbs8dzOJndslPIb/nhCYvGVr0YZ8YmXPLEUPwOsANz0T
d+K171FCzWswXBh6RuQCEXYNid2JjQnxgT7inZcufbOqh4Ml6ii3HYFEw6E1zlZc
7OWwF+0VQlaHPxjeFcs6cHUbVEW03tXhuXjW+B9FiVKK1fqNc2lxMgvG1pGQVB9V
wwsAm1tq9BYoTQ+zEHozUBbb2RvYLlPLS1UZfQ/C5BgyG+YKJsWEVuPcz3NxA24I
1AgN+oGSTGE5ihvTJnJ2YiehygwNSw2EYlih/6PlnT06SOOQyzzGp4ed20Pjki7Q
4MvNVy4MN2pUUhQYmsKpuDNxWS1QIYXrR+F5vqLkaWNXil/fEQUyFW1mib9HXWL1
qtSc0ieC0U2+BJzEDk8n7sb0WQauSPn7SE1vWa92GZezhfmFcGGZ3bSXjLtRpgaP
ddc/AvjOzJVSFwRQuTgfcyblB4/lbY2fw6dJodeKZ5iB03AavToyfxUGnPkYM+HJ
WSwg4q4kA8TjxA+ABQ5fKQAE1/sG2aQ9OdgJRIj5bl5m56oRrfk6lRhRqHCbDr3a
TIwG8EX5K3kV0/u3wshiyTL6fgyreyeGJJyYlZZT0vKiedkn9W8djy+2USfEmGJg
MGFAqCHwO1fCNGduJ3uhJoEZL+tcqkByOARQausHMJDCw9Sx4ddJIzR273eRUczT
1uo20mvQgG3Mi1zXsxY/aSns/FkScqfi6slcCiopUoKuVfIu/CxsJ/wQseqdzpIn
0bGG47jKd/NkOWeUd3fG8QO+gNncS3IOzmIGHjr7uNHy+YPDsTZrhhEEJ8fQpzlh
tSEHONp2DiAD2r4TYUpHoVTjCAPikdscR4OncVV+j9pEuDgtt4Jv6RT8tAaRGcOZ
HcBKnDCn4fYQzc+d07CY9p0STBJM+W1YfVP8Qx8RCNY3dRxJ5K6wcQfT5z7XqTxD
9mUEnXDBkY4sA+M4HuvhUBB6xY1Wrp42VAiBem91yLRG8O2qsUiBxg8JdfePxpRU
oMg8Qd/bo/Kgn9pEaQdtDEWtPGusG5z3uMX359j3S5v4H+ijTTDm5Kr9NYcQyer6
aOwHESuNvtwaPRfcDNJxdl3hOk6XknoXBvO2plTxTNR3zZsdzYkRD4BPSRgnxnrz
u1S3nggHGt+jZcdGQSg+eFdxN1ILYOLHtJJBuUGSU4f5qSiHtwJVBm12qMe6up1b
5orsEpyNc2axws7v4oyZGjWVj77JsW51CZCzgniztGU7hbWG8K88f1RUVm3Wl/ak
p0nAPZELZ4TfCUQE3AOWL6LQouDROhiXsMVl/nrwsTlIoD0JlTutvEaaYsyZ3dgY
t2epNjWC3nvi91qDSn/BNMOG3P8/9T6CuujhQNXO+SahMbMDUHKnhZnXjVLXB//8
0Jk3uwW7g1CkFERkX8nu1JuSZli5Ad1o8FQlNn/9egqIbEX3XCxHQv4HAVuQdpyM
9E0UJt7+CuKTDPZhg2/hxv1CXvG4JjqmKynApHCTYNhrk3Z9wFdDRBPO92ioIr0Z
g0FftO/nHIFXF6/GWSNGf7247pamzZK9pa++LdPkfRUjycynRmzWzv7MJ39WhEGL
I4HGC+x8hWJdjVWzGiCDWEgAjDL/n5670drBeCSe4Iy0ReWMWbTeSB+FmD8QVn8P
oCcsuslRe8DErxoVFr9UrLbBPdg3+rVgzwYX+4GTB0qrRm/q3gh5lzDGtsKJ1Myb
JiyHmRf75S2JB5GlmRIJW5a7MuJcvXkyGqbULMYMK2tosHDE6k8aUMgl9YXwd7sr
1ADNtN6Dh728D0xYALFyRtWVVkqKDLrRwI+p1N49pDA00uZkIecYLhdJDczoZzCL
36+amZHK2bJbN6xo8D8OjkDa4BZQYHSBcd69pgVmCNkW3jZa1NjT/uufaAnu1ZTW
FbeabnRbdkcJNYU4CyfBLcOD1pX/AVrWwPv640N3Nu6/LUnMgBmVtCMKHArqGCta
MLVrITDJJ1PmwBFSWHIF8uf5ktetbIXZuYSHUCKio4K8U9biZjVrQwbvBJHReDHE
Ojvq+PWNVnbAZB3Hl8eOZWeqQBbwlFahmPDmQMOfIgs3Qi+/SzmvdvIv1seYJTRh
3UouGhimTWRw7DCWvxm5aO7ef5Rmo6f5zUs8LKi+Rbu4JIcyvvEz71f6KUAumPT3
6ZMvXedDvl4xD2u+QEtZVi++ZSPfaZkYAgHYI2FljsWKP/HwxocOMJ9I+oG+L2TE
y8t8Vws9Ngp9mI97hRsKKh/iiRSK5jzovqpzu7yGLyk5zIkuUpBF0q0E4uavfk/F
aYlvmaWz5O0kfan7T4urQHmgC4rxWPjCr6+upomrhUBfwNUsS91nhk86qoVesF5d
oMGec+blN5mEcma+Ant8+vUoKl+PPGtVy9uHZAdmrOuXSYlBg3YMabq5OKIOZ6C4
H+A6ry2Jt2hJ81K1ZY+dOThr//1CrMf68HpFZON5Mi42a6aYvBnzHZeueFvxzEtp
nd4lLq4Yvscewsi/syYIV42ETd96+K1GbEPRteZ2eYOc5gZQpzhxRqpSLB9qtpL9
VvL/FY9UlTXEIb0CHZaYFdEFO99X+YK04gugC9mxwKyGH4AGy/L9E38gM0Bh9YrZ
lsDGAxyN9At5Y3IdgTpyjLYtzWLVawA0RBAw7ZeZH2GrUHBuFlqOItJFc4RB8r2U
4kwUOvGWtk+lgKPTR7VDNan7nRcW5Dfi+cQkgBhwZM/2ZZ1Nxwopx62/G9uRTsAf
qYUnIt7j0Deg1xl1h8xTyxFpO40wQI0PUQfYE9NTlN+AfG55Kcb/tc0gJOLwrmGj
l0SDAD5KQe8ReU7zRKm0FJ48QNAVxCkIA8oPM473CKymB0l095RCZhH7osvybcqT
+A8q8c/TcBijKVCuCo/koJdRgmavK7RSnnrML4FGyC1RZ2qhOYlVhurt1wioo9A5
RSfR9mIS/XVVpCtqNp2FEdVhzwO6Je3sJ1n7aSYqYl+E11KMVm1Edq1h23BBXqOv
3NRi8hHxZBNhXGz1XzGwxAv/n4BTpRCWc6p9Xx4RhhtNruGrej4RdulrY+lBmeWw
OMVWiFPbAP67KGYP45f7xguJ7BrgslFPMgAwrjXPOTDI1TJWzWqq+Oi+rpyNXyNg
GwuGbJOhz1zHKmo+Db1zqLRl0BTdsMrcn0rTyKELmv7rdw7rma1bM0ISdCPSa5sE
qU9Evkq0YYdGKjWIL4ktHczCzzPCOwhOMN8aiNgC083lVnKlunhdtrop2UJzaUFi
qxZkSn1gQpWSRUMIASIibiRl5o0Mf0jz1eRxgLpGqGry6Tx8OYpzLvVcRTCC1fUy
VHUyA+C4FdVeyjah5Qjzz910BFSnxQixE02sVAQm9xaJmE2Fo/2ENn+AlMVzCk37
mrfpchHyfg2geEqD/kCMMEx9Ff6BH/+enMxT2ZigzDzsFBkQPOJLKGgixHHAJIiF
LzsoERcpzHSC5ei6CHtr/halgPa77cevNUx3889XKMmgdPns/aHdQHtk4+X2kYih
zf4Hx6ukkR4JEZVVbORKsVf7wn1y2i+Ka6+qJdWBCdLR2TfyOq+W618dHdoq8Fk8
Dwmv3qFQrAZDpWNuX28KQkWMdT4hVJxsQ4pLsOa1sTTLl/xqcjo6fmv3z70S/lr9
HxU+Mo6bpuNZI83St80nq40N2soS/j7ZsnofjovKCJ24KkFtHxaC9LfXepC2naYq
SvdJb5X2yoPdg0WBGjIAyYkVXPbowUFVxzAxiys3S6kKHS+urETiTv/g0Ypy+aQw
ZJjN3d7PyMFnPFIONRWNAHUVwK2yFT0AfyRY7SmloZ/Behej6quYGRqby+ImgPY6
y0O4juD1Fudd3YyBZPtb/uYAs1l3V9eHWUDupRiTLNF9NoFb44p0+RhQ1KM6PMne
s+1yF4xOoT+n+K9ezq3HwbhUqOdXH4/QpUT/XOkexCZ4KNF9Qj2/+1CJZ63Z2tv7
hPAFmH1D8C6DRwfQiTftq7IEGaXtbNomayq47p2G8Vvu8YLXWKbnJP7B2yl2DenA
OgMWsQtuzmhORszgFP6HPRVnveQCSvj9jo9VqNYTahMlcllVN90Fjj+gNhgY+G0q
gRdy9DzXcX53cLZxnArL6Pazxxe61WdhRqJ3vOcVgN3ChZWnXzHOb00qak0ymsFq
Sqafz5VmOeL10mpN9cclid9eeE+OZYuW/JkAmzVNasgaW8evWpaIv5nFmqpck9R2
iJv6qxj/LCgKoGUUdedYO1Hy2I9Jzmcy7MUwbRtPqmbgz3e7yZD3Q91KXPS7idRP
GYPg42V9YBlF9xA1HbV0E9PaDxiQc38Sx6jt3ZvqD7/Fr1HIHQy2kRYtUmZivKok
d7Ts5YaY69XhOcoVvGnVfzT0GbeCeYrrM54/jyhzzkgljC+3o05xhwXI/q7krvrM
KLCMfE2A3JSpxs1k0EtbOFK4X/DqXuF3ZwspO9mxxCiB5dqyzV7lWZCVW+VE269e
blGeezYENArIpWpPY007tvadMi3H6W/BdImDIscDwYfqWsAMYnCJ3BxLdEZ0Qr6C
qwjchFnY4Fiu+RGwGZPdvdmQXs33EM/YTO+e6o9Eetsd6zJi0bT+DbuP74TeyZXt
UUYq/1ehyVjcyU6LVxLJBixfjCYvuuaYN2uLwKD0loQ+noFMXO5sObufUqSdRS+C
WT46qp4UuK+FpR7QqIbhg+qC7JKVwJtNhWG7nHYhZMVpY3ZIffEVmcY4WVy8hsNK
+6QQR4RQD9Nqy4GtTEBvUUVL5vpv/M1qz2kcgx0uon7H0VTuGvkrc0gfSpXN2Cpr
z6acQQsE+FUitOGKPU+fFh/oNhuSX/cgOsnwS/WgiXSWsV3mGhinr7rPUu/QoXWD
cYU5yxdpE4VKXZWMTt9tS/riKNreo77Bv0KvYx1mURrILa9ZAjOGe0V2R3Bcow3V
YqwKUwudswaDJ4D6fmdJ7EVyQyjGD9qRHVC/G4U1I4UYwbrpP/9U4j4VJKoMwY/F
5GrSDQZwiq/fIqKnTzn5+Mn9hPI/hG5blVE+qk4iBKu3IzRyYNjIYMIGJvAIJI98
fcY8ER884TZuUb1j0xCM47eJr6X/7GQHxwYu13SdrKFOWwOw9Hk406zw1uf9zk3F
0wpkGScv8w5fhjRreRXHKfmNhJq4sVfHi8oLbFDOTeKPsQz01VCRbPv5t+u4yf3u
tsq18IgpmVc3na7gVBOu/z0QtJUph4N3rU5dUcBLfVu1Xevf0gm3K+vhqKM+C3MS
MlKgvf4WfuuLq0BKCqOjFXyItBXHK64BKXhCFKnuvzi3fRjwQAfT0S8p4RB75cdJ
bzlEo56NFnaVKUR6jNGDDb/wSYc7omaX8QbOhWmPsmRFhx+4G6UdJVtlAZc72dpc
8mk0LCFnibOiGNKQ0qI/AFClDdrME8tIi1CsFbUFTF2Zo4bnI+tlErkZ6XMNUp7u
6g0EoFdyVmQbHk6XcoBYbR6VDETekW7wFbEz1oCEECZhVabTIGi1OQJsX86kNryY
a6T6V/i4XQOxoerl6BvlSXe7TabDTIGzXL3bCbpPz+38cb42C7VmSkaGkmyxZcE3
KjPSZQ5sesqSeJwDme8vze9NPruhXbipChtB2BBaV7C+JZXVkJC8bxUSd4o+LhFi
Qcb9XmOoyTCvI18C2MTvjEhTdpCPRCgjrsYbPbkrVD1494+5Q1s2kkk/L9u8bLgE
PUKekHp/WVcQlx8waDKEoEP7SB25HHOnZcHF6kfOp2k2VAP3jsfUF8eVX3QGELxf
zw3ZZ7XDlaeZIudUQht84dlov6ldQWoiFQMrcwcd+ej5cvf6nGqFjkq5vdB0aWZ/
XzdVy1bSf2zZ6psUkah7Rb1+06SBhe5oe4gG/cEI23KfAOzPOHxTk6S7FH3Qfz1C
T0xeyB8ldx4HxWLQOaon14fWDFhMh6RQU7+cAMEaJ81SELpbg9pR3gYr0+R4gqnT
qSabwaGUEwYIDJZXJ7TEYzyEYRo4ic07dGNb48td1OE+jCESTYif0/bBaCQ0/Hyg
jtSdcATVJXWPx4/1gQsoPk+LWv5nSdNck8EU6aMFZ89B0rOVzTK1xc5gDaaNNg3m
yt/UTDwa1/pnX9gQruu1TKNwDBIr89ui16TcwE/CJ+eZwoWeDsJ4pDLCDTrXlmwm
KVKAMwXsOOEq0SDujje6FKBXAyGsm52mgvWd3lrO8ItvX31NAb9WWSKUhqilbLEW
//1BxyiuDcH/wOdjxXCan3OhSuqzURJXDixz4IGAijGC4SGWFh611zyM452+arv8
lJNPeHWSCqptVy7AAOAbzOnGWlopewDR0MZZsjvUpeYwmelVHjtWomOmG9kyl72T
dpF+qiBDgkrKFFGd3rLwU2nJhrUvDdgKa4knBJH0Aag8BAgjiVR44M2WdyeqPS90
fkk4MDPlxXcxzfYNX/2CGdKsrjCA0z5f1bh3BSiE2gNBexymZbWje9l4iJq458Ye
Myg+xBL/SKnpCntyBHJESY5CT4NI7f8MyFRB9IrNxQQb8OJH/Fi8tE/3TxGggo7J
zxi5XR0ocxQuHJBFrbjLeLvFv9QYBIC8in0/tMoSM4vMM5XcPNbkykd+FgJLQSjc
arQki//ayDHXJxNKddX190qYQjCDl/TVMBo3vNOEmJhnywiPuLn2N64eEbGss7ML
bv3hY8I9BVUfXQ9YAJQ/4F0AJjFm73BkK3RM/QN02d+xdb9lJqti2lj8iXkQPAsU
7D6Gatp3Y5yqtXxLMGxWrMLiH+IhBPsQgxw/SkeKuVkExf2kchpc1f1XVXPLfiaq
q1vuNfqiHrSKwnAMPmtXh8JlVCew+xjuLHtesGSgq+a+54mWRjoVR5h18kRHxzCq
W0r7W7Vg6xbVoQuWBSGBgCvm8pPyeOlgyIZrsYy7TrRKzHHYAH94rv4ji983J2kJ
HKFBS7tYMMwYSJwsC44Ho16J4bAw6XL7AFCM52LO76F1qOSsNzFPujvzohKc+oLv
ymaEUTRjK8ZsWJ/N00CrgxNmNmt2tQt23K792lxLZbyfVidGB1SdjI2wuBcjmwmF
q0hQvTQFh7PzSD0TCacERxgtC85+NEjSjdHvUHXhZGUDR9to1Sfc3rfZze+rGsxd
C6zXYQILCll+C0USRJUClhet0Pycdygw8aviSswEiJQPZDsHKxvYwBl6scGLit5u
sd6N9LI3d+Cjk8Uvkiio2O6HJJ2/EGRydmrtdxZmYku72vZStACvG2k1wTgGAC0H
ER3oEimFzf7os84G8hm73kqyDxEMy6nkITrCG/pHiMpQyVF7eQpc+uTbhQjtOIaN
EsDkawq3y7t60xEAa3djN7lATszRz2Dv2zHk7In5lQHWLaRKOy7kkVb39Z94Dn9u
l5vLsxexN2ko4Wp1oUuB8q5CQWn9OkwWQ51DTQt4qNY01IZGnqjfJijfryTDyF3+
HHyaBGaUWvGyMqniAF6yGNYPDTJI6mqHQBgJFOJLSZ3Qt0fhal56cikvKCR9IUAT
TE9jHI0H6jDJuXz+tbokCXHV8tZssBzA/e01pFH857VPuEoWHnqyXhMjcX1ISR7V
IPDJ0AmTae5Pt0UzqiXo0kpFLL8LEOnMbxk/Jeu3qbmZ0j8VSLHINUXASG8m/A0s
2xB03PwwN/1zCaWIvqOund4fBtzAzZCBOB64YPgbC/ZfFcE0Dbu5EXD3ca8lZS63
s9BNpieVRmqrQwo/FixeoI4fdBcZpplgm35me/F+7GEv8LJMmgDS9KxH+pV36KNQ
eS//Cxf3wFUbsgYG+H5vNEFzlnAPxeA/4Sye3qu59crdE12mWpChQpN8vqOKjwgi
pFZwfrDsq4FRbZDn/KilDRXeFEZ5KAVi0xn2GeiVc6mrj56EHIwBMhoxlq8GfNq3
8s03mB+1ur2a4q4aXMJE3eUfj/lhFF8yO9wUZihGCd4t3q0ikqeevDUC3HHqZSWL
WI3kDOQVk8PeBYedKPUXcuPyiPx3NnrmjP8uZtjRY6bkfVWzlZPcMwZ/W5xia1R8
vAcvDIC/GSZPY+BoMdRyqJENgxnJRBFz79O7eNicqRh181GQy3M9R26+Poc5iC3V
UMdfh74n3fc3Bk1VhjZtl6ymGnXUzsS8MvYjIJyV0dYBC147BJm2CvOCoPmMA9wr
MMxvBKkHYoGWah5IvGZl3ltU0E6hFBO5HYqhlZ/8Sz9QBcXpV19MjpAESmIYluq9
uol2KgqeRyUGTCvuAgoyltYspOv9yMdgPivJdZEc+jdbKdFsv9SjepV0cj+ug1gt
SoueApZT25Gq8cGXZTWBM93XaloxJhNIQlIv4U0COoaECjNLjQy+4eJG0UmobYG9
2eBXsJta9jVBjxQhX7+0cazSZkFraxrNfm0sGAEmIFm4u0gXku2sJ74UrVMuxHRW
vhv1fVEthxuOCP2fjn6Iq2vSJgUVo1L65zsrHeAdw4fZ2NBhObYm2rwjMJTG/rM0
G8Mtt37bnF79ILQMVSpfK4VIvy8C6up9MoBpHaiiBsToPv3cb6dyE33eEmEHfw8U
NlkWDOrwxHUy+di0vf+FUtFKcAr53scs+1Vbg0k2+cJv19V3d1Gaz552cl9ZZN9m
B6TlXkDVyk1sbNA27+b1pFm/AIVvn+Cz0iUwuKyLDnmPTOe43Hfa8E+/xra2c4CY
XaUC/mBfSnjp16WQXOCDGK0iPQtYEywPt50lMqeXN7x+X2a/DVKjccePT/TBvyFr
0IUaNVZz4iYoRGYF2ywR4jxK5pRBfMw75bfVffiiC59ndlkcmVXWZIRkCG2SYB2i
yozgNHPzRl1I2fSkymbgO3+SCmzllA/kFkGefJOYoF/gTJOoylN4DJw/ArLDhZUg
dKtS+ie7NgYXwZud2tjnl6Is8pRrvckK06xYxO3YBav/R9J3ie6pcjsG8B5cIMfP
yRPuY8ib4V4KdUzeeyjm/iqH4HA0TWI+jaYeJATivmVhw6p/PSMfNnvsx+QgPq5X
qyDj/8HFSSMDIuNuXpColfzFfRMBNIRmu9/eTFIV/Nqcpd6bTsx3VQaaNp1qdDMi
9RQbry63zbk/TCUBLBBclIurpvccSAmNUcV416KB+nElHB5xHE26slAhS2AZb2fl
Dpfn22ulWzD1oEEPa00cQw5WmM1GVuBf2F/Dej4tqn75rHPbTuy3cvLHU18o8gJ+
Ihj/ks7qoHKrZc69+Pl414JeGZO4UviorQ7lKlQscMqbDPFUxoR5jabliybhcYqz
liA2lxDQmLRkf+4D7RQp82570o91Wk8xu/AaeyYYrPOAVv7j/mT2snNhQRZLIqql
P24iNmZ9Gggibe9a1r+mgZAH8ZoxZDN/kKOOR8MMw+DsBpacUxFfDoEQJYREEu3y
DJuwiwNXHPdDdEwDhDLk9mTrMCjsNsJetvgkHqCkQDwAHO4M8NLZvmzNBLb+dgYT
uoj887AIUEXN7DTPVuZp87cKT0k4QvNW4wppXb23++NZaizWIYmCks9yNTYoU+Eb
/0ECPteLpoG2Etxz3MdE10/nCmeVEbKaifyap8zjgMMOI1393goHDJNNy6QVM/Aa
qX3lkXNx46yH8ON5Hb1n2CVArpvDsAkKxR1nv3hXE52fxGKcJw/3P17h+q5JfpRl
/OCVQiAFhAxCndLBAsBLQ8rwc6FQw2kp97ad7Hl8Vu3e5Qjsn+qKb5+r5Fe1WtJX
iB8R6ftSkKSFfkFOtwsz9CCOYzCKVzzzTOzephjkyH64jb0XZnYMDJ960WcZeY8Z
a0PqocbdUbKgRbT35pjCrMeDmtR7asmEB+Od9OEJVFLkfMfCDal5FwdFah7m56My
8ZdzMXu+tcfcJJxxsV6thdQDGFB7X/EhDwNINT3MX4bz0tZqRlxIeZ7r7Nx1QD7S
sNyRdjqFFei0enzxfoafZET8lvKzt2dU6a5CUv7a99V1N8CaSLC5co0R25KzEN+5
eDNRoPoXjWmS0LqCwqC791ds0a4vAgRsQl8FvpBnZ0wwfhKN9F7M63siN8XPGf1L
vc1lV9NlEzWvRbK67iZI6dJi7nT6NBwn6is3G6cSAUrst47O84hJG5LApu9Jmfai
Wy92sUVQvs75c8nH4MkYM7wPS0+CkA9+VZnqeM3iO/MdTYeVBSkZkezOu2bBkNAs
DhqxGFZ8KqnTgrJsqF2SlqJFyY+M6CEGAnAjGNgcgVdm3QQ4uygHIDY70fumCoRd
ibUk30T6vd14ri114a9mC6BGAVZxDPm+XviZq8GKZV032UFYbhBxETNqlYZhwwr8
O4M0z5QvecHT0pD9nhWG6AHzF2BmZM0p7fIo+mhkOCXqbsTPO/IT/cawsa1v3p4U
Ao4NYqr7m2pIhK5yfMHlun8KTeMpZ3OUNYQMaVFY5zyjtK9xLtQF+HfGUPzZgEdT
xneO9DDeDjy7AyUpoVYJrKNdtgatxKCI+QiXBOGXvvIKcHT4kYdJ6Op6T6W9zvE/
6HiQB8cAO5r1S1i3kIERn29JBCz4We73BlUuh4+60hPY3wKeVP1xNSL/fq8ryRPE
GRCjkebWGcgcC6T16mCfoRl1Akdzk9DaTTNq46XIp5Cv599xM8V9OoHZQCCTQ0e5
LnaUpRtyH17S3XlrEF5ktbzkGMXOk5eyTkZXjdk/xIitsbWUiLjhYgiMfVQBeKy1
t4aXz8AYhMRnkOS5FVO4/YrOcsu4elxQks9hDDEkFL+AITwYWK40F2y5MEbEayUK
GITN0Iaca50yhZAvdspIOFNtwDExletwnF8I4vwc2fBP+1JNf3dqXBJ7aDXQRGeU
66XXwOaf0AAesK6OQpVrrTXo43DealkgFwd8aWkUlttR9bf1CS+ClsrioOXfulJ1
4MVo9ulT28RYpeX9VugvE/ZFVu7R0tSIvLqiS/rXAgm/ctT8pDKlgc3OCh4IH3/r
zxnV47LSAqaDBW6vxlkRVeOTrIQohtEtuAKZlCVBanKBYSTBE2Ku8zOJxmKCRxqP
2CQFBfO9fE5yv050h2Vi+KsuAqDaU1nz0t8Px4GAUq+uU/squ9D5RzDmD2gn4nDd
pXAuJ1ZT5c7LWLbFisDl8NJ/lv5GurI5l7fSITBK1xmSayXoP902ZmMqICMavxlp
4LO2+1U7KCp/SOuAMa21Rb+4CogLW5D32Yj8gMB/2rPyHphF6cGCc6cErHN5/ejK
E5t5Gd0RdB4vIDiPv8inmLX1vQoQGFOEVwg6ZFpZCQqMrLt/CuwkZnNXSezGFHMb
A3W84Z8d8DTVUI9lSimp/l1oV/f6qnquacNCRSFTFbsVraFzvrv5jUIhwqLTiBjK
GHOgZNQ2GVsexIbvw7ErHfjYAAWD3TRhGVgzvRDEGt55h8a0L8j92tYiBTTFgXfk
V72YR3Fx2J7rVlqDFRAzKhzNZn9EX3fX3/QYN1z6Z1rKwr3EZjXmaVK/f+9wvylD
jN1Mu2cgMEKbi1sAZF/YRgWF+Tbk3XtPWr2Y5aOtxFvTLZVIb2OkXH4bs7X88EUq
JWi70xZ5nkcXfVCFUXUkRAbBILh6dZ/VSeDaTivT5WPu1rxgI9h/Iv+pGbG8eG8j
4fHRqZFe6VQeATVqZlaDorQOSxGmwYJ3dcrI4AmqD9X9Xjk6WjqmQY+lngkwubKC
TAm4p7CMkg3l5Bxh27qU3Fwa9sH5ly6iAMZ9WfGam3VaXRTbZXQTI9RBPNtw0kL1
2Gg8Zsz7QnOUMqs05Y/L5FcPuuudI8rfIP9XHL9DQcrjMuqvQq0g+vPAwFRAYXjV
Au8uXVd9ex7YIWaqH3LOBOIVlhbZWObLRKswNC+T0qakgQy6tedYN+AIUtJgGy6M
mb4QwJNHnd2/C1Ero/FNPRmLEpKpY9+CkeD0e0OZZDtGIcV1TLOrbf/OxVEa8t/T
BN7q/OlkE3TayPO2ZmwZJ0yILTB6r5NMBVQXrB4c0C+LYYNMWrpNJgYyEwqN1Pzf
gGf2DVRZBAbQ7PvdGz5UiZ1YpZPcs36SFo+sJ4XKSAAuqGGbNZugh71QRa5GpJZX
3fr8mkNW8O/syPkrwHINNzcb2UwX4+SSF2buSqSHPYOUnU6nylY5yj676WkTqgw4
8L5jeVGpgCMrCPal42gOfFf0orXNgwLmoeA/WfS6n3joKa2bEhPOmRjBjj6Qr4dk
sVcMqFvI2uv1sf+EHKp/vLhrFeFPuxq2GH1cJDE1ihnchLkBBMSAbLiE+1dvI7Gk
ADBBufd7NMYpjgJihnGXByhM6YlkpOOuVY7N0cG+WYYVkIrytmKk+KQQyRf2vifN
7ZxxZ8Q9nrzYhAWkpVNGiIHkwdJ5tGHUZ/7VT5NrTT4QD3pPd4UyuxKEZvbXu7jP
QU6TgtNdFy6YLXGvTxs7vI0LeIj6XD0QlNOMDxW+Qyeitx8ghsRXFPFuibIH7D7D
ZX8OwV1O9bom7qWwEYbHI3DdtD/5QdGNwDyR7QOVY7lDfM7AbuXOcWe1nWS8JqTZ
WLv7UiZr52CRuAZNVArf97fe8kDdq23aPIALbkgONQsRdjljei4aQaue6kwZRWQv
utmUReq0+aByt1BGIBWXW23mG2YSWfIZklK5xHGcPBxt3erW2ychz968LoIW0uui
eabp1mrHKKnhQ218RiIrmIdoEKp6OOpyN+k/ToZbC5lnJsdCHyy+KDZauOUBTb7M
gV40zGZZODuiYJhd2H5emd0Yhrnswt0AYOASNytI8uFX/tz9UTkAA2LaqKXY7ckk
/CXH8VaQ6vUCt7bjEUUK217XA3l6s0dLOzkctlXSdqOtMa5je+uiO8O7UFzB9Hmi
Zj6QuPlWUOgI8cnARtbcb8IdfpHimgmIiRfjG7U9fxUyQ2dD9LDvcwGprkCA/k7X
uEQyZ1KGCM//4gje/4qDY1sEyTA67YfP2ed1aYAB3DyGLSQaA5iWj+mPaE5yxBmQ
qIwDuj+ygZKr5sV/v7FBTUo3+66H8vp/U8cINDYL7Gb2ehAaWJqqaH6qO7SCSAt8
4xF7TUeQMAKW/sFI/17LS05aKD9oLP3qEDhcJL0VYQLcGjh6OIOqVA0P74bPMNxT
q36xtHHn954WOs8xmg+dxBlHv/Va60ZTshvff7Igprwap9NtnBqcYdj3TdU/rf/T
7X0UhT6oc4anW7t3OD535GHss8ErIlVIQfvqKxEw+ShwYghLgRbdliTnOnBPBiLj
qCItUbShHwmC+JZWgzRHK0Fy2ShkukVNW4TrUFRsbFYmV2GCTaZBbbVo3n6pOo/y
yfO3cFuXDVtNeJ4/9cJe83yUTf4BOUSUF9S+jat9uOopdIkDHNozZiY8fj1dcNTq
6snD+46W0HLi88aDD1UOLOPiL8kaERXN2vKPDyvxj/HYEhpHG1ZKb8OmPXnLor9S
FG4IlplhV5KdTM3E9C/Vq+Xgxcxb8mcY+NBOTokNl+/0FuIAIjWVrLjUmk0qyFb8
frGpU1jrI2MsdSZydTvVCeru0cIa1utw2iIDS4QiWa7+hkSe7bRgjho+QmuPYGcw
8iZPaC9PvhoWee5GPeANUIK6ZhJww0eXo9GqImMfcOUH7Uxlps7eATv1IhbkhIhS
aHHYaLpefze0YFNWohwg9SnhxiJGKNW+aYhXtzzuMsBYr38xYdRaqIBNzpufl39m
UfZ0CS1GncOXHRoLTxwR1kRW5uqdV6TbWpDNslUOLbooFElFKt72/0EjSR64FGLx
3hFzMpK1Ak+7CqDA/Ez0c59lSvvuznFqytsoSg6cyIoMRpJZjf00wluekK72dpd1
XdtezJr5SftYIcq2BZFBNm+pv7RbDvjRFMtsI/H1fZl/nKdA/ZpSmxD5+0AYuyqD
iTu8d8/iKr92TFhipshkhC4rz0yE0osiy+/mSCEsL5gJnZePNhby4vLw2pRhNznT
lMjO0FltubeFZBpKrAEfq5hBoIuxn5EERcp1sxG+/AvidKMMsBdFZAnV55uem7W6
INaWBiITco/wLZrcU6SN7PXUEqx6X50nyfyHVyyW/MrSlxL+I9+V+fEMD8WNX0MO
sIIupPajd8hs5oxR4TiYErocnEAhURUTF76v3QFEml66cjXJFt2Yno/ghOQA73YP
dRPNwwnvFEHrUdTw7lFaHFC9f3IaMnL4j3vbqHK0wbN2Xtzzkh4ICinVRCbFiY8l
/OAyKdL7cr/FWnT9EMwaoPB/XxRKfCDlhXW0RhTxnBvVID6wlIM41HNTADiK39qH
jZGd2AHygrPqr+rh8My9BRwIMlPBK+79ExpmlCTKrvKZy0hy/N0+tiWVBB+rjb81
UR9THdFUfePmnESD1tiAl1JU57MChMVM9Zb0E6tQhiNdip95CwKdztTsGHXXtT+i
fIh4/cEoOst1Ayft9XgDNUIKFMgJg+miDvgSMIGfWWL7if5uBp7/Ki8fVYaAUIuC
eFKzTHpoFfzcZpE+c6Fcz/vqClRd9z/+RzDGEn/Ueigh++ROnywfXCtz/DjtaFII
Iug3D/RI5gTvTDTUkv1BSBa4li1/a1DMDI5S5OGHaNvSRRgahs+7EX0/bhfBD1KP
iJwS6kCPH0ZGwVEhX1QCrbUulZwl9ru/SKw8dYG6pFoMIDm6EA98Gj91fr91cBEg
QUI96YAO2I68mO3aPq8bbD5QZpM9jJikj1IB3DSZSBEWaep/hsqmNjpl+nm1V0nf
fIvYr67m5tYeAS5QS93oowy7UHh8jkluQAKTj0T3gkBSxCP6biYtrkYPrAZVxfec
nOSlSo305hPULiSQ4Z4m7xOTQkoeGAnwP54Ey5jAYP3TVnDI38cJeBM2tX3BRAwz
MlVpC+EwvHzGpjqw0V9isiffGsV7iph+duyzsyHkwPuw1k5URIjfXDADsERlrBgZ
X2DcL/FsTZkdLkCwcGxkV30U/BFyQXKyaCQfmsNjdZS3igzcMgsM8KNuof7hovVC
u6O1nhViB3GuPerUN9AMybfwx3apq7TDYHLqgLjmMqicM3xX4doFkeclw7MURioR
Z7w5+ZP9yB7ysX/zGk4gWrqg+OO+LQeWktWb/BufcsY6cCbIkSx2ytPlwSjcdtii
VBn3Q1em7bz1e62MtWOV/V3r5DS/kbOnUGOue4T8Rj70xJvQrsz6MT+umeCybAyX
hIbfK7LsC7J5dJ4NYggltSnt0lKblPI/lIqK2FRZcroURCvtxgiQYEYOmc/hR5+f
El+WBURjzk7+big25sAa737hSwKOrn8QemB0ywujw1WoTFkED59olxnREG1UtGbc
qVN+KrFf2qZ5gQ6r4pTjMr/z+foolbWuTvt7HyYysRsN5wyPcJ6kHW3Ggzaw25it
MHlzUXAmh+8vR1seVIyV60pX8+D9a49eRR5HARxbXAG55TqeudGmqqjRud2jhkEc
yDBpUPKtIQC0WwMIBCao0pO3PtEZBjDFAjDVt52fgZZlDeLddxN/KM9KAJBmGm3l
JcD7BBELhcjUQRiqy+Iuri3m1dV0HDR0rcPW9aB00VLi+fsTV2ssl18M8Y7Md1nx
m97WQstJhpiQxewheRMAKHvg14EIrE0I5Zse2Ab7PWNTnIbNJe1Tm0VTQQuAF5tV
LtOhcbS7Om0Cv6l9L6WulwBvI0sh2q5fFHrUpalOgMZ0N7zr6KNd2I7/+977UoNW
Gsd1yDmummAQrC/x0yAxphpWv6C8L2bEZWjA9BFO7wER5fnTGYeqzSkPwxxsN4AP
ArdV5jLt7jYQ99YLP8VDCAXNYh5rGLAOjo6zM0b38fgvGxd2Gg0076mG9cNZvViS
7vL4TJ9AWac6vbxU6VZG34Sbj9sPlh3q2pLTjBGjWQzVTKDKY9cLp24R/fDxudB/
W8+tvBMWwJzUOIGNW1H8voAogldjQuxZtn3AwmjWO2p2xRIo9XAmf8KDjU3n97k2
ppLM8Dv6mIdWXyFjO4j9hMyAT/Fo5bcWmGa2mK2IAfpWXFKon8F1zOiU9NQnzseE
JMwAcTRF26Gf2aB++t6nabKCCTHxTcxu0Q/+zUy118dKszOKJayEIg/pW3lipor4
jqe4txQtOVZPFzf5eM6FWVroID56Xlc9irvLJr2xQp4fvgSF/1fZlAmoKjl6L6/F
Ri24H2EPPV4taSg/kyEvb/FwgNgCjMnNiMBdAed51o0npSZnH1w73Tbbse+pNIIB
IBAMIml4QbnuoipBxznCHqkwga56JHdyIljlF8/ujrdG9xjhk9E0lSaCoHkHSsHW
WMq5RAz+axHe0NwzmzdqhRnVs+V7Hvkp1VNAJr3hZg9WGQ5+QTK9yB4drPZK8JiX
3XS8CqIzL050cISNYNil1oxdlPbdzg3Jo0FZmk2xM0Aq6EiwV/3J5zcIwpBLZnmg
+rxFJo+s1jiFX1ppIn9sfB7Rb4gYWW1cfaZ/bsMzKN+4Yx7KD/ckylUL6gbEkpSp
2MtQGK2fnT707pqYCeabPM172+4xCzpxzZFtgOcag5ZbqKT5cWBT3E4CB+U4BzE3
gGfY6M0eXvkPZUZKfD894d0vAdGY94mzX9X1Bs18JToLCj9YWXpd3i5/SGR7YgLP
7UGGWrk4P+Gdxr2mAeTtesN8w+84/gWnH375mNApdJD6TeUG1EF+BJ9YDQUEZYYR
toc4rYt+3ifZx3jMMmvg1jfsOc3IZcoRtenN5wOFc5x2FQOPanZCSB5E5eX7eDKI
LNRof2JQcR5RpCiqd4L1Z9cST5k/sSQMy3F4HAPb6CfXEEnphmLVqAitO2Yx17QF
0U5f55kfX4GNCwVy36TkU89RMpF7Aaz06t6k0J9ix9nt3/XZeGJJRS/mIT55XVyt
Pyz4kzWs2Q1PcPBf0Iz3iM4j1FPwsu5M+NasrqBBiEPRfhMh/fsDg7xMvsXH3dl9
3Q9TuEA2fpWhddZPZgRTIlSsV8+7rh6ZHHCVTkTB7AvwxAOcnkbJkdwjLp8VYdDN
LW2S4F7+mEilBUKDQd0hVB5RxFh9JzCvEM6e6TGzC+qlPoZS8gdSJT5y7qetZWYo
29jm+X88k0cqtjd0cH0DQkHE0UbCoELlibmgIqG3DhTm5UAdgudFnPVuFga2AVzl
D+cG3OQbmR87DZ+uIqC9+xYhQm2PniEfidVh1UDFJdygeES1m/o0T+0BCttfjgNw
94gqWxEckHN7YmSLJvSc+RkWHeQ5K0WEd+dnOQ/KVHJ5eZnFw8CfFN6kPMTGO4p5
X3lo6ww4nypf1hJItEj55eAzQ3BTjQBGIHQF6fPBjVMeuHij+XyWleCQJwYs9uki
FB0rb7Qv0r6yQEKLFU9FzAM0iJIlKmRx65bXRPtsUOx8DwqRcsrgBie1TOCwKAxR
KYMkIouw0etj11b1WAqYqgUp/y7d23uJDrex1p9fz+XS9msH9J7OLQItGcnQLfUp
ngO9oYZdl4Jr36ujhG/j1JDAi6fMceBTOWrQg8dX7SqnfAyyRUvFYiQYTxtQ5IdZ
m0/93C0ZewZW8Iw88GY1XFlUSFBb7O9mnlcsWu7jg4L7/7VnEYGJUG1LwWpZ+Z7v
XQn1ighqdzF9yU2hUOHjkdsb3cqtAZ/IsXfwnI9XHv8RRRDc19oey1QENlQ9yneP
fQC4LicFl77qQrW2Xd6OqmmtU66eBkFCglgZhIjYnGzAqeqar/8W8Gv6gBfHqvT3
D2vD0UzVkGo9z9YXuHoRAKXSHrAlcAM5o69x/i+c5hQ9vq/EuvV5QUKdMd3axnG6
bHqRQ3PQEdpQBYKwf9CjPK66hw1ag4xqYHqdokaZVE8zWPuHFeACBgL6alSOUZrz
z5pWn3RxjnR+6qdnrdd+fPrSSj+5OCHkmhOp416tUtoftveVzn4sO0MTO48SfAK1
isRlh6jtltA75DKW0XqMk94w8et5ZvmfDnivy8J/4W5Mte2IqoddvOCAOg20EX2t
F6sBBkoLXLMYVNv5wkIpgQsoQygV32qlgwQPM9KdfNO42G8G42/44pmwnuYC1YZZ
vRBSIQkhfukXuV6zAvI67t3l/lX4bxw7U3GdDzI11RRtWqOMCqJoH76CtdoQ2RVn
P0XgRs2Xbr/73NfXSSgNPvoQLzBOKcYqRFNyz18UtW+d7cVifPiXHxXwwxnXjdrx
ZQsz2KzkvvePZR7xlP+vadf06EfdOG7xoiqXDL9PW/f6v4bdpoG8QcKAjq73lnV8
iCPFzbn02oYdPFl0iONt990dP03AWqAC60Jhq3H/jUx1/CLYWZI94ZOa6puDV1zP
K6pkoL74yKZOey6l25CnuppCJ3r7y1nZFkFJR3gq0MunTJ2OZdbjZWRFhnmbf9WW
RtgcN2LEecdjPqvreZfQsZOq/sCbvsOXD9hkO51VrrYRf0xv9dsLR2NieiqLWnNI
4psQdvlckP1Jk1yfa5ZVLsIfrdFkkW8WscYVMfbdrF2QKj9uCuQ8xFSrzK+egi3l
yTm2Gm2emB4mIS+QQmtMpOTGgHxFQJM1eJ5/lLLazynAZx0OisdQ5xJyMsbNayr7
f71frcbEL81SU/iPYUd6L5ArFpUN6GS9RXw4+1LfZEs5N/dCn0GiPcA9TfxwALrb
erbaRulEFClw5zRoEBMR82yT2l5C1b3EMnfNrQWOfupVhJx2IO4XY9mxLxjaLP0Z
Ot+lVqODQLQMP5bsV3km0xlrkhB6Hh/Zmf4BYegkWV89fCeHtnSUpfW7LQD63RJh
RIjeajKOOEHVTFLntMMeS0kCuGi74HIGU6hjj7KZq0sskvAJHiZAHohoYrJwcN57
8f1rl0JoodlRQoOrRbLHQR+FH68i8lnWfo/RUGh4rgl/hHpOKjDducpSUfupk3Rt
RrIVpXj99yQvkiCskOVxtimuBODE0s+orFkiEMr/veUFP+eNglGJeya6CMGcunUt
v65+Ey1KESnkL50Ggc8Wr/CoDaINBbHyz8ZyiOY1ymD1JTrWmFm8G8/LA4sQE9a0
Oh1mNd0AMMpYqWacql6VA/DRubd+Udq2xz0X9XxiyXd483R1DsNyPJWZKatHXwcI
zNx9A7tkxDOQOwJ4/JyKQZsqWtPGjkNEKsdEPkCldvkqGVVRK0KyRIoLD/xTNFE6
UKLdTB0UdcNF5QNscfsLDxajCQeP4JaoCFSNM4qh1OsIC3SiEG1qEDo+0R1KfQD7
/4AzQRMBPwwwcv1f6TxZNi9xF+DiXuh3XpdNl7g+er9wgtRK4jgt33m8yqZQhm+K
yn9mRRB0s1W1WM8D7xlDXPI0taRBRpsgjQpTKqw2mfYBGOz8ABHfonvGs9xV0aCm
rgI38amRS6zTt4dFcFnbn1yFifnp5xP1Fjs4jGYIOjO4s/tmvFvLn8ogyxvbkGFv
ZAZHHdOH47gZ4XV8FLTy/XXI7AMA+SNAzxDcAXIKVczhYqtS51nyPvoNv56jHSto
DieTonUnbjszb8VhO/cx545u1rvTIFZmG2GEiNidGOZn4XmeP2YhxOxkskxbW73/
3xtpGaMhmHIgVIbrPOd/r3VhJhaLGQQIX9mv2Hv8W1Je0k5Kg6WHhXko7Q2J4tsN
gKLxymCiKFk9x9aKYIex5LvsyMIwNGqGGgelh/pVkoEhWfmL3EDMvkd8Vaaa+ErP
VYMYN0ueuRoPKUtTI3u1yDGMFi+Qk78m3W584sqKiCplAv/MAoK6bDS8SOYAHSXO
Mzm77ebKaKYE/9s97vL0Xyr6UKa5ayZs+q58ePz1hI0PfOOO4ZKQPNbZf2zvdjRy
LUHgOMAJJi3B4Zj6Taaefg0lseFHmZAdpQgCcM/tWepxAc0SWtSkHOU/8rpCBEho
KO4UPPOH2fbWtSAxZlsoinFkolP3rDFb0W7LfxL7WgsiXFlHAXGDZUe4WZEs7O5O
HGAWCPW8w3Q02cj/6v5UG98eG/g7VXyo6pOClsEYg7oNWukTa/wUB0GSj2eDq6e5
2S9q+JEYG//fAiV0T3xrKKHqgTopLtbf3T6icRTPU9SeEzYfPihtQhWsOJwcuCdG
RYuvP3odFBaiXHPtNyHKLIl1+OjPRjfNxeKQDxtiCaMAFIvQIFdb5Szf7u3BLjVZ
EiO2/YxdUhyzRREaapgy0OPnaKwmnu6ENio83Mtk4VzpapUcgZ6T7MwDvhMwlm6P
BFHefwT2nGApYlVg7bjNbPmBxrPm+8ffKMgnmE3Sg+DPZG990dJllvbeKbLAe/Ew
HryazvC5r5qszi2eQ6JAzLCYMvyexJXSd/ui63sj+HTG/fiGihaBZ9c2wvFMmCB5
SEA6we/ttaEHj7BZRwCW0bSBqL8RhbIQClSLH7n4apNfeESQ/I30eGnl9QfAUrU2
nBdcbQr2iceaGJR9DF6+GuJrjV910axBjDCfvdsS7ALijxzdTLbbhFtuDAU9Z77f
uJguZ/wfigk4mhCqEv3olcyAjeYaQp+V12HKDMCDWj2rmWOtk6BvN8cFT+c71xpD
c7bToXfEMKinjRv/pmmoBNeWjJ4jfSDeztEAcZvyCb5Zwpe6hXik/NjziTekkIXC
hrIVJb2HmR70ow2gis5dHuly5javl7iipYdw2wOb0Qyiu5fWn/eRJdAMlabeWj3t
OrGedmSqw8p7kT+cH3/bRfFkeZsuUoITGFBAUexMk/4/MGVIpU5fEttP7SjRGWvV
jbFESxtHqqnG98vVmaAYb/X4u4G4iHPyAzmhOQriyOR6SfD+gEDStzzDWzxrcq13
kYMKYCmzUBMD6WaCrIyOhpq+VyK+L3PWAdkYLTrmxNfTscU8lZiOtqTRBO86GfnH
gpaH7jDkUy65hLBCdMZa0azQxekTFyYjonMQjD98E/IzELID7Slqe/ghNenlRgwE
4032oCqYohUUine1Hfw791w1bFhCDrb5dy+0y33PVimTTRVOiWYhIWjclVcrJY17
A2B/qiizbbIytZYE/uJwSyamUgyOVUufEjE4OLXtoz4IGTi/ugwAqH/1kp7/Gq5q
JNXP5kqWOpfR9oIfhVTLM2YjtiQ8O2iRShRdZe7jqj4/+Z8lUbZ99FIGHfaMq1pl
ArPAv3nHJPQwv7QAoVl7HwxUUTKpI5QU/8379JGR2lNtnWMopJl39t+zkIrr4lCE
5Z/pcaYvp0ylinTwp44i6TVTwkxhDjpWVRnHW/GToiua+dWkYk06z96xR92OfqAx
dLdxZzj5+V3s3G8Kr/ImUzaYW0yyg/oJ3R5dc8tbqcdbvm/t0kA56PRr5BZWRSjJ
p4KSZxFwAVCv9zowhB/eYRMZkDJao8YXQosUIJJEY6iDIIQr7a3dDKCNxDAZwanM
19Am4kdu29S4Ppa4UM21qhnVNZZZozNuKopEySZ5kgG088eMwstQxFrewO93FrWt
Z92sbefyIKl4Mi4jic2KWYQOYAUs8jX7ChgnRR+bFJEMOg5JUBjaKFkcaeeWTkgo
US0cQwTFXkU0Twx8vo1r8OPKRrMz3ZpFZ64NLft2mWJ9WjEE35RwHbg4CNg1F87e
v6fi4lMjXKydugIxZx6FM0/ONZx7hOdJhSkDLRtnKKcDKHKyvDsDG0MqML0rN3lq
a+9YlX5QHd4MZ5tlDe4kWmv8YXFBIQ314BoW7ChHf1OWpKQS8RKcE2C9HXmI644O
jjPWMK3fln6+csE0MTddpZIvI9P1XxqrZ92jtHgVg/Akv+VkNVGG6peE3Ncqt3pF
qHJhxSM2raHCHde4or4CDlUjUdUUCVEWLv19Vezr7D8NkfjZcm1y6gdKT5QVfS07
rNtV8l3LehIzuLVTTETIRolJVDiXy6gtAFvo9oe27ljv0hCyR0hz+1AmnGYDLLiu
42ieXmlBbuOFQC7g5Pbsf2rjC0FvMSfxDtz6sExw0qgtkSaT+DbnDFZnSVGgl+p3
gCtn2/7BTzd0m3VCgRxtu/gmVgdOXohLghJ8iIXMLMOSUat5etfHAKnCUukAVO+j
li8SL0btBr03JZS0vqLOkMHhLNc6PQ2rmav2L+GO0paQAOYpIobCcXz7fPWand+1
7ZkibAje4T0BJ7NwhSSOtVO4FmrgCVQRXDmlK4wlAosYa73Js7jldN63D2S1ebB8
SCpLInj0UbxhxOyNJ4h1VGLAtd3PTQquNashZZbRkD5PoyLVfTWdauV2oiEfTbBT
NFnaAJBxVlx0g9T4plJ9U1eI9q+09UE3zc3ZtQ+Vt7cMBL2VAs+6C7gAFFhBAX7I
JO1WFFGSpKlnFlEt19abuIUZK+nVHHFoXvlBaZLuwS/gj16aJzD/V2sUQp/63iO3
J1rq5+vHcCD0AlgTF+WPEWNmWCOjc5hoWtGWUsG+K0O0TGKIP0tNFLuvt/0Kt8Ue
g594sZrUwkvHJ2/g8plF++PoXdXI7I0nN3wU/rZWeto/5oIASgLvtkcNhZS2NtA+
MGKjhwBvYfA6jZfRbpt4USm994Qa6LrKgzLSEUQGCuRfn02ZyOjAtUJxgTWjdcJr
3wYKD2CrmIgR1wmPOsaP2AbW+pQw7G06PXDXZIbnKXPMAXPs2sgMG/4mwte5id6Z
hqTrPwgMWWtSXYjBV1eFwO7GlaxPPDX2/yyv1VREL/TdnurwqG2XDSen0mqJjLdD
jLxHNMKX4C9v/lYkeOhL8nyWJeYouQ/TIbzyqgIHANVRA1YLQlaoSV10qifzhZkl
hSjL/dUbOEd1nQDJNtKFMhU6yPdYEo0TfIX1IK9W9uyo/vmdpiTFeOBePkxaqjGP
PN/R5UnvlzUJwjJlcmeMeUNM5CPOHmF69ivzQ72HX1BTmiPLONkRwaPz9bsH27vz
3iT5lcvrhHMb35HDMxNEya58iq9afz+BpbjlcAJkS4RJmypo34fj8tiDguPd5ivj
eaZqcWsMf1MOSd4O6YepFpWgHnyT5EyugA3WzmUQp/kbamDVD/SS+sqlquV8whcB
S1wSJiSOxjO4ExGoMnKie+wKNnFkN3rjFgHmek1sGgaPrid7y9Pq+DILxNm/yIOJ
/2MHIsu8Z7mmy6d5aFdG8wK/CS42uU3Hk4W/hIUdNU7aZNLnLUF5otUX80ugIFiE
+3QxU2YYwyti+YkaOY29ESZ9dzaVEbZL7cVQIij/TgVeHyvFX8rvhN6B7qbtO3Ne
CMGjv8ZLFxIymurSuFLp8NeHpY7iQAySgRwYpslBggtN+PmcXunywlbHn+xcx4Ej
knw46jAs5y4gYIk8czr3JBY+Q4qBNycBIOzHPnNmtB7Rt5vcJ2mkmENJTsJoO3RD
NR7YEefwl/3m94XSb0pRD9JkX2zGsmLWwaGsXB2ll5vkGK8ligMuFxCtZJmEPTEu
+kg/gaF+j+Nm+smv8nLvsM2gaonwG6eudEkEOsq5C757vKxhz0SWkK4wyDE3S5ly
qztfRSzGL0kNPPnr1ksrurokVlhLOeuw1ptXt/0fpm5JsE7jXZANn1ntZw5O1U0Y
q7hRxA/srdV/ZMY0Z5a5z6sFsj1h+DyJsnlSGwoZrwVyBNqZd/qTtxPELxwQ/eSD
2DFIL2nRUnQUc2iem8wgL7reCQifvcHkF3spMsJblrl3fTJa+naOSwaGn0IXBzpf
bvgMLjuMKXz81nsatbB5Rh9attqeCbC/3/Ru7kWj1fkdAoY4SHvFfcWdqTdTE5Sx
6FZksVCabfpAYw8iuher0spr6VuzLuCwjy+INZ+H8sr1fBV8RMqcUy2X+sQRo1Il
PNntwC0cjd+SIkiSjEA7+FLXQOPU2B+Jq+kp/PHFPqtKyN6ljNSy2JcTFUV981D+
ugX4Y6KKnjntE8iBr1OYu+qVxivjpkbgJlGUq/A4Fo9jycoMFRABmFcauY1Svprs
iRrl4B2JaQJ48McctbkFwKxeaKwfOwVKA4IBfANhjn0iRkY+4Yi0RMxqpZAunbAr
ys31W31TbHGy8YhsDl/zSRuRkxIHj+gy8PUNsoWr3PQrywbge+SBH9vM0nMSJ12h
viBomu9rNRe+W5Vnr9OP5S0GCSGqGkpsDRodxjUxtIoJB8qTaP/aLZUJTvWPEpEI
2qGhZo4mSJr8iT1WJYnkqexGbosKb0E/E4cZMBhaJ8Mma9+MMTN3hDT276MuqG8V
+WanfyeSudpYxy9pSk8bITs7euOn0nCdp97crUKa6ZJDg+h2BoTsOh9bl6HM3wdr
LTvhBpOyT68QkDfGXl1DG23JoG0kpwXuHeXMIGJE24fcceWSpN71fJMkU4meip+O
PdCAOeWmzm4t3swGZ5LziWfRIcP3PBEpyVh0eJgxVpf1XtGsw7loAvYYQrVvRVlq
2QdhyYe7a626qMgi90C8CM2P5snkjD09AsSOZaB6DXtj1L27U4/7M6UXeWEHbSB/
BTlwlZzZBBSEcJbpH+sUJRwx5/izKpxn1mnn+v30ykL7kzfDfWn3BZp9sQOxmE4E
Bo98fPas8Zv3i6BIdtlQCV6Tkg7vQxCUB0K+4hLqbvw7KHBmYnp5voG1YFq+RSUU
fmHDyhYxAF+E47vqGXuwpR9K9vS1Q1MSP4Ux7EvJXy/pMIgTQI8vAlDvDye+2mo5
a6TXMLOS97sH8hF059ZtPaVJ73avf5pfuaVQ+3lhM4tTgJ6vreovSZvWPtVZ/PTC
yTDjuup/s6RlO795ri+cbVeLaAPtNfKSrWVDG66IX9b8M0EP6AHs3N1gq0CT0RIV
TacwT2M/1nPbMPFIcHP1Zv7H18K21k/qjFlCmFV0TpHjlGosVXRiztpEfV3EJOFN
IFDi/oUQDBCxKvHIBCnCKhMGOvWgZd3eZY4C+JM9tgHVisB/T4mod9tD+gYIrr4D
HUoKcGsH0d4whnemtnnWp6YByi37VgiTw/HuzzW5ojM5k52OA9kIlvxjX0xPKzi8
XBfgTqNd+uDZ4lMHSsbUM8JAw/VSoImgyysVXmPdENtemD8HdKa+RWV72X9TCpi2
OW5kNwNSOZvzyIMwgAJI838+KUChklVAIEviDLJwJ0PyvBDWT0oPUDYVJjeH00HY
IwrwhkzNJPe+6tILKF0nsJGBH8W/FfWsJzmzZUA6+v633T4sB7h7kRPxVYGcS3dA
R6g8N2zisatNcMSihk3CcfJxYKk7knxqXUjWw/PghRhaAk0yWyds/NQAKBcyLXWj
WG5ySij63zo/M0vgPdMg0GmK4OJqHrrMg8pdWTFbtpz49V/bW+RhOyY8AJteJZcf
CL/fYS1GNtgOPrBWIMqFpxOGT1YQeAxJbKzogAlq9ssMGBnlf1qIBbUmcSECiENT
JkIcXLDZxeHJsOYOerTJY+DhwNtVVlx/wOvyMT+wZZ6o3c5S8n9HR2jWBD6EewCW
GTrxf370CvLcpxB3dChnOFoRUJlAW9unos4VRbGO1o2J4ZCav1qJRK14PkTVxF34
QbfsP0mCLEvkMhurIGRXE05ywH1k2KeYz3BAseTxAgg4tB34XVT9GtwQzEocH7hh
5h7iKFU6K41Qt/qVHdBwFcR87e1rFJQuddeYpDuP18XPb8CtNvvwaqEL+0CR7LTG
9ynFBN7UPiiOQOWBNATevNLy5hc8+z09DfkfxHqKN2UEqW/4cYTEy3MJPeuDjYDF
ucXQmTc7E1SWRdyEehUB69eQDuOe38uD+AtxGChRAU2RAkCeHUK9ChGwSCuUFOry
eTXjxX4ShL7NSF2Xa5xKA4Op5Us5MlOl3+RHKj0VHfCZoxlzicJPZ/GBh4R9EzvA
wZv0hteS3xpvwN+2D2dKnZ0+y1K6m458JDa7wTfOaDzQn1A+ooM/qOS7n2O3lAW4
gWxcsmnImwIbK6SEzNCJhglzf40OhsKNMsQfGjb2LpEXPupDhecoy9En2HbniaLW
eNQLjRxSfWKG6ZAXKnpZiVOPeEN0z5XBUM8njJGaLUElWBliMuVKs6MmFzyZ96Tf
inovTj3wsDKrrW6YjIIu7mwKoQNLBI8U0bTf0Xhyndj8f6sY0Wd+FfBCX5JNy4Q1
uRQl9Ma7A21TzaVQs2lR/zK+znP5PiCzJNevrZSKv5ggKlPK8z73abgurtoG8WeV
ymox/LxBRa7gJ3EJN+7IOIl5vphRB5l1H/7/R72qbrW2Jv0MvBd7Rcphh7YMnCrM
p2BRSdeGP3s6Dhe+zn4ASY5OyQDFTWbUrj8w61muhkvHFMVA/OQ/h3tHtPHCVAWt
hWrBVTvaT+2lQ1UCKhRPPF+STBpTGhC/UuY0tpBDX+vkhyZYXXXQ5wVWs5KAHKEH
eqmM5ifCs+nUT2YRqdcZaY+CQ/dShmdI7CE/HGriKULM1Y3Qxq/SXsrNnqNuh9Xy
56V2WFL7a3hhcZH9/q79KVD1raHNLrOqQ9f3qHwZ30E3Qbd1o9VrlOSyoW4MtQzR
GUI/xRlV6ve64NqYFwFDYK3m7VEIWcj9DxcmUAzfYQjVLBM0RqxL+SNTjPTFNovi
aQaXGlm93FmMDq3CibydiVi9gHkCupnPOD35ru8RJHKW1XrmpZzvOiYEh1pr9I6B
wLoXf8DFfe9n5BgEWgbzLVDv5pqjd+w0WjfMMgJN63kYRgWyQpffJFXXmGxcET1C
/NPfs367AZjMQqMYPuV3z6c9o14LZDToD+PyxyUXTMK4p4xwFfHKUH4Y6ipJaO32
b6U4lQYQ//nvUu201gFeoSDbEZNwB4RipIEEHLZUq+dTFCqke8kxH75oh0U7lmaP
WESBenX4Jgrf1OCb/wbPP1AQl8E49jxIL+m7FnM5l5gjwBdb5asGG151OOs5gzoe
939d64w5B54BQnaaSn2HifDZJrzzDUkA/cVLG9NkPyPanbwhZ6FSc2M+PvVhK9E8
BN2ALHEsW9jKtrSRXWj6f6aTr6a7qhZgYQLy3aap9PD+DDLhHjxA8z0Hyh3mo5zZ
AcI3WATjMKPEdnJoyIDxtJrJXsZGVLyG+GRFXu6JDs3DqGB9DHxl21X1a2kFQN1d
nBiZFor7dVyeGx0KQZDzO0go3yBREPxWEExMlh8nAaofGvnfO4OF0RAMao9Trn61
kJnc9DkVGVi4MEKdZTMIBmxQxliNcstrUGPyMYv42L11md9cBuUPgCKKGEX8LTT/
zGw4Vw7y8Fl21l23D+lTta3MojchmD5UESXL2Np/vFd8YxwmnLYhkzx0OcL5KZcC
hEd6slbjGmtaM45IfSOeI13TRR9+PCdJtLuzXvFo8qrZzsJHJUyDmt5IYEhECodC
vW9MZNsEfoczQeWP+UPoS3yQse7nnGrT7KfBkuPDlm4jhge9yRWBNgOBrpeJbnJJ
V7U0O69GMXBAyIfiGMhwizvLJnpN+FUvUO8MS0kVCvwCrCP9vBNTHz0YCo4FNWQg
lQoj6z21v7crJ5PCzLHoYiqmEmMwhm89fl6w9tjHTLTTZ8KbCU501Iz0L2DZWxH0
HvQUZAPJj3pa5Hv/RwjdoFgnMhGg2+9IL6lm/EkBG5swjQJ9zzUP+4icZMjSB5E2
k8dnQ929TngdzPRxzW9ClZqHC800YKXhEnIhw53fKOXXfHBbkXMW06Rk7PqQD3gl
Aq60Kr4ffc9FgPJrMNj7cvWujNngC3xpwoDYbHKKc690oA7ovW6+RsqmR/xMjbS2
3rFnkobolFJ5FTSKyTwZR+jmaunLJHj8uLqld7ZnJJ0J5UJlX2NX3aP3kRoOSxYn
ftKZ0S2LFC0jDsyZuKYWMijFEgVq5d16GoE77H6RxUUGNRjrfSrCXjT1FJkNWCYt
m/cvXqLpDjGRK6JJ9JH6CjvFiSzPO2hFYgzSdL5+cjdXvy9s2aMQXdkE5afl/z0V
tHXnHSIF5ld+Pk9g2gyRwFVT+repoyfpsL+mshBoALMcjvHlp3tT11OAwz5CB9+K
EtOfYktk/b8rRztZeQcM5xUVkys/iys1uCLlV44ohf40RhwHZpCA3uzB2fBTq6c5
tXMkbJE5/JV/u4wawb/hUGCalhsezk7WBDNySoK/qn6hbYIrtlpcH4FE2SaTZnxn
HvgiU1JTaW4yxJfCkhqa5MAWQgORfi1VqWnqz8946ByLW2CCgsePr38PXAcRPeQY
U0qyd7Ttj+uAIOgfnTUFMZ0imG/S60m3NJXEerzAGYEO9biSLo1ORNWnX5DkFySp
vDZrnY/WxoiSQachXduW/y3diBtBxtjnchwaBDySfpdWJFdHvfhJVV46dCNMuTty
wwYjxv3Uuz2xngrCFqk5T4ieYETTjs3kQBB3LziDPUZnhrRCDzvhwHzwcp1KAg/i
w1oF1C06QAHMOodk03PX7d7wsZNyxnbICLO++a6xN7C7QkU14ifzUD3c3OPHBRmU
ydcGBE58D3l3d3/Zk7ljBMCazdkF+uQQhVmYGAJWu69OgW42DsMqk8EgbGEYE1c7
KI2oT+kwB7t3nCxlc5SCI7NYIneoM54lqZrTP6PmLz09NKqUk2vl9p5QQ5Sl9iD/
MPO4NgY2+5UfbuS9wkXhZq8iGnBZn+YAmPRBk88pwRHnrQFD/3iM8z/NIkKI1Zl9
gDNguPxOb9eTPQrBLBOQi5xAmpqfqItdMAASJeerMB/KRC9+YvWLqqw/z61kMW2t
IZI/taP0r+xYTI+lNceQDh3zQrG7lw/sPPknwAooBIor+/dWM2kbWReVEhNaV+5T
9kLmsqMA5QVd8zuzZPmKO+o/tkRc3zC6nfuqQ6RBfFsxZUtx3Nn5xAhIetPCw4Rv
dy3uBb7xpofEGvbhdICH3YyZQejahwQS0Dnpzwjj20gdurqHfGs+oEV2nfOI61qn
kVv68vCW6fkdbw0mOWW/KjVYtkvEsQ8uY0W3ciKhoG/5H6UyXJxBcZGOCMNXxiNB
Np/dKnATUEJokb8J6GvgIFTLkkpF6wszcbr+9boptFwEIQ4x3/3jvOwwwm1yK/Me
EmvnIxlWCKJZTsiJPH77B5Melg7jZgQmBgl+faZE/FOp02lXuV7dIgy95r1kxdl3
lfG5/FmOJ7+Vx5XoXraPEjfsmhNy23usbD5rAIPuRfS2TrrmlGzxs09qFdJ6C20S
osc071m/wXMLmVAitSDVykGrmUGiwmP3Fbnm6llyEpy+IQn8D9I+2GTvQdpSRjgE
iKdoFQaN/eIe7ytFcG4BCdX8H+/00ii3IpJBNSlO41Z5K0GpoX0ID+Y5QJozl0ax
0RHtFOjcx0JLZCqHlhXB8JCAcyHXXp5h5mjOTWoCjz1hjQWWwkZzBfXhfffbRGXF
Kkw15BDo5rVsYO7Wrz8BpXSyJZVAvQRDZb49eV9qwZIKw08YvvVSOWjoJkTJQV7z
ys5UBBmwYRaBetqPmWfAQTvbN2JVp95q4yXFgI2DE30BCP5aWvQVymPUNKZ4RpS0
K7QisZ1xduoV2A4Cz4aCp/H88GD/BeeholNvQuIruJ+M0G97ZAm8rRxsj5jPCCve
xFdRO4fzDRx8mfHDJgdPCsqs/b3d4TL+ZGnoC4Sq5L3y5kC9407rAqyzwnXAfyEZ
XAhdTVrB8sZU/n/sTlMWg79bN5c9KSXfXCsJCpxRg9NNlIX88JRSHOlQbi9u36U3
f+wHwdEaEwsQuXBV1bMuzl8DI4NUpnl/GjZJDIbUDNiW6vmeRV+HDHpxyex6aA3P
f3leQwRlDLz+zL6ifV7eqcU1Qs0HB01y2rBFoJ35ZcNefsgYpXXNrvjrlzZQ7TpY
t/vgtPGvq1QJdSSyHRD/yS39txsMQUGmyPwmjI+VJeuvqQDDTXOXQ6ZXw4XWGlNj
RxCE98ZEPBehCmUOnNPZsIXoNBbhDJ6tu8eRN9nBGl0zaBXB3z8m6lBQtlChXcb4
8RDpO04Yw/6mw6VtrkGptLh544ws5B89yJE9sfHW0GbbLFx0CGMcoDAbMeDlgfx9
X6043kBKM4pbyOvRaG4MHUCgFb0W58uAhr7s64hjL50PWslrw8zjyUuPuoFbJMi2
xonfEDFdf/T8VwN8mgXvhlVp+Qrnv2xw5KxNW1t85yk6uSHyRC6U7JSmmdzlQp1X
bq5VNPBOMQ7VR3Mcl2Bxkkr2iE0tSNfTFX9a5d7INMLjbCVyQ5zdt0og1O6S7r6X
Gm/MKDclaRlyqILH6OvCdumnB+00qAYDls3UFnKdbmCRlYotOlnnfNLQzibqg4az
TBGBwpnf0PTBr+vLQjcT0COD0AgGs5lqLVMHaemk5wRQoGEoaFjlS7xpii4yZkRX
F9o7JjmSnggiHcvoaqq1xBTTY3kkzagKyp/M/v7V9GBrX8LMmJD3xMftW9kn3tnW
wEl7IJncOtBkaSp6EB3qpWQYD75Fxows5KcCcDHTipXh9qc+Iup7rgmPCm1nQLDl
BJf3hUsV6S5sDz6QNOald41MGkbteSvR4v6d9gBlOtmasPVnG3euD7J4oyyfB1P4
FVJFqhcNnkOvX1ySVfRB/uL7NN7XXtQMmMCIdjbOFQV88zWM9qzhO4ItC4djZhMm
hxBCpQBhK1j2TkqhG39H1sgNv8lVy5o+UDPi3bEiDkxATb5eOI1quLGyH/whDvUb
EYUxvE0f1YbJinL2wRTKQXlSIEJXYobJ0Wy2ixrXtjkHQ95pj5VDzxOI5O/7lqAH
uZR5h64RvYq11OjP+5er+zYa9KARWQ+1rifRQTQa9YnkyrxlQs5NWVfLlsBj4M1a
9EiJCGsX7iWvM1b+vrRmvsbXd9XIYvfAZL56AATRItgzimkiCtnzKuezsd0q1fPS
Pw/XxbO7GirN3pLL8+XrkOX3zDV0Tk4b61MGG+PyEOwgQhhuDbBqXoeWYLSQUUa1
SK8PNs+J28LnypjshfLQE0btE0Z61BeeamXjUYeZq42oiBt3wZ+N8q/DT2VRI8nz
NPmZtI0+Uf5JnOPrw/J9nWTYfcakByN49L+3RXkus6tvOBvlQSeckpe/xMIkI2Sr
VcvHtBclJ6t2FJY+7Sf1ONN79SPEhLttc2j5ExhAGNMwYrWHaiVFpuxAp/GIy9Bf
aO18rGwm4DRVCDV5BlqyC00l0E6A64plYOUP/n1dFxI0GbjakdIiDJMwqGz7vsnh
BstLRQbmRU4HyoB355Py7IqOL8hFhym5JBcNLQ8UQjchACUIcp+mE59gxjB4qa8n
dvHd3YvxI2vRHGPkENziFP2/U5PNwKHajaawU9Cbs11tSBv0R8xp2mgXCKEozLs3
b7pU9THJmk6rrGyMmGJ2RrWai1yXgNKmDf+6s8vJ/15vUzgFSRexoPNAFXI5uA0f
+Q0TKiSmjTF0AD4JcUzGVEI0E41DNxqHcuazyTMtQ1CL5b57uOV3oHoYwf8zmPFt
maVaRkm/l96jGCwocXvXVJ3odA6QNiKT3Oo61xH2IH9ZRBGDkLciSellXwYt0Ku1
9dNOKDQXQUUPwlxlgcqL5s0aYQaDgUJl84+044VKSaJVzkVUiJidf5B5bfISW4AJ
CpRwlBv6B+24TxwOTvx590KPG7v0dUi0dkaf37ASBrzwBwzSk8T7moXqhv3IbRvC
RpTrkLr5Z/rMjwOWztHvZu3mW3B48nFwe/ogEANumZFcfHUI4jiXqh8GchKk/5hR
eUSJduwRCSNshvyQn2Ek6RK0V3n41NWchm9+WufafCP0wFptwpbaM4zDGffHOrvq
INxMXBnNWWiIF8Kn2TOIeVmDp4Oden0701fUUJgCLk4i0Fj2iXCZxhpQUfifEB93
o054VLHMj2XUNyqXLIrYO840R/ekRhqMU5M77ZWtXO2YdsUzucQQLQtUNmSJqy5k
yWiXXDEkoBAr45wYnypjY3NNtu8SCPzglidgfLc9v9bQHA5+59wKyUaMUHcxQ7bK
naxWe0SnMt9US755Te4Bi4t4xIjOnEeSKc5YwwWHDge1hiZe2JgG7gs1RJpAfrKI
qBdoqclnpk7GMLMN+kuNPFHMPju7ZNiaxSr9D2KH62M9Lp/d61/iU+HGsS1z5qSl
hCIYK4vBPeuH+16ezx5LCYtjFUO01zexnMI5EtPRInbiL+NJynVlN/X+ZJ6bNd3k
OPir2xMkRYITWeUIrKJE6tquC+LJS/PEY0DjmsFse9iNNxACD+9onh/9kyMvh/tP
38ESLy4yY+LN3S0BRwbiySg3vVKjDROSgZfu2lN7Msagdn22hKeOc9xsd7erTpm3
w2mrGaj+m0b8Z84w+U+4jueUcKer0YkWwkOV4LzPXnzkv5oq0IPg/g1XTDnPsRB5
OZi2nL0Tt0Vo6g+D7Gnf0yLIXLYfsmAdK0XpANKZl3UL3WOJe4sPBPpXG1YZSmkK
gGwe/JA0UZh/LGIV3MeEy9T/W+oJNtIIBmg3loGLBm+6Z/pklx77BRJG1CxMqNpR
aa+78lADDQiyOvXTe1bWJZOyO+K5cdKZxY0ztc49uRJbqGdeEHyT02axnT3dZ1H1
eE2WIkP1VIk41C+TrfC5dXiFkQiV2KkVYJAANBzJNe+oGySRZcdLwCuvR/dtPTdJ
VYuJwibRyuqDu1QUckBUaHd5514ux56zekpJSMwl3Z8/gCa6KGc8HL/1ezB2fy8m
t/4cbQNH+ACEnK0DLF2UBrBtHR1Ax3SrA88PLq/jJyhyyEFAdfMed9vBp/tiTA4L
pgrFMmHa6mwpJ2KkqwW8xA1C0WGHIaC+RR6NUZ++tmqH5EvquU5u10Ekzqg3tePY
v80IUGf1mA2jsn+7y5Uqf1/0J3XczjUvpId7L+wsMI8OTvfEouIMWXLhZkeY6L9p
PQLGobUm68ORspQKmjTLTXVqg2IzhQphVyuTv7HQiZzxW4gXKF1acclQpZulxg3V
jOU97r3GS+EutJNMomHf9hg8gAXHbcWzGyLJW3Q730kj/7WqHmMh4VFxvTPug0Nu
1MLq2U9IFfC/EdoeTRgcylYttk6C5ufpuZKOe5gLfYxG9Wir5q4cYbwlwkX4irFm
hlFqIZE9wRXimFZCFw8eTKZvVUrj+BhXhtPdUPZjSMNrDU1DBw7MMdp8Sw+S4nMP
hrmS0t9FgfJa/FRgx1y7ZR22TXOLqPkBHQd63pNOtsCHKjpG9F0kfZifT8sx9qVG
qvcebeGPldRUjthXgrjtHOGHOPHNYcle4ETyqlANwIcWucgb5NwMWMNFleq6cNuH
l6LzWguBlze3RePDSS+d5dU3Wrpsv1kSn4M2Yl5IrF1fY8mF7g8WAlyzX9bGDB7/
dI6zuhnVQnz7MVTNj3UpA685n47P7vuDdnjJNUnJIed/JB82S6Mk0CSsZov2RJW2
qOM+TNsghJ3UwbQoNSFpUqGfMZ1e4tMHSNyHEfDxb35FYsV+Y00ramlkHwVgrNKG
qODBW65FvHa81oklt9s+7ECqrKaHBqEq3ph5uNBhl+osnnrz/+ip1DzU5+uy/c9h
DlQrnacmHe+WV/hQOQXfin2PzRgzgjg+W4NnKX3E1lzWFD7P+q/olaeBiit7HJM5
t+51dvKJcaIdjQS5dINlZewmuEaaSGBvTQpzHcHF3YkiWmjaoiJjXEtQrMmGDP5s
K2rZckQY+2bKsezcztnwPOzcGYPIjtyjN7eiOmhqYtOH+cNPU8wCcYKH2DphJSkQ
upU+3rIxLw4Fy1pQLM24LCb9vJXDqn3vCPTJ/SB5Egll/ZsIDWoQaoOD+d8LRoLp
y18ZnOfaJfHS9J5sJsjzHzXm6Jt4gJ1qLXt8ttTHITRA1Oa/p3MowST1asAt5GeK
q1SdYoHacXRy+0A5jY3VfKgsyI5uCo3CkcoIFE3s4T8codPDcAOLFD4u1tcHlhOX
usx4XoaREg+S3EMQR3UIQH5YslEwsp/k/DPaUnuGyABnTshMXObp9xttcMMq8Jzq
fKkH90udmmoKX5jYD8vP7JclSto/tl1R9FqAMB40sxS+WyHAn8Wc271J+EMsvjjp
krjnQnXReo7w1o5zvGWiuPuiCEDaQlg4eOOXFVGUk69xUdnkRSCBHBNF4WeIxqKN
VuvOH0lE9uSRsFkYL02F23HMT8J+l1NTAEUdb5C+OJM9Ge4Xk3wlzkMXjQ9eoYig
dfjLgRXDq0jqQtHyEai6vuvy2XmDiEGtorcyU3GVSHtnfS/gqV41ry79MskBDoy7
naX5j1vOE+vHCh5tJolHuCvjdNaOL9erLqg4qat3Dg7q2fCOX6EwQ4Ymwg8jUnJ8
j46zcUV8AqfxiRlx0zF9uM5PIEJBlNmYBBD2Bh0+7xF3v8E2UgSIbIQ9QCZZfM8v
eC0MDatu1ZkHiETj2N/TN3zl3RdrcSO8/dNURJpp9YR2oMavR1Fvs/HEyi5eAvNF
KURAQPSt/gu7Lgy3w4gyXoxQVWcwFJC+JbRe9iMz89nssxB7uMlCvIyS+Bxo74Yx
r6xKC2bmO8XNmq6sng+2MN3mX2hZPlpFZA/fwHIWoo8KTleIXCZQBfDtAXtfLMKd
HoTAOUbmK5If/7sUKp9TTK27D5uEbDm6kU7A0YEEDIX18LdPYhKNIspp04rYTq6Y
r4CStzoItT9i1QfLC7YzUkioLS9VUeQzYkVSJ+aRn4chC+lC02W/ZE3LyzPkl3Mi
Ji/ngrNXD9Mc2rl3VJw3aDdSvJdeaFw/rb7Eq+LekhycPu5nXZXCn1Gfu9xpY3di
szFbZ25troNJH+1TfqG8XaqhzIHI6imcHyLPixc2tFk3uTLn8RtpXdH8uxXFQf9s
/zz4kNyH2MmVhAHuJ3OFD5aQG2GwsLpbJn0TloyB0bWg6U74cPJyPgYfS/YHqaYm
wocrLVJzOyx41TJnwePTkE7cpqy8vUlghIVSAC8lHxx/IiGyTwlTle535Mxh2HTo
fKpw70mfSmqlXWDYFat+McaCB1kv89D1swEhPpKK1GqKUtojBeN2SGkJ0mme4Sw3
oMqXtaV/UzJDxMULogrwkWuysds0bJlZB3jUXSGbYo7ccL/J7DgdxR+OHfXg/4A8
q2J92rJZwnNIliZ3LjKRTFGS5aqpigZBCw+hVRxMxURCoH+W1H7Oqx9eL7IGa2ur
2LNZoxi8Gl0wrmvvkCz1wvMaklKVy8IpmSxIAQnrkfMf7Q6PsKWPo++xaBSufDWu
YDYEso3vJepIZq064IqwXiXVnHSPQpd17Hz+w7+WCY3McAaQbES3zILKiocHdOum
mNelMHWz8WZJVBmXqzOMos7vxr5tbvoQPht4E6RUeH51AfElcw1ls7/W02B4UR+o
foSeybuXWwszUKN1fQ8dHyao4E3dE6JSHdqCL3br8C6IpwM1bv8agU629ksJdBRp
9jZKLBFRL4RDUogOC1vCafDyef9BH60VUKmid/HtqiWXMHelnQK8UKGRIJrj/Z6v
1kPWCVAho/arnUZXby6+9JDIKNP0YJFhxtIvN0668upZA4p/83SEaGWNys2GrOC1
y7D9U6bliqCHT2pUtuGi7coArx4kO8z5KzQ/7kYfalgDOlqeEqhOju4zcMrL4yOl
QtS/zkK3uJwOu5sy/dpnXzyH9FZIxE3oKBb29lkIaa/YMabNat8pTXdSdiIAoQLN
nuTzn3TYOCcOOV3ekLg99UMoev2JOj00Qjjnwb7NfExaxRbuRmiw30r0gGRJgDWm
1xhuq6aEdFz5AvYDc4nll5RjI57t4VkbpP5AR1fLRuoN89W7T0wwsTn2kMFzAvF6
bM+0DKzV7lFm8StI959VITHuww1SGZ2wPD6fRYlsfK6KDh87Kr1X5/A9e6laHFt1
ZMXIILjOhZ0a2EaE6HFk77WYhoNrQiYaZmciwwFYN1NX2lEeJHq/6tR+BFvWRi46
lEy3IFs3kI2m1u8C4IVmXAIMFfqWTxRse8GHMjKO/UBqC45pSwppoS1/3hoV9fIv
zCZSYNTDoByK4Dae/jop3xqkDQdjAMirD8YVpWKf6BYbzIkG/XkpeGjPVxWOZERS
IzxnkAiHXF4Z9WjfQYwQS9uSe275ObRDMgJIvw9BYwaLymURMDYuy8ON8Vs7+sn0
mxI4nJcHsYmBdA5LphHZitSxfK0AeP2B5waUEP8ZCBt+1xVJXiCH97AuHai7lRbH
GQgqdCfMhqAXyV18Dz4R3HukmS2tSkH0fsxBnvSbOwYRTFN4+rmwbMURL9P4c5vu
IAG9BR9Y9EBytGpkRcJbq1j1CjZpT25g1PQpevjUn1eb6NdkCEu2Hafa5lMOzpYF
76szBiZuMUIJqo+aLIuh1unc9h724CimHYniduJb+nBG5LjJA9DrIj8IGCS76927
Q0c0WdOhaTcHhEIaH/GAL3OQBFVRfzAqzUslK3CkM796xwUG03oMhwgOAJI5bT42
RMIfoBb/cc1frOT3Y2EuABteLilpN6gIEksGskHoDQNVuyaM8eo2OQSgBU+5pG0b
CDlOo3etD92t/dCy5+HEN+igGNw8Teesy+nBytkCKfdtHY/XEFBJ+pgJu6Hd9SB6
IVFF2KwFN073i0enTMggUrcWS0hAb11Q+B1rQZX7WV1L2c/4BeFBiT2gF5Oyod06
FfovaruKllBT5yKVUSkOkmu5v8RO/sLRsaWwVQYAjyyPIfEKBl7gY9xVGZ2I+xxQ
DD6qVX1z4xkxNcbIvkgKzA6tbEOF0lH6E26VutkEDrpsw9nlziRnwwFG0QOKj5Z1
BDKnDWnU9MeaCtmxxpWWH5oVbg9Gt8cDHAbAIvnUJULG0kCtqP6z3aVJAzXc2FkM
42vw+YukuRJU351ro1VHMcDQ0FB8yMoCG7CY+VjhF9wVPBbrAbMX9ChMN4ymcTXO
FmlC3FbYmi+0bbwKa7MB5iV+BAYh90pG7fRXWf2wbLtdSDnE1z5WwowleLm0jPzE
HCxo2BFJGZ/zLwvScVgl7u8Tw/MG08GnoVR0GaQia/uyQOndLaNcQlphGEGnsTiS
q+XBTVrwEb7/sBIE9nYTVf2IrAkHH7R4NrnNFWlUBvXGxvUtpyspHk8V/UAnypZi
au2vSEMaIABDG0HBsOAKBmV5DPrProL1HEwZ5AYqkxuh9acmkFGQOGPuJQet1CGE
JEPNvJhw/ha11QOhV1NjC7foN1kuMXHkbjtUc9veQyJoyLeW151Ax91QoczW0+3h
X1c7cHQiCI7zu1sKrErK1KeFFdpx+dlDa9uVpLTrL4Ecl+nPBFVMzYdPy0YsVi81
UNWIgV6ody0ClCH5s9bMFnO17W7mf0Fmd+ESMC1cWeK8zIuupi2KCZK5QYbfCxvb
9s305dLhhpbiXAzcnwvq58TlLUoXvDRWlcQ4rg2mxwpGCSbjIqViojV1nt91tiyx
Rg0HNCG9OeT2iDPDoSIgP2WvSUe31iYOyzU9F11qTpE5Zwwvh7hCayo1ynyCuYu+
mlZSpI3nnMHLcY5sx4t2J+KodpsIS/Ry0KQt1c3+a+1B0N+r4uiAZ+86jF+MwyoJ
8boXzzrN8wkIB25uC5f8tJX6nEFkgYVMgwAW/H8r001I984oeNIMglqEr1Z+TP4+
H7/cLN2t3FV1lhvxzRp74ZwKqMFFWEkOdHOOAamZTFubFmR74qDkErQWQPkn5mkb
yVMkdJw6jrlLMTlxSqoBQUHG0V30GGmY9QI9T9YC+aPqEeSwckG7iRkB+DLW0Kfk
69XZwMIbPpz7XGbfxkKIIHWy8CQtWxRvnepR2iT1DsD4Xj80lezh2Lm7hO9mVDvk
8yMJgULPJDJJScIRCXxqs7gs6dTFR3i6ch/M7mK0F32hGRGOr56IawguO0zjfsvo
vQQgMeHs+882V0+X80YwhzzEBLn8R97Q41gsR9vVGYQCKPpVwGKyDNFgeEtXIBm/
kf7l3B195pvALEQ1KZHlO/dYk2GoI2xUA3iw6HNMc4/olz92M+4eKM5sy373jFoY
KqZTnMXClM58BHJbqOxFsBEZoEqb9/EFj8jJVVyWBECqg/t7SfrCNlxzngOq0a9g
Cl9Yb6XQHmEBDthX9rb7MW2KhUt9+fh2WhPvD9R18B5rUw5jSKyJChZsqOdtNSTt
e8OIdmHBSeBrJUXKD5QZIXcv8IR1B2U17hQn3hN63REw4/VniTTluLZAMgtcfvLD
Lz2zzAObKwvZcLNZel+KmxihOKldvENNX077F+FY3zhDRFE88EMDopfBqemcPjnE
J6M3VB6lETYnZaWu5zsnIknTfx3uAJNQ48MEuTJshhsE6brg5ddJwbokga88/MFn
PRVEqW9M0xDykpFou96tr8HeCALpi6PcMHFeVE4aeYHjCSB6BfvVUS/jBTGsndYr
sBFzJ7s7KQEUdE6Vy9px8XZrvF8w7WY1B+wSf2ohbdinzx+ueIISdtwvsmKQPqWO
OsxCin9GC8hHES0YfhbZbL44gWFuNkLl1sHqGY5i60miZA4xNDp3l+L7mNcwoJzr
bp1w6MS52MnB7Ss/nBhfLWu8VyjZKeM+83MtktC0OlUcTPuiRSvxsqzOJvNg7CSS
iNU+HaLdCjFwauXbuhvbQayQBJCyd9CWhDuGy+VoF4r0H5k3uOtRDt9VlTODn2to
MRgzgw8wfbNYWD0Lb+8ZWXP7zWSrfQUGZZrHzjsW0ZGtou5bbKDQ+fHa+WgV8o8W
yWBqiS2MPndBLkzv0Ru11okrkPCUQHTyaWcY+W0PyJ7EBuBSrw7/cEDAOeoVQhT8
w9B2L4iZLordGfNsws+BMS57rpy06T0LP7iNEVoXbuauJFtYlwm2P+hOBBbWusWA
SsfSgL9+nUBvothJI3FEHxUVtF0ekneX2OImpCbKkR0mopi9ieFtajuhpHzc9M9M
yvK9Vvbx39pybnLifAzMcRDSdr0bpMmtbOpQVqohMoTN5yYI2APW8pcDluaEDyRE
eJTkdK2kgKI1B71uDGOolk2oCDPeGjm6Tw6PTIfQYwU+8V3xJ2WMsVgrMtqHRHb7
jEJGut08gfWH9eDcOTqtlrcudYMSh6ixvSvocUYtxgZhw8zpB9gVackqqWzafc8C
Es5/5D76A7EFsFzkPz6UuiI+h8MvuaqQIY9ggcrRbIuAEdyCcNUYIhFggu/2UwNB
cceY0MluvWOE6EslPzcPAGzgC2lsVBlznQz73FRg2D349NDLae/WLb29DhLMFrxu
90xEAlQbfUhESjU4MjvslJe+Crzwjl9UcTzAcIhlA0NJ6NjXGsE/SvxKqakvb6lw
2V1audyiWqHyLRAvjWXoS1KmByk+6QXinHKRB29/vtyVNxaNMn6D+isA1H5ik2qb
vvKG+lDJ1CStHsooY0dYmp+6Qnl8t09rXOyomznyi5NNPs49JSKlseKqfI4reHPq
4tLA0hNBzXfSym4vWEHuJOu3hTlDXBXtdHnolbJkDTFuzHwFh9OaDe5i8ZQHcFgB
Zz9wrX7qVUiZQnUsXErRL/1E5x0clanCYlCHSMahmoefZrLltYDM0k2uQt/2m/aF
9gYcPwT4BfQkWIZq6OBlT7pOtSIZV4u2A9mJGGzJviBeDOl+m3mXC6atsvhYNDqS
OA3aECcOokvOfP+2UsczHyndvWh1c9ReLzESPbxphMKEJ07RBqc3BmSsQGORiM7a
aBREzzDJnuZdIqOr7e/ZOvmYufzbYGWF0XjqQCw8XE3OTHhAt0i9m8sAkz4SCxre
xxjC7/3rvDknGOn7G3YzcOc1oHsDmogIhc156dwwkXnAicdG08DKP0ef2Mv7Furs
V4GZ4hZfntvtmLwCY/Qfa2BmcuhvyldBvssoDPsWKysCFkiOmxj/wvPfPOT8Kkbi
p8r39Y5gUbl6YmJuiHe1vKvOje0ytGJ/Nbfmrux4kGnLOSpiO4gXvTQygvlTLLRB
U0pZMUzu7m6fLMPncF7Pvh/dMl2Qe9Ktm776UrZivIw5Y69VAId/NC4VEgU9DYuK
6NI5uuVD2v6F+PNHGILnKo/9yJcG7TGdojuyzEQObdSc6KKNFrkcBIE33pYMohvI
LWgzX9i8iWqJiGnnRW5lE89rDS6cV+lA8PekZz6+H2LlfAhTmXwfMDJaeS+AnhND
jSlaOfNQ4o250pWQBGbxKWiUGYBC5HGl4Ml7e7wPDdWQhHo8LJ1JknTfohv0Sf+3
ydThvEejPgTh4AWblWc2ieuCOsioVz4MPcsXQFcD77VKv4dWrTJYsxH9O1IzNtZn
Tl14jpLJjfBVieFabMnUm10L420I31tOg7sR9G/gb5u/adoIHnu/LsxLGd2a0roO
FSHLwdTgN6rw9mPvb4R7cboCBfhVHuXK1toUdBHnHZcOdbNO4QEv8KC3Gvspe3ie
F4Ex/JZOHFzmkZ1xjIs12tdoiMcDHy99mTmS9zHxw+L2KyKgkCRpTdqvpl4C6z0I
b0qH+eoBsJNfUpQltv+MypAK1E4cJgp8u9+dT8VIVrxM6T7I/riFFJ3DvGiNTpg2
KXFLT2psMdOyUjTcEX8GrseIIIp4UMswEM1ih7uqlaN77XQL1FfbHRxsQvPnyuKF
4sXwIBl8XH9BXK1sdOcgrmxrS7ARasGK6+DxMm8HKqfDUcRMYG+U1hCHkYyRDlY8
F6lgZ7FgyIwBQPq7Lkf6D3tDvK7q0kJN6PV7NdUSYYSdFlhMHRH2EJOD2jscnmI2
iFeTENxWC4Yc2xpU7VuTqpf49OBexdaIL/VwyED3II7Fpf7Y9pwIsSBVktqJge/g
bAHKjebbZFqtDHPSEot5MXd94hdaVrDXWyJsKM5n/8Vy+RlKyLOpk6Rlve/gTfNV
p3mvk9xjOd18YTzTZTZiCpmSwXXwSmlh95I9Dwb5MO0e+xMPpJsHyVFbYZzWJwu9
kim4Tdja/4T6iffzOIhZk5RCFkp8j/6uz1IjYqB8c2Yy/zZYuD7+iG5wh/OZ0wSt
U376AejNSDRvBZnJIR6Q+mKyJi68VyVXFZNNAJrTMfA9PBaOah63uHm+kdPRdsHx
YIxeGRudvxFwngfjn/U1mXLEMzVihljXoakQqx8TsSFr1fmYt3Br4zpivajFQdiR
PFMoZ3o332LZG1e8YDvQrLCK4pwu+SA1JnFP/4YUkSyGWpNZCOzqyvvNda2YPde4
M9VmS6xi9Q3I5IAqV8PHL0eiueWQAA9rbqakYCLXK8F6NXECymYJpxCWzmu56GSD
f/kLBbL1ZtaYfZtl7LbwmfNVqJxCEaPwt2ATq5VjAjLxxYhkqod/rcAB56124BUe
rUgiFusumrh5Fb39WeUfByYeFoZLORHpPW04PEYD0GLHdPBN4x4kxF+Gyp0ZsuZl
VZAbed1NffATs1aD7jcujSWbp6p1390DH09g58xBOorTK4sfWNEatXdkhx2QmPUF
3/gt//GirwyPkd/+dGI3UcsRp8vdNE4J0+oTlhLDLTVunNspWaMkuOXH3kTq+agK
TeYxEm9cG3O59+lDU+MRIU5eCiLUYqmx21/RtrVn9alw9tgPjr06prNHj/8+qQCY
yVyDGA3mEP8WaygIsvYRHegyrv5Y51lZGA0drehPdmiWJr48NZbsgBkyLXvB7h6K
m+eevz2gbTe99bSEv7qaxKcSr6GmFASJ2HSz1ATTMshocZgFUVlr+ugWDqFB4yj4
CJV8Hg/tUnq7NE5wmoyKomQESIyKmkqYvPPsFwZWNGcAJ5U9FzGeIOlt3L/oYO2/
pqkJm6KfP0wK9DNqxMhZpJDOFDhfxa+7ZXdYEu2+z67BM35aAYSbbl1p0OmKOVd6
HIZCkakJ2AkSqA1eKPRzy0GjHe34Gw440LvT5iQmyA5zggOzn8vI4a186X5Pt/M6
W6OKzwNOxn3d7HA126FjYfbAwpcaejn8uXXHSHQdAHrwoZD6eH0tTLCkZl0sd+45
OLT73N2jafVPdnkDYGpeq0ldZcxcZIU7wv7YKSTFnQvtoaKm0jbVYx5Bjh8UG3Ps
XGt7LmKZhNy6wFi1rKDtOfEXNQH9yLpxZ/GdhhGPBdbn0qF5yTZ7by4XcCIBF0pT
Vzn2cRf7C40tFtjQnwr/j2M1MJHExeOFCUzHH2HZSzYySu3D8kRXcXv+3uJC8iyp
0VHq7E/hUCsjcePFv3tsnWtAfDvczFM9GEZjfA0wOLf54Q5nplSVdsFP96+G9BYx
c9uEQpWfg/Am16cYFcoh1yqsKLmd1bMV0ZM/aND8tUvKr00YvbiHmMx88zEqmPSA
V1cqTxlkH7Ql1m1RL5CPkZpF160fcmaJ0jYKjSKW80WIylTu3Dyz/nKpSUZoLkJc
1Tew7aDwCfkf30KOv6B4LgIZP1qllc/a3sNEqncXOOoJHaitA/O/RidqTkLPeSXu
6QOunY/9k5lV8lynmBa87Tt9qOcOmI6Qp+8lps8xJIJ9YOUAmVhFymtIj3Bdph66
Oa/eqMWpxOUihX26TuB/Nk8mg0exCo/BCqOvdL0G3BJTERS81++1dXVCzwIyS7gj
tQqilyHNs98tGzoU0rMrlrtd2u/XljJw52/YA5Dg6vM40qw0J1N3d6RSqSvaLJZY
vLzSt7emwc4QLiyrC1WEmjwqklIsVIqcKgR9W9H39DgQut0h4XVhnPhiNB7S4SUb
RHmY/FOp4E7C9C5XXaKLBRZJ2xFy7B5GNURonFSSLvkXM6AmZxy6jNuLhA0X/dOr
9ektw3hXeSb8VsWdwBHwAIh2+pVL9t6tAmUVTIrT7jh0HXOMwPV6y7idGmRLQWgF
8tsSm6HENA1wTcU3bLuG2PEsZuc1mg8Dz6h2cEhO1cQfBa+AV8Rt0urvZDP/uYKk
jBE7hssXf0Ey/8tDePed60DQhsZ88DE9X8kTG3SiXs55qgzXfI+ryB4Mj35E3K9a
vY2JIWsSHM7c2V6cWdyPAymGkcCPgw/X6uZPTjDpyF/xr8ryVZGHmVg1U4EWiGUI
GuVJOJ7fBxJNIiPOsWqcg948gxhNI+8MhvWLw/vj9DIfJI5DkojHzrQ/NJKm2Hp1
x9wMxVjonqUJlcrJqL9vQFEqZmEyDQebpTSw1U3HeHzggI3UGFR5mE3L5XcZ7HQT
B1Q9YE/7EEqqKR3RQSwIVOl+6iNalOSq62GyIcSt3ttDSNJHycOloR3M5FKBb5pM
pV1NGvCj3h+ngn5QWGgSd1aM4J5EDMJZqfSzZdSOOmwaQciZDXLlUQ4XPOpcvqLc
feCr1GN537FnzSMHgrpTaarUPfzMnqvGXEM14oxl47CICml4SVkZHexT4FZv8q0G
+jjjX+o5ioulaWYwZu4FC0A1BduXhJMTrtOTOChpsmBmYTA+21JkMHTOWwhDNVJt
mldod7NBUXux75nzh6OnMpj1PftSjAMy0zSz4wZ8jmQhsUGH1XDvqJI27KX23ouA
jzsrSdeypXiDkry4ktgh0t31m4RJEwK2i0SAsT3atXe2+I83053dm+mVPokt5kFS
slMY5sx1Q/GNYPWYEbDmmDkmc3mqgvvBK2dozgPctdTRPU4RZ/Fqo7xceKM2qoTo
eHDXduKlnV5KM0wKFshwPigalzq5QU1aeY3cFzWbuhQnZTvyHl199rOdK3sb3Gsz
McdHBwz8iKNwlPsayEE9fpRipgREkvWLib8sgODiMI+vsy+1mkJ/RPGP/EQu7psB
6b3VZOHXXgc8V7DcMM4Q2o8JqQArRBtBt6Qq0jjijZlg5XFzN+/GBQkN0m582zvp
iRpBWnCf8yMzGnu0TXwLJaFg27CqlU0FCcf9sbBVQGR3i8UOK9/+ki6GZIo9bFvV
iQnVHGdJ3ddNhJjNS7hWEjpGrUBG6CL/bBc+RQkQj3frmAGDpZe59UXYvLRwPATW
iXUdAi5r1s4eeVvBMOEJ3erAP20lWpr1xep7lZRwLj1J3xbmwaOq8MCulifMk6Tx
EY97L4ewpXEF7NYBuHxahe+Q7kalxXgUAq4bX5RhAH9nsEKaGp81lmXTyJWkjJRx
j0zK7yVFfZVfOpjn0xCjHIqmQC7icG69I9itaqJZtv9o42TkcfpUUWABCvH52kLd
uijHNK448sUXbpyNb39uWNj4NC1nnUf5DdDfWNiOGvcm4Z8uaZjayn/8BvROwLfN
mBS8vmKwN29a0CMVvgjJ1DZ9hyeEtEOUQEk+BkcGro+McJ1UnLCYt1NQViDYCEl+
+JksSatAet5myFWY7LheuhRd7W85FKrKDLykZ+xFvogeseXFqn6i75fIrAy3iaMX
n6eJphlX+fW0YbRS56PT8hPzuYNSXnubOIo4SyfqiKxLS4qWEveMLBaLX//loS3n
9UgzbuPtxSrGIXTr/1yFSm1sV3FGhL0eNTy08pst/hxs9s0VhHqxLCEV0+nxm9v5
YkrHqS5H3JGcuOIurzX3895mPx1zKLmaNVfl+vF487i7xom2g00zXxLUJt7dXwIb
qfHORSN/QwC0f/gy8AYsZmr1kmnKQZvS5TsGeXfmeHeQgPbYw/460D7tVeGMD1Fw
M57dKJMAjKtjQVs90tGDc3bgHaG05h5hSHvrl+tM8HmpK3dXc/LNZA/L5ztM9loo
h1tf5IrJaJv6NedT+HA81+sS8q9RzYDl6XupS2amxrAfz/XDFYIS8mXxmuJdJhX5
IfMMtCR0HqxLslBUQWSQlGAAhHjAZzIZYApQ636xefwyz0xMGgJmfZi99Uaf7Gk5
H/aHG1TrRXVc6J/jPbnVZZMQK/RxQaZigPTuhpvll/S1tL1eWyxcB/huqutb2BlY
oxVrGH1A9B6T0y5UZw443OA2DO9kx/Q79a0dH1fPkKpCmxPgh4e+D0+utb/x5JQU
dC4m5bHejzPr2PcaXn9kbAtScxGYBZrfZuTH09NmoAS9qG37zC/7/SLxJEeIIRqM
9SHUmpasKUDuVtwulO/hZeZwx0cZeJSQMDD9uE3e+ibejNd5bL8aMAvXnVKX7IrY
rirtYUVJTojp1ZfSJ1bd/Q6uk5mK2HSGZMaPFIzbPXJjWltPULaJnJL8gX78yTaV
uMfAkb4KlZAPxuyIsZn+Q8ApAUttQCRtm6rg1TjrDV7vR8EoR63+5P1O4V6RnUkZ
CoEiksySBBvqb2VClYSgsWCLs79WqnqQN5UucrDKP5zbiPlVTjmmKrmD37c1ubBU
0DqUfcNR+Z2/pYJwGbQQHasz8mf02sDEGu8vWrqLrVuxUFWimp2ZsFikA+/IStHM
b5v2Zx1XFYQBtb5IC4A98xhM2tbVDCbHMBLpVl3HTs9UtmXQA1l1lu8Bd5sY5xyo
N3lyrlLjuFWSH5DtMP6CuIYhfpDGe0t/NsMcSNEiC7wS4RoqYgQcWLBqY9LV6K5N
X5sMzEfl59Wn0xOVLUkEeRuUvOm2wHiHfftTdKOVsNv8Hot9hh9J6Vgn8DsLLgKL
fkqIjW36YT2CmO2sIyYKE+RryudDLOMKOaTZN4MTj1VzsONj4zmIqZzndYKw3Qsa
h4JkuxccedYK9iG1Yem+k59JqpK77Edf4RcD9osKjFEEOAea7tTiQw61vp2Ylg9F
a8EGk8TIlatohNpzMsN5Du1CsacGtUWhzWS5nftL1IJ3fziZopitZvAm5xTtzLAn
5x2U2LUOnmaP0yPgS/2XYOrC3VRHw3hUZLZJaFagdbCT3++UQkjLGV6Z7aw4QMHY
r/U1Nexh1PpqVemtnIX34nKJdpRut/cqbRNqZmTQnv4dYI2Jy+2ZsE/OYD5HGc2m
inBBZA1155yeZmRVP24kCXoKU/ft1lJ7OGb0PrJ00wa7aCfDuGIyDu4jpxaFT4Ae
qMRCygSLMkYyjv+DBT5EYNSW8jB4ccpc0yXgjgIEbjpbwTpF948shkmDzGy8ROr9
u4J+JiAmUOz8r8oD/2iW+O6HEzfzONTompecFvRpi/rrLRs3T6n91A0zp5zGvAOK
5GYkugnp8r46TTWhh3p/UHQk3FYyspnlJwD5d1hfIh8R2r7b2ZIll2jAILeBR9tl
zDvbeLDK/wXoj/HQcJG4+bXIXYkGHFEVoqYVnJROF2tZQWkFbrxFLp22srLXZorn
mmb0tndT3CciDmT+tOLaUQTB+0AEh6NWf0g5uAu16Xu0gaOCHSL8IWPfSYJ4I12p
KzSVqxM8v5DBw2XiW6lkkrLNiI31QXR9xaF1lAaxzG+22BkGD6LmeusU96OcwPoN
97EIYD0JIPYV2J4awD/y3BLaJ/yf49EuxnGifHGeu2Qm0Jti5T3YY6TsrYuuAc5g
gDTxfh2LwJTHAAhf5PGFwEzS3U0bxgRU+uZ5WsG6fkSjUYvcEOl+J0xPz+AldXSb
yaSXFv93O0MwpuZu3spNRiQuPnjELsYMiH+tz6KH0Otj1FEOosLmFWSeyP63eBk7
2k6y/4fg6sMdb1tb7sKAZbCVQ/MlVg8ylhXSS6SBBXDvnLooZ/0uZTrmYk0diWji
o411bJmU0UyVB/8ZcDYSpXJCiJ8ydXjxgE5OxlelvQWtMjSUVrFltlR4xk76UQcA
qtw6TVusDBpP9+9eWMXduYe5pb6qP0vooiKXvEq0xvcfbvFl4mLnp5HhqsFAPZpo
H/e7p9TmbX4ic8Co3/cPUnOtPmdEudoAnqbS51etz8puR/M7DzPZazWU0eV1Xj1R
wloB7Ufk4b3mr4Av0CKuK77ugdzvOgpSYY9xqxHx3gu+T/ID8kqsCuBbg2ND2arj
k9/beuE9gdpYqp3MnAGlwQpR3s9acEukyLd3bjnvMj1YtVPaGYD47gTxXLZiZDuL
iCumdPbU1gJuMRWHm1m6f4WC/PxwXYUF5iZgY3JbCM1sVFKsBZnaoUDZ8TKazC+P
1REoJ5p1IoWWP4MuQrJkT53NBUDjhL/Vh0Hs66Ub/16z/XDmwQ4RD9clhJTGR33M
D0oWNAcJlA67fTTvI+JoUB1CVJtBO4fkFjNDHBC1Ak62M9oCcNIGm6pfirN19jlw
iTOGQb/4IitcTXbGA9NCGwMzEjF5jEpzXWh1q3iCQWNvKNtoOoiJZ03rYDVtEXPB
g/qz0Vp0n+F3aWPT74vxmRE+K2fLGT7I/RjffL8Vj8o9RLD59dsu76qiAB0egFd4
HIPJWBiSS5ZvOmF2DHFFx6pUgf3VrLs1rENqO20Otm4Bdv5ZMOSh5vnsfO8PhIJP
066se6cedhUSjDDW1Hm3PWaLIq0piYcssgLDCxb0PUKcX2dFc2fUMG0P7bFL7P0g
zZqjfMw4DIXMiru/YwaKkk35X1LX7y29P03rL/Sfixwst2u/eKratijYV+3wloiC
STx5Ti3Q9YtTmmFtQog+3ROAx57p+57ZKTozpnBFYVAnfmbiMzJJv0J8gZ05zaky
BKhhv5WcR5ol/zegWVcf9aypuzd56BCKYE+IKUxOYHlRXLRIv4oFl13kMJj0gYxs
GVr/JNjG7taPV2p/i3otVLlXZ0vq5RfKwWINneELQKGLItfmy93la4/XjZ5LMGyN
YsjMAsnTKyJzeKjOST3rcacf/myw++XNJcD3ADeHsbs0pAOUMjO4/xi0KaccPJ3j
9YmKldXLPi7JTaKTrkIEcUr/0yePlRBzNEg+58dc4heEu6zkLxs6mO9wYX6XGXXG
eIFLKE3DBgD1rIzOCXImllatxOsZJbztowPlZj3+JUWr8gmlAcP4cAaRh6q6aENk
iq7Xi2yu31ZlOyYsVfgX6brMaIj2Lz+DPokkTBC+dQIghDNbv2K+ujuEZUncS9hV
xFIA4q+P+y+piKknw3TQYDXNtXEAe16UVa3qc+lM7NmCtzqzTHfVJh4zk0S+gtSr
uJk1bxFZdY07ZXlsivri7f5aopv8oCT+zUPNEwEFT6N3LIA222EksLjlclWGo0U9
iwN7n19ONIEL80OkYpMy/aRYlRXM81p7N6LlTgLfKVVMtXrd48o23HWAAzeFPR2u
jmJcgREXxxCykd31dxA7I8Geocr63cE5dKWnujW9DsiVGNmBihD+ugK3+KzIOrbB
zAfwqPAhrsyNNVoOX2qod7BAWOwBwEeIZ4RqTQ9xySds2bEHw6E5XrRbaqfoXacC
TsHTrdeIEYOIRwbAypwZ6jvb7Cyc0WBVgdQtXltfxRGjrFipgiRVzOagnV6hoez3
iokIpBKYTBEGyzDIoLOQr4aekdYNJ5IegIA9ehXZSrEcoh4Dhqmvi3VP0p6PEdDl
GBovXoSgTPz5NzXjCjSZ+cTJkCAOZS6n/Apc1KY3llsB07m50MenBJYQb8lpbUQI
5beoKRL9NN7Xcb3Eq7woLFmnxQRGp4tRmLywX6BWTWzw30l0HqYIxhegNrAMfkX5
xAN04Vd/BwPOhehrbkTN5RzBeLurObQLAIXbW7WASmO1TzQZ0Jj8p3ksRcKtUi7J
tPpwUnDSsRTOcycMEK57ITBqFXk4c2xpsDJYs/XUhjfhJVFmjEjRxwtGnlVAYflr
EIqKisjgHUxFqApoZX1H0GuAvHLtXFgmK9b1KTUMoJbCLrl7ftxxWUVxTvnH9wSR
Hfvk6QqTIUWdj8evaFoScajkAZB4wOcKB2m3WoDvbpUvqywifmlS+im6vLG0NSaY
ij1Rh0C/G6Y01RQZ+IHIIOGBdA0TfOJolRjKIeUgEVgygqHwvD3u3JxVZDC43khr
UXcgFm7PjVM9BAEOFiNd2amrL3udw2L0yqkGpaqP0YtIGBwec6awCyjJhWhGuH5N
YoGgs64SxJHSUOP2bgnWotkqurpbn8TmLovu4uQUo29U+KcKp1n5BKC4j1E3uyw+
2TpltehZfAAUeU1aXW61M9v1AvPUbqTnYoMeSEKW0zLsQlZjvNpAkW41A/L7erlm
SawgCZTG1WiOVVnHMpa/sm9gPPKVOkluJWK03cYgz9OiftlHGqytvTFPTVcp8qGm
51jWOZnje4X85EyLQUMUz76Ji1bUyf9v+RsMq+CkiNtxwhpe1hoaI4JATum0sEun
Av2LpQqZNr/5TXKLOo6XkGnPLQcuV/O5B+nU33a0xJByMe3idiZTIXx0Nr6GCP9m
mCvkYLpfS49dEI/Jp+Dh4FCRl+d6THfgjPOaBaJJnhld1uWyqN3dMc73KXrWagwV
aFkJXp2YnkfnLgG0R4BEAXOCvR9GUHxi2Mce9gnCfpQ9deS2SknOPA4uzn6ZCCIQ
GmygqfEHe4QpBJCN+eqnn9e7f9bLGHpK2nMa4T2z+GMzDl3H7jfMScqXjXVaBKL7
mSnWFSucTF3Uqk2olkLhAImGS9Z2PsHvKADcbpL68AiZBvNsbSnQq+2CszMCYO6w
rDPiyJjLvR7R6OChCQiXyA44ppcuMmpnKktLk1adpRXqeYY+uB+RAX3AMK6PFQgX
5mG3bFXATY0q9qYEzovyruBZateCZTL8WTRl+cIVYbpjGTt/yc+odro7huSoRA8O
jBfo+mRR8fF5iZWTmUW6uI5zeBWws5cuwvw3Y9Ajw9DQaWaRpmfsKWupGg7AkDt4
JeaseVXNDtKWVLivtLnkG31jxu+uq7x+1Uln+89qa/CuVTm5nptr93tQjpG3K4G9
5BUJR4xPePDND4KKqNsRELDxTngpPDVDbHndvAgUZmRXUVKNx3oW5T3B4pq9kQ8W
8t79+qNQ8mrgxvuDImHGQabTiHnV0nmBZDMfY7vDhzYHyC1q5J3vHfiSuveTtHio
ASDZ11KHddiLGqyhXq87a8FqkL1fQP74YM/ajUg+dHnl7gJ1DuZpkDzIMjy3tEjX
WyQvRGF3HtbL4xlhhgwXhGOIhrIUUVlk5yVDqelk7PBfoldM1p+SOxl8gQUM2u8V
NHNEHQ00g0QPljRJ0y8M3wUnmc+rsM9rAhIjONFAty8kEt64XIe0+SprPWS/S6Wg
YdNvgRUcISKynmpMMig/MoWzCyhb98tgnrNHKs9how7Am+/tejgrpJ/RYeDgTL7R
eduR4KB+oNZi/VIN4uB8CUR5wMjeBNw/AHdfPoxeMAM4Qn2nT+Bh06jB58lupooX
kgs16JX2iTrvzoZbTbs0oOT78XlLIpoXl3PPeckNTsjyNFtQ+5M0BIMVKvD97kGI
fpac99MxV1deQHNfs7irOYpBi8cTQhT+pqt7pakAor4qpSCrmi5O80oB0cjMEJRC
BYUgKZkbDONgX1/7c2Gxkq/lgD/OsWGYXcCF5+GpS8VNHlrc79WgE5VY3mLxcqkT
hRa5TaQsc1qwjKv7F7JppUtGJhcNVCba2VKLqhakmta8UY0+/B9DygpaWqQdIFyq
dP3KUKEbWc3cW6eYez25VHpqpFIYUFb+JbH3cUhrNNzoxxL4djA9n8asVa1LkJAG
grcivUgxSjiYMjMju0Ycx1Vz9BUwevf6XumFyVqQ3XWjWNmU5k+Pw8tw21x4Z2Cd
2mvImqbi2hc1dTjMx3jOr3ljylAjF5M09/dgtFkho3cyriWbcQ3k0ofKwSve7vdt
dHQL0n6f3YFlaYnlUu5xvK1utGYIOf4BZsnKiIYkft77BV2EBED7G19g2Ytfrd33
chrn8N/JqnioQcHDLPVWlendew7TLdUm2bY47E4vOMrcOCDZgcxTvWO9FbMhu/Mi
ENWf+VcEouprYs/u4ycoa82EhpUjlaKPiRe9gTEotnStPzBMEexTVT1jDUfbnzf5
IoHiwbhqBtZXI86PiyO2qm7oKecgVL03u+9LMGUW/J+NEAShbYKOVi6vYmWJa3ji
dqBoIbzpwq1G9bwz211wPlqt8hQcpJZx2P43pNRC9gVuCzHy3BlQCF4NxjkJzQF0
4+H+HNXdi0zNn52lmBZS7WcANKP2x0l3Zd/9WDZv/+IuU1C4DuExG38QH202GbAv
4zaFs+rxpafFxrQfWMmhL7lF6QXn6M5Vor9UdSQ+GR03b6wBZaN1ILv/hahZvhJh
FsQ+1lborW+A4/dcT0zfFiNIF0vO4x1o3h8EFYqtHA4sY3+3luh/4KtMV9VWHzun
gp8vRuSFHzvSjIIeA8iHLcKPfuKvzS6UHQX1E5BAEW3v3yYjgRR6EwIw4tk9HXPE
JCMhsk2y+l+LxSx9ekDQ2WIFH6kWU5xeUlqdJFNX2oqMZiuq7EPmlS7SFOQn7sfN
FO1sO/V4bZ/CIaFTpYkiQ4vjA51FqnXendqaDhJN/G0N+PL+P48gXtqULXwgWFiL
rULGnQELL6lkEHbozcIZ3KbTzxTMMH+vo5sdLcuoqeuwkal3MpAzLnwS8RqFrTkC
grTtyCjkVq351lKG1aJcSSpcGSuCzhrVPImkjnmQ4s92NVnk0bGb+do9uImeiy93
SRTU6IkVOIa3XXB8xVU46MNuTeccRua2MB3S+6uzapx415kCSGFrtdvzOwr7/bw/
Jxqo0my10ZV+fF8AM3MEvX4qtyYuBMeBseKPJ/N+4LZiRbmCThXum3uCRJPs1UGg
efcEy8SJ+AAQ88cuu3oeA3Mml6uvyKx4iUdTtld2Lq/3dNtzmV52+cy0KW6qsfQN
2DHYVVmc2WS2uPVSCrLNGqDpc8NK9eiY24i2N+XAJn7MyGXSgAr7JSVm8fbWEw56
uIl4RuVxpJQOYHsyGT32KXayn5lt5JD4g0n6CNrx5uL7s5X4elSsoRuzwUfiBB+0
ouH6kqftwJGZ5pBo+Y5Ryw8Ht6bxu8WSj3sWRGkQHRbHAU/evdKi5e8XoqnsJLDP
QOsjr2ujnZnIO3FoefpdIzeARipPhrHEhoR1A3k/LPfPpm4xOkePAgMoSTiCCF+a
Y/bHl/W71Yjf7ogMezTQ6gpRmL6eoXTNv6msFdOFKPD/8oRtz6KjQlt25vFOLYzY
tuKYhj7kp4rHOTHn1+5ZZF/GE+rZPyuUa0Js1PuJb7YdBHKSOmh7jhuVh6GXqJ0Q
PHXq+DU2iIOyMUm+skZ31PUuIafkDDewTwWOPNzRAEM1NyH/OyWShM+1UfRGvZLP
5uLEh9ktlqA/tHSFhABKMYrKT56HCWDuLfPyN2BBI/FPTNwAl1QHNCsKRqOt9INl
z1WGEB2Ipt38RNA2+MG7zH6K+L2r1MER0iYq7y7grwRiPK8MF/AJNPojUeY+HR7Z
eG4EUg65XjEWEClzlby463b2rEEuzgWHVyrowEF6sZdKTvdA/ifANTdLbLEHoSbO
7cO/rwr48yxr2UHrKiQrV5mTA3KXR+LqSxReTVBHNtkAWPMSWLniVP22bnD5swjm
U+z+May+YJdMviMSItv3Ci5cSvSKuIqMPO9NyF9HAki3xO00o1w6OTy+BKKZrl53
nbUVYgDo7iF6kJQrPIpvzbYoyKylI0KfitUBeHuxmBNQBrT3XRfi7w0oabzK5ftn
O6po+HBXP8lbPWMXIfZtKaXwqMUZ75nJNMJ1Pd421O3+jxFcOkpXIEUlG2kDnzas
faB5MOnUJBIPDzhsN2m+qpm7q15ImMRuwBCUc2m2KgopryPyyxGLjjQ+Pyzrky0R
tC+65cikxijLKSQt3iXLH9cYxkDYeg1kPGBIl+vKANolCNU0WNGCtSjDEh8niFr+
BBuWmFNsV7sDrNpA4zl1qjyTNrnUo5CykmJmDWSHtGn+PaUpw3sDu/4suoU0XlKk
oR9KkMzOWtf9Zqj9G07ChgHW1SdrZQHqnTYVNFAtxYioLr03ZnH3r7wg9xa4z/C2
lHpJ23ewUJZj10IP/nr4fBRBO8spEIDazOyOtwS/SJYOlBEUlupnZxxxm9mN8Z0F
DwJ3xpy//jobjxg/jZhn7X+pphDEuaBUOUJNe6nTKUKm98r6JpDOZ4xTiOBWg9NI
trATj09HKNZmTEyNWv099oUcropWpU+6bHP7hDhi1x0umbbsrwNnJRR07+OHbzax
XNhXKBRrU3yDyJTUvWDuw82tvdIshq9H8aWQZlbw9B95vOC09TShzfCna6peAlfv
LQl/2wEFHBakP5dBvEnemNj68EFoxdqaZgdY7OLv8mYXKV3rvvGx0RIvlzKQl1DP
xnbKOFlyx6skx1yPHdEIqT+oCNmsV4CRxxTMAjUCBrHUa1ZC5XRYCMm7QEB7woX5
IqK9x3wX6aTcbK4O59r5rJqNIUDh/aPcm2APN/oZZ2HyPE7T8kzOklQjLhE9UmL+
f5yur4fZBsdLGZfmV851HPHqXv8B9OF85orkiwDdQQUb1ObyxKooynafzn1WrEsd
W+Jm16NPrGqT0XF+f5HK5brXrGGyn6lG05EDyVbRy3ep3hA9sq7A/o32d5TIpw1L
7/3MR8ToR5qnh92ysJ6fpuHugEBJ+jYTF+U4QT4ZDSCoqatUIvgHV92Kacibw7y5
N67n1ath8zv0vSbO4nvaRnNflCP8rVsslxkZr+++2Zllr9xTIhqUQuJXjKVupvqv
xmeY9Om/p0HIFYMl0pCjgBXrIecfz5diJ1jYu8rLV1fkQJSQyD9yr70WgIWfG2Fv
6WxaFtxC7++m4/i2eVmpFr0hCje6s7fnlZDA6PqPP43JoTM+BI3xr7x+5BWT2CAC
OuxpOZU4QT5+waC2c5pgxwQthSsC7mEPRLwDSEUvESBUnM15HcuFoydaIfVNAjgS
DBsYw/7iKX1wX0IGOKs+dAVljrzSv7mQTongdBup59BEsFjKdJrXAOHtJoS4/zcx
6NdTeLxV8IhPqIiH2ZJ1R0e4z+xukl9qvywPYrIekcITBjK9XmPrVacecgE4Z2P5
U9KLHHzAXjg1nNrBas4e9ISB/rGMYWwa4KeaIGnP67sYWqJZVPKFNYXchwv8BlF5
LmTY7znPH9D9G1Z7CHEAj3OTqZT5nTX7BJYv9ZhYdb84UhZtRQeb8VK+Y3CEA8iU
UJDmkOM0na68U++l2emR049Z0PEy46l3RqhNnae3c1TRChGNMKZIAj5sQC+ANwsX
pQw5uIQzXEbmpryEGP9xFCMFElv3G5I+4y4CyDdCOlRt6PE9603V5xsTzoVJAsXV
ElnsD7OycieM0fBspj3qsFB3ujoEPWfXJhAUmriKHkgtOXfCGswSd2GMYzklf04S
EFhtJbvrFU1GyK7CMFZZiGUH1TdNDE24V+qYU/yMaWcx3Cg1INzumXcvia7Rjnwl
P5DqYIf8l7ff5gdbZIH/wiSs/oyJvKJp9JozDzd7FqzWTv1Pa298UrDXEhKg6+cW
8FI42ZU32oXtz2jsn85EAZvKTtCaHJwg6CrTe3BhBsyiFR0agUAlD2ZD9Nw2/Fzt
4jHF3t2n6set4qbqqlndssYUnZrOn7qyb4zCW/C5ARtT+1WXu2m7xNHmF+ZiFmlz
6PtfYrDYpWRrzoB4IQu4xI9yW1iFAQFGwABjwLj5COz/PST6xlC1k6/eBrZOf7PF
UDMBH1bUXNNiUU38EslD9K69B5qP8QVtX3+0RB292QfJKaw9VXi+xGQQirQkFIQJ
MZ1kvZQUlaRwgW0Gg6uCOclln5Xoay7zLPtC6hxNefe0X753XprQpmVbu9b5AOXF
71h6dZ2N7B84nC+7kcWH6qOK8AIrAhp3uOMyjmjUiac6vb8LFoKkIe7U/oqaTotJ
BHeoSLUPMIr2/50UfpCLEjXqN9uAzgKMZfVRwCCK/uTHm6/r2ZlbIwMQLjPU9FUu
QpoNMZT0x/OV7Cd/BXSpqMUbyOfKcKcl4T1/jih3CV8y8u6V3Zu79OHN0mtO1eJ4
psuKeS3xzZE3XXWf5fGoumwPyBZ9DtXg4E34SIQwcXcJOjw9ZTf4D4fTIiUibC0x
X27j1eqMxtwqJK4pAUlOc2rDyMjRfmC88Yn/Q09Ot+QUrEAEhtDz706o28uSc0dH
4vZ+Jj4H4ifOBIqrjyELuSTfZkoC5ogg0wnRN8s5y0CUjP/k116dh/HYGdu+XDta
bi4jVk4IK8a1SOp4zGZyHKPz5gF/DErv82DEJSvGnuce5UZsWZpv+CkeSTji1d2K
pJI1ta0eT7+UwFonQ9eKL3p6bBlH8b38ZiU1W9UzZ8R0b36qy1qov7FnXe5evnYm
YDP1Q33UTazhvT76eUg2UxJn5wUOSbMmNzP1FJlPrbdQTlzRtFYAwXHVeh2lF4so
2kZz3+PtzRkm98MYhg6wyW8JIaNGHzuidtrnnpla5Ajuk5wPP4lhARtcv50JqQAZ
e/K5DWO36nnwTG0WBfh0Qohf8Y4uWXBo/hl58nrOWc/1OEVfqoNqxZvzAf9GuNsI
6WH80oy2YI4KFzZ+/uhHroE6ctLwRcnn9HTLGPbbJwqtyxPJWx4exUlMqpkNPT6v
3BdMLAiG9NIrASH5oM8e4k0KF0ggaQa8haL8Y2BiTR5kOf6gIoUKfmV4uy99HBvZ
/gSv3B9gP4X6sVzNNjEB/x5XfyFQqvW4CCKmaCiLsnSsddYleVm9eDQt04B9NfHS
C/7uQUZkAu9rMLPfFoWUEPMEJ1YqYGbJ2us+SdowT/UD5OaYuwSLPTgCEGrSV5f6
kYX1O0RQLEt4+yv478S8Hby6UVGdHP8fIGCHhKcbdE1TwV4ohp519KUUuxXgbB3w
5ekln7jwhtM+ifcNsTz9sgtpN/pojARtpFJ0oOKS+pLMEHLTShCb5LV+ByzRgdKQ
UgKLK0tUleFw2gZbgs3Ol9tnv8eMcOGJLa4eZTyKlfNzHOnjCUx5tHF6Z53uFviB
0Ylf+NykJMx3/35wc5pQ/XGk/LgqU38irRv6LJgNOdC3jD9LK5jZZgBKcbiRfV6q
lfOyss4bHe/D7F9UsEcJW2depXJeLr2f6aCA4zNTs2PlgXb1gmJ8pmdlxMrKrLcw
T/YETrCyfZztXMvQB6ykwKifJviow7zTc09XvVsmzYkvVlBH+18XtnL0fWgiNoqN
/H3Tpj2P6uMvw/9Ovsd5I8YyY9AnBOm/QtIWgoHxnkTRiRYV5bAs1N8tNEEljXxB
zyGrbTufMJyGnS5N3zSgPI9I4hPe+N52am/3ZD0T97Tu87f0VNCmjhDz368owcjT
aLGhxbbYXEUAt+Oq5oJJZlZDZ32qtC/OAOc6nyGRhrhbtwsrCPbByoXUBAAEyNN3
+Nu81OlsFISvOvBJd5YKLGKhv/2+Oe5N5qYee/3Qu4W9eUilYMNBK3CVZ/qNQ9Af
DLTNrN2pLwwUnIb9ehkMJWrZKGO1/PbkQPsoQdst3yHPBG2d9SW366LYidThGHFA
hYwfDZ5Nan36AeoZdeWGPlRNHWv25SZFBUe30LyXNJQA6hHzhKLDYDh4dI6OYsKZ
Ca8dWkcpHRGSAj783h/+nnrCBjjQVnYjJxRHbiR7FDtZSqtuFiHTVQ6E3phEAI6k
u+K+K0KPXjpMVFPPMO3widoih3l181XABbKSY+6n3hhMxuhYvFcMcjcUVDdZAUlG
ZsfFsYa3JtXKtuaoRO2D1n1VLvr1VMgThxkrlp2w1Wh80hWFF9/rHvgn4q0BxIGW
DDh76zRHscCbwulBVQ3PNcl6PEMeftd+8tbeLhFJhmXek1RXIiiGBOYZw9Lf6OOZ
qVzYzA82+/v+id5Xu9F+h/FYoqEtSMo5gZ7vInCt2vzATtMZ6uYjCoylQTHRxJyk
obt91LFhtthKjJWHdiY+MT1/U5fXVn+zd/nsJQai4mWROmDJMV/Cw8qxvmMX2RyR
r9+SIokYb1VXhLBANx040dH+LbW3NKITVeeVWYmix4xhCebYjJ2Ikrk+IMnhypQn
ImtQHCx6wSBv3ZgsppW4C+t1qzZeFba0dOGOHjJrMFturcyDtGn5tMGSRIuk+DTL
03ApzTofMsHI4cTw3CCE+vCHMiysaUm4iv8dEiIhgOmpuGJGDJyWIhZVoIIVv8Fa
vdobZEt33m5fusAnrUBJXVmPqDKq7ZPoY+TRu5XWoz+2DJlMBNnAhBnSpSedhiIM
4B7hT88DLZGgss4CmBJPvP8H4+35ANULvvQh6NZuhtvzkqd3oSc9PUfe8W0jLOg9
pghoMZOieqBWREL+WJQQxDnsm+B3ToPouAO88b3MOwAO1mXLfBNsM+0XsK4AsUA3
5/+IuLEji12ZZ0mYF7kSU+Ji8T7n+T1ec97qY9Uz1tBtpPFSdfth4f/0hCtINkj/
MofQkD0LQpwxeJfhESLgA54SMcAPGxnSeYuQNqjsIeFm3EovhJWIyRTpQjVFeFYQ
CYNDqOP1g/VecBBv7QIac1DRx1d0tK3xNeixP4UQDx49vCn2G0a6HjHCfOOh3Ad+
T4wIjyM6MZKZrl2QWXMLY3kgIlBRDFqFybtKiBLoZl57R/TZu0jtql0MHt8kGtTz
TOMEJks3G+2qe1XEMkOBXJH/AegCyHjDQ6GSkkD3kyHlDIFmGYmSfj/QMVGlrPDx
oXaCbpEfj116QjS1vOWEr4yatE66KUukgoX4RySsaxJSAI8GQQc9Wni8PkaN1DbG
yOamRo9uJL1vNjZBnNziw3uEWYCHzXAldJVClmEspdbDYdtfeFIHjr5vK0B4e+AD
7m6nEeTSYpC6zYgllQ4M3JO4CptJhQ5In/QVoRAyXmolGLaMIiyGzYfD8P3S49Q/
1s3ZYqi+Qtd4GU6D9H+NSGrdVC9ThPpyfVNv6RN8Gf7OJU/XE0fZMfWhTn+AZu6T
KXzJ+PEJ6zEOpurv6BS93pHpK3aQGrdD8Kn9EkI6xLVpxqspo8068eGcAuB74oR4
/F3G4CWFJ6OWdVLmFDEEfa/2BEBjdAjI3H2Vb2yghaFIF13o05EwA4XljQncDQnM
Y8tVbgKbJRXDFLN32nG4zK9u6NJR0c2glQOS5nFstFiakRSbn1yxQ4YV6Tr89Fx8
vYVz7xPE5ppW3+S2AzGSjbErwITA/FBiHI8kkU2P0/qnWUO7JFY8Tn9g0T9EguZI
wYvdMOG5uGMYnimWAn49Y1COd4QG7XPyVfwnG/V/c6pkhKy8gJhPcX2onvVPiwxw
fgMqbYAbHX90cIkJ9DIA38Si8Z+FTVC/GGqqf/7Wyy17v76SR2GcGux8dEQ/XmPM
FdId1hq5rOugOiGhBZyoWGfMSRFOgDWJ0RUv1nBXcCscEE+GJ20822+3715+bEVj
1UlPoFps+HENK3eB35pJHmg69aiFcf1m8ozZnKvh/PsY/XfbjrHE2pOkGj2wF/Wc
HRDJo9XFadred4g3b2K83fPJVb8GL45NcnGY4x7gHUSPjlxW6x3I5Z6W25aFGrwI
BtYu/N1Tq46dOA8j4LQ+Of4EDuw5Ofa0WyoOMFMrhEYFSnIeKWnhFKV+tilqDQMK
olxaQjcNmzti98lZZu8LGhzG7Q+u/lMfRSouu4ltqw5RZ4Bp9VS+9l0O6n34tYBP
bWLSiD8oGJUQMg9PDXP6Orceqrw072sE0qZv5B+XN997oawirkrVNgEBM8ohsMHn
82pFv0IlCQq52vyJZ0p/lbNcUg4x0rA1GXifqe2Vi1H+ST+j811cbjHENHFuoBZJ
rzCf3Wo36BGSsMJemL4jS9xcFEpbVAZVgVq3k3FdW4WOzcvvaT5GWBbtISmswH6I
XlydcL0/AkkDN/bInFAGI2ezKQXG1TA+GXnf7DegoS1+eR90psbEmHE6pl3OHHZ0
sDRxSEb+WlZx4lN+aYj56VdmuCRKEyGYOP0rUycF1YSxYlZbCNYFTAhbW5yUIIKg
hMuzyYOjU5UWhd8cIPHNunLPBonhIBWa8DJBgwTNkF88/3qKD2uBw7nyq8h5e/0Q
WMDs2Keh7IXf0jZc9bY+SidxMXpmjdVjfi32Z+3/pQ8oiVT653rWKL+k228lrUxv
CWuLy6x0QDi2ji1hCLe1Hhxyr7PSywdVvptigwFG73szYCdWdW8FpIeTpuIT3ihP
6dCM4erhakpMrgyabFZh4geh1a4XpVrcNPkHMbHLm+wTsYBv5346/7SHclmmSEDD
VObpE1JqgeIb/njE7u/VkZGWSHQ4KUSstPJAO8+3nxokmQxE/t3sqkNVdClbcYnd
yaDh8Lz/bTgDbaz9iYTN9awmbz4XgBRl7xtPt6y5dVUOQDkzl41P0NVQ9xpTp7+2
ZaExlz7JMeluEr/zLMq6hpvge+iSo/Bf1INEODUHpsXBtTMGJaukjb3eNY7dPbDX
73c0Zrr9ZZStV8silqB+ihBsewoCUH20GRib+gP/O0i6Td9xEYecOmwf4X58JUfS
WauuYsg8TSwWoNnMeeRFLsf0LXvqHuzVwJGrUQpUiJTBDeBPSNvUsUTA86bjzzFs
3MM5SujY1lwZ6vAh7yEnBeMkOYrkCsFTQqOJjRGxaMUPl47zs1CWsRoAdBfsUIkk
WhnTSTyrk8akjZypZAszmuXbhIoMatGoeayHBOCtuRUyXyb47/UrUglGAqhkD4op
PurjAeNphAKmZSVqeGtDd9xe0MfIBTcSajjkPqvN4ZNCTeoEECkJEXV3Ljncm08n
ZtK6ez+jHdwwgysf+3tdjjXVkN4D6nehNiSPr5AXp042z0HfPqaC1hl3zqF6FPX9
KiMB0h2bK9L4bhvOWQQhKQE7XwROv1UPInJK0FQy+BgNBd28aKh0PKPfIlSil34n
NCjJrch/ca1at0d4YWrCip+ckyM8mKhpivfh5yepS+N//VhsWdYj7jF1COsbCZV1
x5tuZFRS9tYGfy/eEWnm74v6gWHZube2MMcYbIMvPFMa1Ov52qVixh2wCi6iKuXH
MhuoMcLMi+983u6nzxWmUpCUWbWXMtflmf5aCLdR50Z4pq0LxPVma3oRaXlxe/QP
gI+6U5LdczRl24XPcHX8ByR543t+d1VTR9G+5E7WnZofXqWInmlnA3UPsY413kuE
dKCp//A1crEryGWdrrHT15Ug4panmScqgM6PT1WvTH7mV/zoxomu2tU/7GIaH0GD
iRmeswwDpn/qwrTsNnudBNedqXAMLe2ITRfjrztFi6U060Jv2RzGOhUf5ROK+ZZw
Y9K5eli7L7Cqv0/fyW2scxyiM2GSw5m9lvuOwJFLwszDz5nO7Zy/787onOiqN6Ks
SFjeW2hsH7YledQ+EkH1VV5RzA/WAuYZOPXnLc1x1EslJp6q0gOANJbXDSy+8484
+V3ePeRfkms7XLTY3q/POGICuv8fbkJs4egWGneLWZ2axHVXzKSkiZsjgmTZTK+p
sIsDwvxukxXYTsECT4Cqu4gIgS70519eJHwqa4CG6LiGk23CDavm4IOHCWkK2RON
X+zqf67QF8jF9zutev/2yXVYj9Zn+D+w1xZKHZhr4CFV9rc0TFEBAM8l+Ntc7gG6
IyKf/BwuvyiqLA9oSmzKajnEvywFcT6rvFg/dXph32LShVaN6WDaauIUug0DxoXE
6mTCNSOkUZk0O5gassSA5Xvxbqo/kVwbw+MRoI2g5FyVnDs1wQWVnVEx3kWb8QTP
YuS57Y+u5h4NgLIUacYJc0fVp9mofXWkJp0tuKvauymzvfPz3hiGPMEB6c0dwDne
80fiZYm4tEsYx8v9tdpuRXhztcy4j0+YpiGwb2yuJXlYy+Voeb7auW+qgsW0ny4P
Y9yN48RuKYYnO2RBg7LpQEUFDiaafU9fCe1f0F8jCShMQebX7fPAeDW0ESPXdN7e
3ASGd64Ympx3iuk2wMqrA22wsubGK8GBE0GalJLEOl3IciU4vvYAjHpUwSqECO7I
7IXlGMDhDnOwXyGJ7ps9RInq2mhqXfN40kLJt3WPIEmHKqE9Nggu1SyfaaenFxjs
AzkSKMGLRmaaJ8NuP4Hx9ktpT9R51Zjib+h0AJyROITzXMLPwklsksDb56k9cbcx
yV4JgO5SlsFzS8sM2yrFgZA9eo+90hn5OjXuZvSBFzkgSfn9Lsn0bTz2KeRuCzIb
mZnsb/I7zcHfWg4PSwj5kF/OxUFhZ2RwKJhGrZ/x5zTTPdj4qqkjh+MeawJPLc+h
k1lAQdjNpROUg53rMnqFrFHfCdOCYW5x02JP15JYGhvUrCfDeeMaH45Iumnmus3/
z0BIcQSOHP+h+b4YoxVQWKMCoDBi24EvNdieZNifU9ysdMutvAgrfOZBiUBd0Mdj
IKsNF6XwRQJUaRhgpEsLsMQWO9MvRzUWXcuQr/xYk4KIxRIzCzQcliVuPrPL9HOx
1r8NcO0+jCiIZHlCEOEEfKOW/ud6/H8eMIvFX9VTWqUUx33dTSzTnfH/R0s4AVpk
91WEPm5UcNqX3imGF2w/xdBu3GF8ojK0Jay3/8sKyRHtgHH6n+IiQpu0/jnXiB/p
m96skFB2YclkTb+hgQHWDWNxjnfjOgQL1quyOBH4gI1eTsGqKWL1L/XGpp7tXDXI
ZcCMFaxda42I2bd/P4g5G0AbLVr/sO+3HhppG22014oNd6CcU3UK+C4PKuR1++SH
oPtJVy4P5iRQCoGIxp/EyNyA5u8NeQeOyFZvd8+7QQptJ1RKukrlpPtOj9XiUdsM
Efg0aO2MaDpgSd/kEBiSQ19n9OFbHjzQV2f1ZCuo1tJSBabGYHN6qClICD6qq0QK
3iJ4iqzURCOHjHy0K0NhR3tGZYBYAH/1jTFP/p659f9pY9vK/y5y9sHYG/6xV2E2
VJPS4iz1s086s+Abi4qB+aqRhVstknNmH1NlXDJlwVnfI/fZp3vHW4/wqby8M4Sm
05Y86ayV+PDsronxKr2e22u07nBYSExBDFJXt90LUcuKxIJ5KGL3ljaulUZCugbC
nj9qJ9y7LDJyKYQb2cT6DTYpeJfoF+g96fTI6isilnoZjrJtQV274LdKzUTg03T0
h3zcaoa/jXX5ZYdfuhtortxL/Mw6OmpGmQU1wow2f9thUIbBx9wDc3K6+k5RgNWu
S/WouSQpJ9WK/QXocN14U1GBwhSfdI/S/+cm5xy6X6LtxQ0a7n560ZaXkkOEOIV2
OyejQXfEbF99cyXhrM85v7HFjgNBXeFIiBJxuK/4ORl+Kf3qtoFyfvtXPp8eTHC0
j3Ed3eCroiXBHraXRus+I7Vmgsrysg1H/NxyQkp5h24BNUAcCPpwryK0OUfpB0OJ
KenBfPBQKQIUOnaCy2RMSqizISxCFIBXmeyAFioJIqcWrh/Vv277sgv7zJWS4gKA
H+CY1/eUcDd1OlIGug9js8KasMfIA7gKwBJWEVCu49PAtb7GxzN/wgxAdarFOPNF
gzGHN+RdLJqlq3VhNmfdDVOYDt/88gwCLCkOUKbEngAmwm8uiYfFsPNsqEUBHkxF
gup75NyXQmkcJ5Rvb1cN9d4he4xoMSseUXWMZDZ1mDXaEwyUx3zFCaoNJGcBUpa+
yt8uzQEZ3lZKdrRN7n6m7LNdIq03+n8cCL1cXgx+EeTOZ4wpskJSY7A8JgZofc6V
swk9p+Fg9YpzDSpa9GYbyT1JVXl4uOX9eOh3Yca7TdmFxyC36pNAnbr92Y0C/AOK
Yx2djyT3wqkbq0341nxLnywKBddwxoCW1PEsZdbSThHoNNY++tGEBrEtcwhe9Ocv
+bEPmjshrbZpajgzcXr3SPNGvgJbTa/gYQScF9aYn/ramzSA4WWBLP1mNHelT1XO
7xyZkcDnqRfSqvry9jUjysLsf7u+lfACrW7ajOMT7xd8fLfWHWBAV/HJIV5V2kLf
dOix3gqPUhxvOM/lSkNYUzZXgWFf4ix/IixlScj4AeoNgB/pwfmSThh2/0lc0BBT
R4qVIADN0Ib922lgPUcu/4cMUuqgDGfGhBISbML4uMQDEZcOcBMJqHF/qoEfO+gR
UGpHnrfn/YJVOV75UZ14BTIifHzZk25qydoWmJ4D6d62RhbFsGeIrHo93GkW5E7J
0Jp66EjOy0kq8F/RknwhEV6vo6lq1rHRbc2qyhSpd4jcO+symlUgeaN6MhSEVePE
Pq8dtuC3OnSqW6MVDPUDTBYbEcLTZH4UfkOAp/netp30NsMT7Ok0H3gjXWfknOIU
mOjKUu0doIErtdaRpObv6XgrBNIRRd+Ee/ef54UPG/mzoaoomQubFsKVU1iG/xZ3
5eiIZYVfMvRIuao2KK91Rmufk8UqqIq/yNAAPFQSHBpXgM/2f7XZ1dPqdJbNCAMM
dn/Ge9aulIIrZuD/vt9VGh4G7kdwynNECyUDyULOLD2pAEQsw9Ap7um0jXRkVZUs
ucTCmmp3aMRhcLqHKzYYrfcCkwe6Qfr6jPnN6Xs7LlWkjsc//RjevsmASR7kMPry
VOL98t6Q1kWzTXeZ6w03HL5kX7G66czVReUZd0uIbjWBXGnexzV/g/2Gj67xB74I
AJTqwqDAOIrCYcEnpnBWFIcaNQ1883MDQt5eTiLxjW0f6Sy0qK8H/YUSAuuIP9vr
0oRPP5avOMyiOSib52Htaw7JUv29NrLgpLc99X9HE8hWSsHyOnD+2lIzKIAe/5+p
bxVlIYB95K1EFduMmDwD9pYSLaUrh6DVPRBvcGcv1Wukl3XmCvwNJCo2p48a5upC
M0OiG/6t+hwVPyVSxAI9INisTqrS0ZmBsCtrvxSxXpM+lMGs9YseFCIcAn0qF9nU
hWy1hwE6hH13f3bMNmfGtpPpTBBpCu9slnM792G/5lNsmI9m7Ly5O8rxrQT+STs8
Kf0Ofs34b7Ac1SlLl4+/SXwUDt0NI7CVxLmPyILC5Hr0iparWPvBsRGhuwXme3tj
YT6UhnLoIOxij5hG6Ytn4XaOCuzQmMRufyR3uemZ/mfNy0MDT2jFTIC91zpWwwQS
WOIgDkHxz4axd2ae7OQBQpY7X+kdLkrzUIJhG0o+6vtQFfHCVxlYNEvWC6HyAZJV
w0QQfVgwrryVnySwjwkD6s2HV8SXWLu3MzrKmIjzQDrI2v1BB5RkHVPqwobFrW0S
Pt1zdZl1CJU1CauXOfA6cq8tPryKp9ZlHS4G533giVoi08h87uAjuBEByfn205q1
NLnJjrhjHWMRwzuqyRApfmGLcQxdxZ7uU6a33fVMkwnQT/YKOqoTHM+7naijD6ot
JKpNAUBnSyGWPN4kZ8Yt6Ac8yk4kIj5U/2pSs23WDEdq0Ah1R/aKIXK/PpcxF9Hb
VE8MS5PzdPRwmM+Trcz7/wPOIIcrxKxMLeOuG3afX0yYtcPP5mBuNkNgpTk9cW2r
I+ADRw8zvW0Ls5ArCagJJTqSyGYC5gywp67AfZbXexBloHtYZ5PQQ1Fxv5ELzh9f
f8SJXwGnBYC5skV/YHDayHD1wixAsTgWy7/RluOcl+WiShu7gZf3Ekfb6+P2HYLc
StqZdXg+86I1hYn2gk52eMaY4cs0mLAN0bUnea/T3vxzi4nn7nOZoxdmHNxKtniS
UbAafKIwjBm5njB91/VCtPztrql8DF/Ak+A2JsSUAVfh+w/YwcTXULxM5faZ+NUJ
SE6Tqw6Lh20/6X4jVwhBHrO++VewBwDpdtIE9iU0xV1Ja8QQKzFhbJrEv9LN6I0s
5Qv+lgNwSZPjR9hfPodnVX/nQxiCX7NZj9zdB+LJbbDD3CsBxAUWM40JWOLAhX3P
bfbp1RurM6/fqNlTnEnb1EgBuIKTF3Ih0CZh9Q5W+YItTGHHYXlNKpo/6qSIdRp/
9CxjuuLA+DgjtSWCxKNKqWqX6Xj4bLFM4BjNPP/4Q9aufYF6/trTojTMglyQrrgs
Goig8rg6kKojEku3SK2Ogkzjb1JPTszngLgFjvI4uDYTou3zL/YmbDWfe7qgf2Ye
KYsGyqC02NeRZ5DJ/zd8kkIv+Nx6ymMK2DRejuiyjr6DdMbq0U4hRcVXc01AqUIL
QtA0pVww1KAPJlYcZIpZSjVPK5IZQ6RX/Kf1XuSxQUqzH7DJGIACUSxi7rmXFc8V
cLT7nfVFA90jKgCtJzIAqU8nzr8Hy5ft/g0uC/TGME6IKFU/QrF7RQ5ByrstU7VA
583QWgPn+8w5paSKzn6DrqzHlNZTxa1DI2I/1zB879ibRedXxVRvON6nxs4YF7Sw
4AH6HGua6T0AlhjLeNZ5LiIQa7UiK0QI4yGxDWZRs4KST4zaIhQIhHQj375T+lwS
oGIC15bFMItAolE+/7JV6rtVKPu+EDMuEBMCqHU48BW4U+DVsJoNaCKSd8Yd6Fqi
CRlru1S6pKal+prt8tgWZHFu7B5/KtT0aKfmaloxcJCpx/ohTNHgEwlNi1Mnavs6
ceS6+2spEtKq9226VMyVTKjAfwqAKOy6pOMjCMjzI6td488zvz1OeWP1G129vEUf
HCNlsj4Mo3/ZiV1lhs90+ifNGhcF33S69GZiFcp6IjMr8nGYZbjpRqBF2wtHyG7H
hDevOm+sWr0HV9JzRM5U8XVGvb2femm1HQoJvtEHxfoY12NWjbE1t6mo/LjNOTPv
AljsKCcEwMd485L3NVu2i0oAU/qvLRRXbhL6htG2KHy1pKCxERfcWELXI3a+D9N/
bWwlMME7MD/bLGn8ayOGBCkR6A0hzrrz3xshy8pf/DyZzGzCb6r5JmbhncvZI/hb
VTI7Fxtzl7VF49JykjWtGAV/gGrX+usi44MYSNthQOptdD3YwaXEpFzewBAhGNwT
+RUPF6E5tPWb2L7M1ydxXMRAFc+GheZxk4VpKlUhafW8XR/7etB/KFsIRu4N/88S
MZT0FOfsKLyXOyH/tGt83A7HyChRbpEcph5AukWF+gAgo1mlA1xS14LDvIAhkh7Z
Ei8Fb6yX0z9E/6LxwwGT+KuejyL8HF6MNX3pFxGBVYg97RB+tPiFoLo8Xuk24dEn
ASCzbLJtTWPUzvAjYkGxC43umpWpyhrD5r4EJEp+enUxNvBDBO0a7StQBGjh8b4+
KAeWZYYTK309RC3qwG8TV8ADOeyFtXU0Z9NlRilfMHwmxFUXHaTRgxZxIbLEgcsg
hHACKCY8UkZeG7g1oKwmUEi0zIUevy6QiROhidi53c7BDjDBgU+H5tmGGLmODHsz
z4HhDlDOVLRWGN9qv8jY9vGqznpsN8hzqNKe28PIoxXzAFc28Yr0Zysp2Qlyjl8N
YqQKFQJ1AcYuqhJ/nlCFLhLilMF+iFgPXdVllsM9dMvJeCsBnoNVY5iTAWTLC2kb
VZfEzWppc4lzIpmQj9aG1GkPlT2eAn8LhRP4XROokY1jVEg9vpB3i5vC+pudbPwD
N93ppdvtgXDGwhlIVhBUQp5mxetyUlK1m8XcId/7iKDv3qye6kz7yqiYUUru6lnt
QCzINKYHHDJ0HyY4BCvYo81Ot2BRhb8OiLRWyAw9RcRt2ocIFwth7M/LQyTwg2Yz
lkDcCgZZLLu7Tgsj/MnxHm6O0N7ydi6Mas2OKnzrvgj5x1aNUoXHCXB78or4pf4l
WC4HIFdvauCXAO9toCP/LdD/p5jml1JEuYldv12dGg+7baLvt8n3Kod5c8eUvBZX
Ipm29YemXICARm51qD1WjESpRwo8CmX3fNCaPzfMpUiq2E1cT33DZ/za9rKba/zd
S2A9VBZKoq1Vg4ux4fehdh1v0zJQPRiUOJueKeoNnALaDlA6dqs0ph93k1uh7XA+
CMGsaRtXBrDyIFllI76/IB6yfXJ2/ze81A4Xl6jM+jPQnBA/XmEptnWcoJsJUFre
5G4O32AZEobCuIyeIsXhMSCPh8KLKuWC53o0atQ6TFzzLrRvM1FoGJsxMJQj5pTo
+fqE9+LiBRaGgeeWxfOjFWyurWXMBRtVZD2hvanKst1LO3FrWFrL0sBiDrYAMf3b
ItY1+LEy17K68WCOKGt7CzXk7Vs8PhS66bCynsbACFf+o3XmPVIsYSzulB1DHZby
wdF8uPjW5jnW7yzNDBFkByqE2laH3kySSXLxrKjoQNEaAP5mF6tCrwvdyHR+fGYh
AtvkD9dX2gIDsfQupmn0IZEzJ1CvjLQp2/CgHclFsguSVpO7jTuoIzByBmCcAbE+
v3D6oQJkIJzcd5hmxM57fJSNTn18DfSIzLKtqeGkw1eGX6G5E/g+VE/2uMC/8uQi
/FW0K1mZMFESPsn6pEkz/LWukork2ZZPtBSU7ktrRIKrix7yVtT1w3Oj9ZG8yXmv
MtPBC77XlIF36K9zfefp8bFimwWM+4YuUT3XzWxgxWrFnk98ZHbvUmZ1pYcYPdU7
ri6kY0xI7dSdQsvU4trdYzs/g3KmVsZrfe1EKpejSzmoJbF+ugjQXtIkBnRcrZa8
81cPJ+chKf0JKHYrPNx1S4VXyBEluSTHxmORvaypfJyPpZ5CUA9yewhWV9r72Se5
g99kIKH+ZK31BZuDtwrJShn3CHauyET5uRKqHACCZ3nVv7VSu5nemCrt9oKSP+xg
PbUjxwlGn2z1GIp9fT6vGpjqW64yNdhv0Jr1lrkQ0TsUXE20Nau1b6b5MJhYjOc/
Fij7Qg1oxOmZGqK/Bmwu6AieopsxrOUxF/ef7KyqlGrCktUpSjSGJ93c8cJFGAm4
d6iPqZIVzMbsRjRslrvmnReH2OAY9yHjxGE0XIIR9uyl6r3OnNXBplIkNkIuAXJ2
t5WkgN6+bND80Ws9PbbFiuuAD4jX7WQ3olGibE8UByEDd9MYxbaXgoMYK81mNMXu
FRBglTPU73WniONGeOdZiot8+l8yQS5k1EQjixncp6Mo14V0il2V3BbHOZt1AKp0
e1jP+52M5f+AmG2oIhYDSDBdoQN0RpG+5J3Q1Agm+edNMLQCdllnf1HYijKFpWtf
DKqF29z5NyHOq8NwwiXKDS12+AZuJcGu5zqVFerRrG0QdJa0V5sGal6TpNtba+z2
ZyBb+krfN3yRn6hgzWVFten8N3O7NwItGruJpQ3VJhmXvkmCE39vJrtuMkGNzytN
cboqXyQmt7GwBijsuXBQoZ+MteOIkSPvMH0bJKZelyAY9u+apORJFag8SOjC3cuD
fvK76hJIxXJoYAAcKHDIOaJosDQ2fNj41UasPUu5PQS3f/qFN2IJnNt2qgUyG6WJ
3hYZwHjSWeuOhW8tkGPpREensEMC4ZVPlOr2wUP+1rSQJtPb8NQPtSGrK26myyIx
97VxlkdJax3LYRv2eunu2Fx9m3rfnE5XOVpmllgtreRd/V8qs50YcYOlnrW12wpU
OnVRpkATYMV/xK8Pm3mn2XmsGZyXJZIwRiiRIe9lKHw6Fao6GkWEJ4ryLkDGlCSC
4uByuerUiBuX5IVFa5mTL+CqKF7yvJcabk4arh2IeoLjl012aNGyi/s2JV9h6FCQ
2Q9dBLAsXltmLfsxx6gL5vcKf7TYHwr/+7HfinFa/2cqr210zlRuFL7JwmNX6OVq
XZt6GrGeSEoyz/WBDuExMjYUxdctMLDFN+m3l68blgYH5UeWnkKir+DKlgqUWEIo
n/G8Ol2OWf799NO9W8W9VZ7+JROPjugPo4+76U7e1Eo+VXrReJ+doVW0IEIZ2JT4
yREEkfam3XhUoGfQsFv3HVxuur3NOg7jNyeIqpj0NzUibXEBs+56gKcaPZwdMYt4
Ofpq+g2WIaBZ+ynJKiBKcQZs66j5Dg8zVpEUigh67VV0ovn/Ae1unHZG/rAUvKzz
Ma38E81eabby0p0ZXXUWmOhpV6AdY+DxjmWNQ6fRbeBACbFt54f4ydJ2i4UWV1I2
J89BPzQ8AIDQ1Od/P0BVpgu42KifC6mhwlmEdgcCPNzS8KR71TJjFC4uMpYc28ta
pcWYVu9Ei+aGY9O6cYSrZ/emIoxEnXiOTi0KeZrMw3cKqjhK+BdMCXDMetdXABGY
kkYoykyEorGiGYJtlWyCRsdiH7MyGELkC+eedpH6mAhWuK5p2m7roFKFtUGa++Zl
OTtW62xBOw8GFEVg51Bb4ghh3Ah6VrC2oiU7rlTcApVDI9imMysXGG0MMqCHe5TW
wwIjMnoQxfQ6I4mW84Lrz7fjcZZUF44YrPXZHF94XT4ozYAZSAtNNe11Cro4tbB0
Lp1QzpCGIK8cGkB/aQ6jQDGz06yIPE55AlGX+VyL4UveaNuwkIAVBAt8hLYffJxN
6K0xHqY7svEf7LApcZ22n82XrxmKnGBiymMbHYuH9MsYMp2orxDWozAZCtX6TY6D
Mplp0Jo1jxlPt1vqlc4+9NvTrzAkS8XqGIzJktbLS1jp8JbdPUpB9uB034DmMmog
2qSNetpt6vAfygArWXzVuzcwbDu98A+srCRfUUYxTX6oQSfUs2bxVwdq0Ch5LWa0
RLUyUTftraP9VaIMO7PwdXPofC0Bamb1EIQO1NAq423mDIF2d2OZiYKayd1ECvuY
KD2lUuCoYbOQe2HVvbCDZ2w9ftI0ldnm5i9knWNbMk8Y5pKMQwXHngGW8lGlsC+i
gM7y1TmsZ05O2L3KjvC47nJ6azDR0mUJW096J7TScVo9sKcsx1hGeUCz4D64LUeC
1XB0Zv+Ebz0ktuaVVCZX0sawPT27bywwBxktKAFIi8LKUqjZK0hNydxTr3Y1viNI
qDdlCm74PAg08UBQxjHnmHsFOXnOd0CIB0M7CAjIsWkyLSVnsGIL38bycQ/utZqw
a29o9cp12xvCo1tZKJ0gLqBbIul40hhiDFszc3tIrhhKSU018VLZ1Sgz9WPstN5i
a49Bo8LKkuMO7fB15lFlkVgfv+GauE6crfrgGyW6vjavjreFnrz8RUSWl9m2iWP1
wUpoYws+W7EDIGcyApMNLQDFpTkfeMvHPZfCNvD997DtERYceBruX78rRJipPV6z
RA5QGZ7HGOF0wOXOVlA3c9ouZ3QpxqY5lNXZ3YzdjDvpO7AKo/EM7tb42lxOUopw
ctOe+C3VN3CQj/sWvaLVuGEGjJHntz0R52Bb8KMTl6FfhudfqgehShhXmc2QiRqS
j0+dc8JCFra4RAbP9GFjBRvjBZPKrsYtyD3LOaRBr/6s+ikxzLjKk1thCZhlggOR
VLnnI/KPtEJ18VaUUcjOCjf6kHQ0ZWrxy9WKGo49v2IBU/t43abRB05uuxNaxTsF
NLo3JOdc2gTjJ/3wNvTjv7UT6HU1mw3sSSj2OFS2b0hby+nBrgRmGC14utBlfpH+
GdQQZD4TA/IILnGtnqBEL0n6P6JZ1Jjzwek+E69J83ScaXiKyN0M9Nkg+PQjaFIZ
Ck6K8URb83+8d0e5PlTvLOjIzURo4zyxhXofgaSObTJhPf08q7Q0+ES8gb4f08Mp
ZIRIDgjdUI2s9PAO41A7Nrx6jM4yByHPMucmcGaorxCp9rjWWaF+rJ19I5/D6GKp
Zw4abQEc9hSGCG/I/r37rLGH3iHiYhSStNM7m3klPA8A2h6qJum08wAjvvGksRIO
fLaAH41GpFisN5tZW+f7+gezn0CEJnqSc59KZKPK8eSiNpTrSlhb+3YKu7PE4990
M//wNnGz9jnCTHpfEACfMPcn4D2ThJwh0a+t2FZVT8L882jHyvnCsp6YoKrakbA/
ed9+lR69ZeZutM+hPETuTSPttZRVSTzM+AmEhCp2paKSqMbu4aTc1dTgmM0CTMwE
0vvnjYOSH58VEtSNzmlztjAAH9I+JQx0e/xPLevXV4OflQCqRWu85rdUHXRx6TI5
+5cvpWrjtTdE1XKu5MrzUyeMXs6jsq1D/VN7N8g1LDnIV618oB8JaEqFOu7jh3fe
SKTOD8ZpguG9yYs8p/qol5OQDcl0LELluCXPAqvgYl+5DVJd0lMjlHd+C07wHo7h
DEXlWfSZt2t5S++PQ5xLiPLAOt5syBPLKEO1Yh5pytKK3ppnvrwV5K+plkqC3e8s
Inb84WuBdE6wzPHbuTqRGwoWu3hYydIBnfHkAGfav4h0aaDdnUkLsuq/5FO8FKIa
djqHjSO4w62JKG2iKgfFOYQ6sPMV6mL5P36LpkqiIVS3FL33E0DVIUE8jDxX1MgD
4dnShCkQytAwLuXGw+Hcxz6Vjn+ZWV8+RNpawxDHjLgM4ipo7lltqLV8aUJvNHYH
4lfiGvA1yb0sh7BoymhhaNfeGdJWGzg0FMb3AOgGI2tSaPYY6gZoxMD7MTWjdd0a
FjPwwEXH6t4c1C0bRJk7hqxUDY0jbgYUvkfExWxl4+rT+amol6AuybRApZYsnRVm
G//9qMMEwx2sMUpRb2M6Yrf7hfsyAKb4wnkPZOUF/m3X4ZVj8scoCOZT2SG90Zyy
K29dN8h58vDpvYg0H2J2CHh8J7btQyi+WoFmuW98pDfHs+f+oAFkeQL1hTxzqHvm
8yhhLdyxDdLxzEekLI0s9xEXqFXBABiEUZyJhWK6XXbd3NDaw0xmXUNx1QpQ+ebn
LhxPE1Q+VFrVu5ZocESNpPKlokzzS+kXQOuweEPVQQL6H/icEP/8zeXf6erccEIU
yx6mAG57qPyJSFiZbKwC5aEZ+rdjDfnGNWGXU9Qh98vurqmisjpsUNLV8fZJSxNj
tYVlaKlMG/BFn+XxmA1CCz/0c1o4mSDvF6Wl2fIbNMB8bOoCR2BlIB5spAmAhy1I
dqfzgfVFtA/sATjMWcGrLvDsUk28/WoJzvVw7IPP9DV88z833XIn0l0bOScmTyVG
sd+7g6rLdDMUrwKmHJI7JKFN74/ZY8OHEFMYmSznv6VbZgd7jju8AScdX6LvtdQk
eXXK8/koyYBt2TcdbqjvCroM1R4DFpVyqgaVjwOn+Jq6g+AbQg0jaEMfmc1CAeIv
9ZcTFZ05DgojZxhnD8KEQFz4drFbZoK17bOBXSLTFGEuzk43AUpL5smfENcOoUz1
mijUFLKLxwYGgTf3mM9TXiacDV2fW3ILOyEGxEixYBH3BJKtQijq97CWq13TWThu
Ena/wwbjcwT0zTNPHIwmD1hpfj0TcCq7x3IZgqIiqDvS1I/FaSAfn+9169ECbbGc
vruv5R2tQg1HN82lYbsS6Zn1O52Fmq593spdSGbN1rXpvfGn8/02nc3RiySKU4EA
a5lXWC732kTksz43Erl25OA6x2X7/aIa3O+WvU82LTpodzUloPQzwRj7kDfdQG4e
gbgY4RdXToBjYw+tXL/5s7KTfBrmkvISRYKdFyHDawgtF+McYJD9Hey0PklqezqH
EXazXNBWOiLgyn7Wb93xxZTFx1z7vKdLTBq6LLoFe1i1qUe2HUXu0Q7zqmvit2Hr
FySxsBIVPjoiNVn7U2eMtfDWMlgAREwnbKA4AwuTxJaE+6oxgsla9eBFRQQKtyHR
2HpYhmDYC6l+O5q1/4cwbE5c6ACCK1ehL3XClDmj1RmNpUG/sAlxL10NSx56RSZD
NqgII7nrIl00/0gaMHQSc4qWYcTIsxhOgCc4Y4kBtvthzWVi8IUw5jGxmdnu2YV/
5dvn7VQfqFFsEzxF1WQBx15YkquBuFqE42Y9DyfDObSLM4MJsRrDjL2tRUTiX44B
GA1uwBunYX+Ldh3RCq9bDoMa/1VWRt2qED53nDVt+ItFCoqxRsdeLQm+X21s7JdP
SYyexb3Fc7v3RSmWauJBstwXwX8+IGG2rEfs8VE5/RukntHdnCIhZh3k9NenfRiz
wClyk1lCxq6gL85QYZ0DW3U95rbd1JXIVGdITK8Ip7dd0MTLgg7yQunGC5s6KAia
ycHwVEPrWt4cxOPDy19HQGnL2KA2q4kuHUv+4A3fNl5u7qWsHwoUllVfXJCPSDzF
90hzrR0ktr9qVh9BrEbzHmMeipkSQnyCZTbyXZgnLxheY7GIhqbaiFyEgFBribYO
1pjYH+1JT+YZezp+A88XXVwLfvMOQQPtt9xn2flsUV7KEP8qcTiVZfLNGyIPcj0K
gJzgbd8PljWZ6wYJO7V+ybqbZ1Gnc+zGYnDVPtpuj4dHArpWX24oHJEGQvHTXoW0
dZ78cJWZakVicEe74YxwI1n48uifXxwsGnTGvQnf/ky8+1l9UDyf6vA1I+70zI1V
K7G7tYdL9n3nu/wQGMiU8I/wUm5V+rgzcS1d7N7o8f6rVHHk1iGAu56lBcycTmZ9
xx3RP9f//CW6fbzJ9w8TjqOiurIvEhRN2Ds8EdWbTbHZlEqGFD6Q5TJ+cxy0x67+
zKnSdhGrrQVsyXYtlZqbDO/OQXLCz/sMaVxUjcUjsXMvXptfcpixlJt9tZRz3V2c
t4mlAMmNjtlwB4xIaWqOM/8KgRcGOcMSUfNbQ7oll9PvGAgtxAQh1BPtSGOCWC5o
rZfUWmalL+Ox4Gkb28MJ+d5LtqbRSgoPpU5le629hCpWTpOlPQSldMpAWW8Q8qqT
xpkyFFP2+TjaegCJLBkBvlRHF7VlqMLem4ppW3mQXP2Mvzpj7j5+h71uIT5ydVP4
Ktajjv61yx4B/JMo3MllJhNbNlIBrG8bU7EzdiwBXMbAttY+dsq04dCvYW0QVK0+
Ej4z+I5qjIJPMl/C23JkEgbMjWkuq7UiBcAF22BccGuB3kRW4YFiWidwa9D9qE6l
eHHc65yJbizKLv+i0ZXH5Ric0Oe7JIvAZPe6i8KdEtXcSmlq11cFSI5KCMB6SvkW
aU0ZARNpXJaD8pesddv27WorRFLXWhg2+h50jWYRV76hz3pKAUX/ZQdjILcRTaWm
lDOxsDk+k5uow/4haLzYLwtOkWgSRzl7aN3Fs3p/FudYnTeIUz1JUZ1d1vBecwfR
h6V9ftw1ZfSyPDbP6y+Fl/hRH/6nPNoUxwaC3uEifMCS48VTU1pCzVK31P43okF+
joFbQ8J6xpPzQZOz6Sfh19h4Im2idWbASPaWMLjhD1rYx1PrWnqhs5O0inijWYR2
TGPzQhftWSe8LgvU/M9Bqo70/zkhquancGt2S7pzr2Kiiduon1IpsihoenPyidVv
/CoGfBy4ToSJKcbjCsiXOPSqD3WWyIX8SNP+WV523U5QdY6CbImruR2enwj3BhIK
Ww0zcYl3HPBJ+sJNvYSDhCOT7aS7XQIKcJ2T15o6c1LYoXwajgcFQvzq3O0MCFMu
fUXA7L0m7ZLCJhXfYIreNy25wsBhGh2O46367PZOmP+M5UsL8Imy90riUyDkKd0K
Z89Al2r32/kT61qFvCJ0w6sXtR+ybdLPoi5IxPlAplk1RdivbBq/sRbpofMwsYQF
EZXYOFgKzPlV6/2AF5F757ANx3/AbScJi7hEYFTv4s5LidLn3zEqoolQwS9enVAb
+Cwy3CkLKxhapTk1Dw7U2Inkgbrm8yIWEANVdksDcC33zMy8ksVdMtLQoAPmmKDG
zpGdGaTQ/P0USseC9v1sWxZoFoqXPA+MPjKyuE+Z89UErkf2VqlMe9f2Wz0iRdob
Slld6T61Mb6GTbkTly5nsuiv9rw8mmuJbPtR9F+aVV5g93YDu0pM1tn5UY4hqN08
PCKwVlPZJcbkNu/APzo4FH8ms2Ix87JzXiZvKK+LQLlw+AvixB3pKYy92fCSpr5S
KeC/yRkGLqxpGRtHNsROKAGBpqZzktt4g3kc6ai2df1w1UjpBbCEeSSVSA8ImUWf
dsjY9STFSGqzIj+MbDP4WqpfBfUEgIhci/NKPIjfhIexnik20l7MxEPQAhhxpziL
6RfMGSVD53wmHsEBJ4HYTvOHLhP7Y6HRP3gpsY/+XNDBnv0y/ixtOGiSULwfdR6Y
7HzZhHd5O9a86V92oTcnQS0wdvVfjeoOv0FTEjR/Xw4Jh2WGzOMCSaT3U7Jlf5J6
avgvfdIV77/7HxUy8huMzbC8nOu9YbyVO9Xaeoc4ZvbSenog08E3j3u5SCbHFdY0
JW6hN0RSx5I7Q8+hdym71PWt4W/q5r4tjeEKht7Uytpq3KIc7/aiCMlvkIL/33jQ
vHtY+wxULiOIYhaiESwMBCYKjc2lkphHnqIVWN7M74DOsSU1T5P3ToXZB/fuTE2M
thCnai3uByyVYiC5pbx/sxFFevtYIWNl3yIkxT9W6hIxgCRNwWKootK5MhJXbFdV
qIbjU9qXln90V3aH0bWGSmsBRu/4HwSDURvGAvCirTW/ouOUZf7giJOwcRmxHWY8
49IG3rVInrp/XIf2YZ5vhkdz/yhGWeh+xHP2XHseuZ7gi2YEkoAgCRYxOFhd3TN3
0Ot4bt5NVTfgiRUTM17seAED6361tQbfmF7OpJN9iuurycwpoDYMBtfhVDc/ebNQ
mMsVNkVQ1AwVL7FPhL5W+FSmHps2Zq/+Qc3bCaYdACGbq/BogVMNc0ZhJKo0958U
mScxngW0/RVVLWQDr1Ks7lzHC1bcfeTTXV3ZQsX/RnLSGFXETlEIy9aiQYDUsPPj
wzvTB1XnQFgCWYUG11817umYjYF7APA2J6lw/gyeCAG5buT5nDDF9gNuHux27AcU
faoeLJIXQk9tEPirzqP7Z33DgoHyr88n6HzRmgaraTObJVq5Lu+5rsqoBtTv8t+K
+gTKGJIqcMFtkcy/tTg0qQc13s/GLrQOkXM3OAFTm2S8CPfr7aB1Ux6mmEcAjXRp
ZY/EgoJUZR/Hz9JxFwrLm4P7kJig/e5SNgVdK8xwvvGZIBvGyhkFdaG0886b5v96
Mtl/VvPAnE/Ulkb1bGhEUtvbd05+Qc4WwO/L7nVsNYrrG1XYV/OWUxu87PskRiJG
Jr2fYzwmpK2hhsM9x6rg0ErLY65xwJ2S4fxJd8cFGxQU+X/n6VTesifq1+QrmZJc
6FR4qr+jcvYC/+Eu5xmZ4e7/uSYcd1IYp5GgzqKETZqUcxpMwSOvHByuwDk5sjyd
+onhj3ztJ3NnJggq9nYWm4SkdXOzEsk9f8af+xNH3XSqjZi1Dp/ZJVrzXl+fKfkc
ggH506jFDn1HvFu9+DaU1XhPxhAvaRAUUlxCBTsIUikeGZ1xkWqb/kKw9/eAYYcs
1vIdMyCd3UX7IZKgj34gHJNRyQ/xLC7FXAcsNxjMjP3TOcnV5hiCbU/PuNuQGiqx
oom+1/OtDIu0vqb5M03XugAVcs6RU0lkFwM7Ln5YVd/hDubpG2OTudwJK5s2AcUx
C6QYhUzjYAjEdZ9tLQ1ngwBVvKdJYOTbbmPjXy/o16LTzWiAwz+igj16ueUlB/jn
SJYgcJXHvbNpJqrCXb2zgUQ8Kv/Ol1VPhVwfzO6UIn7pWba6/EAeFVCZRKVNmAdt
kHlW+Xy3oq2ODcYnU7slCeNJ3ZcBxM23sXe4vXjfF5ZHNgfe7RkYsPxBp5qWBdKv
WX6r1Bi+GjpA5/GX2NLJ4DwLFdmD/2Jmsoha04IHrGPkNjUg01ksWi85JCM/cG2j
PganFkqs9LHTYwWlyIx2u1fQQDbwOEiZccSzf2yIsomcO2IBkolICCuDcTwMG1E8
1450cn+tpAm7VTDyfCDMKWt0yNi+S+cXhZm5mImVzw+lH2Dv81YXM7S+RbpiMM3K
2kDf5m6lPRUFQpUkA0Q4t+K00DWYHV/UfC+qunuYPVhOuWTl6XekTC8gne0g/9gC
M2Tvm5Tzi1gwPWiYld/1uy5oFEQYkL8+HDyTeRIVY9/Ntj4erEhlYwS8ANHxUm2Q
xib2s8s/43tvx1DXBM8zLZumeVtRidgKLZQZzm0KK6UcizTz+Q4+b97bJF3Ornd8
LGiTD6cFKltjvP1VlIpywrB4m718LmCErzZObCL/v3V9CK7+dLYPwsR+VMj9Zz6G
EVdVg5MIRTFBVH5HzSJs9+l6AAY/LtUF0AJZ1cVsbBhrokf8RnnL08o9Us72sqAG
5uIVK9p8cpMhcXX/T0oKVnvHu6I3yo8L/QIkiSpSBwsVNyXTfSKSaw513yOdHRhF
TUPmk+DQ+N3IZURFlDoT2vWYOVB/muwpzw7TsCzKK86rgIw7hcVipuSjhrhrfxC9
pbvqbbW0uROoT1jaQbuTTGXv3CB0o2kW/Z2lUnF+mtKIKkxX8B7lhDlQG462y+hu
nBemepSPF1Pkmb42ovnx/KDMfYsayXBKa8mfZvd++/FNDzNbLRbRw4Sop4AWVSHi
WE+CR10ZZ5ZMckP4WDclSSTeqnyyZTbm2QUCuxxikNEQAr/B05olHWia7eZgfHdU
oZhVfz/u4tnwHTZ3Z2NOAH4+tAfgCxlCIh8ZMWw9fjFdzobmlROTa+dASQxGbU98
QcB7RLUT5FNPw52lwhqSQtqGogYIFXzlMzGw/1h56qVH9J7DBXOIbENisdWnvvf0
Z+kOfvJfaUspSlfT3wv++9pfr35Miy8bMaE1AYN/wjzXxTbEfJWyd7kMi/TkVWRX
b5YFi8TvtEtq4mp97KP206Prcewo1o+HRFcypfDnd0c/y+eHa1g5qZNy1sHDFMMG
qaATqYrAck5fawHfw4af4KsA8mc9rM0Olzlf/K6Awq5IVxe6lollBO4fhMdCtMkD
hjIM3dDHFzBemqq6pkpP6/vl1f/gDi/v6eJ9MP5ilrU2Z9G5KQqVVi4LfK4TapEh
pkry0TAPicDeVVe+tWrpfj+1yFCqXOeYgk4qbWfLQIw8DbPLJBdRoi/DF5omaOkQ
SwRZDEfpdK8PAK53e4YT26jRIZfctJ3LFMGSnaDs1AVr5d0rAQe8DnZx3R1ItBKu
ZhREoXPpxDcD/pgkXScS2uJTdLlStxNMRqjixYM2Gf+lVoCK6e8KhUcrblNVdenT
ZYxBzo35dbSjURnkSU+iMHEKgcDHBlgyUAIyEmuWtXS1RGB1SGerob7W++XTvWeL
+Nzi9eC0hhKn3AUyi8PqV21OBAnep1DR1R+0ikXAIaSw3WuKohnxYivJGz6Bh5p0
QFtd+UwCV6eenbl0o55dcOEI4W9q9SPnZ0vaBI5lb1+zwXu7/lJjhfa27lNKf9T6
FDTZEnUbjAaZXIQiQPA46ntRtGAc2/QD1Y3dZmompj9vZMDiaZ4Voeet0Jn317DH
kpi+9P6Bu3ODUZwtobipyjoG/JJhw4T3SmRh/Z/t3xi6geGq0FYbcWiYGLzCITF8
K3wDfpYGOPbuUSaKykzGnsLhK2r7Htu5iW/lxj5KhhqyOjwOW5HSP7YBOzjQSJu3
AmMBtGJEn/3JhA8q/jsOyKo+N7G6WzJsoa1cE/T6PLTFPz7jmJwCT6oIeFKIC6dY
UDQ+OT+dJ6/BsJjGhqjwz9kR/bGFFoyKi2C1igvqHXAgPzELwTVGcF+h6Bd/s0Vp
Yc4RAF4/sFwYoUoo+4dMpBz2eh/UxElCGAGoU24KZCKLVbVEPee+s2JufKY9KW8b
d9HxR4eGjxNinkdcIr2Vp1OlgSMfW27wKb1MamJ4lktDtML6PoZPe2ojaMlEgelX
87k31KBfuoROspBnGYQRNWTSdFeAmrIbZkHRXFNu0mG+i6GDYPJquRgo4WLSgKe+
aumiV+bDp/H9On7Fjo7qBcnbgl3EE/BcO1Dd2yCg85cUPfP4IlIFuuL5VZ8MTsRH
vZW/dlUcf47klxdL9wpXzxhbhuADrJYYthrKvsXdbfEHYOQ2kiSBZlBLtlTxeAfp
1nYMqFHnElOYZytIp2UODzxIEesK0/jx5SWJ5cn1bn4/IRBQ7CU7lnWwvfOzQsUT
CmP1aorRdqlxajvmmLJFeJ7QWHY40e9kREX6LDH/ELXoOIhHJ+Na0KAO3bnquK+L
CHdbEIlnvKqx0ETe6MwE6UybHS49kUA2Nu0t/C9SI0Smg2RET/vYcpof9TzlGG1U
puwX4IhNQuy1mNxid4COEUyfhpC8A5iCZTv0QYZpnSfXufmud4mfIaHa3yeKd+IE
d8KF9dsqtZtNkURtimhDW4BlolkG++N1S6GdbmfyDaWErskOgrPV4XDof8JgByRw
36kXhcnxaF0LcCMsLl6xzEYXnuhQ0FUG8HIFMB0kNhs5AHWNytuCpveBM8RXr4b/
AlDMtzzEALkTGG58J6qdpV4isQX7I0IQA6oOBUdBHPTSZ1T6lBI5hF51VLh19hTq
3jwEjMbY991YzuNYb86ytCfo/iCvfVtkYx/wnS1A0CmqguNXfcxXsipR8IfNDbU/
PtkI4soSr/SaSJKIT8qD6byUbBnHKeVpqsov/dCa78JiIulASjB760pp/WejdJPt
pwIDvCH0j9aHbr72FzROW7hHuZn8M1ojM6KSdNy//JXyJeColZB+3cDcIHybnaRY
6TG8NaQl3F2NbbXPtfYnIgPwsh9+2zvgflS9bTaWq9VQjoVJuyVPsePXMmrIbL+Y
I0pvIzGy8CaBkfQV3T6xR6S3QE3X+PMpLOU40eMrPQxoGsDuBQGh7F0h9m2ja1vg
V2t4HlX+dB8Zs0N5qci27Nz0q6EuKUrOu2LjPMCUbmmkgqbPohKj5u+INCim4zGj
OYzfOjTyQKI0T72d5PiZDSRpc5qyFRTTk7vdD54ZlPrlHPmsSvy857B4SQraYZe0
Y0z06XF2upUMJueUaB/bO1SKlJGq5NvcwRmoNGDNA6XgG5MkzhJsVu1eyy+dyHJd
NDrlx8ghm9fLjG6qCqDUIBW95OH3b4XmLLCvdQhJ7kIorvuLyRdaLXXBJNGg8hlV
wnIL6pKZoi5SYa8q8jn58+bzx3aNhslfxML5cBTXIbY52JZ49OVIdPlJR3Xw2BOK
UV9/H2VLOJP6DiYLnfyjQ62tAgPLGstHJCZHxNTD+W2ZKyf48iUqHQo5Z79aBP8Y
ibgDZfg20xZt89Jxsn22sXuIJJiwr6DoJr4MYfUQnvsHUmz+Ck7pomsP6tgAFvuH
Ah4BQDTW3U/tGvHPFSdaplrfjvgRqioSMYgCESpoGY5LBNBuY1XxFWAdzsBglNRF
oMAtuThr0dBtAfMgZd31TfzXhS2y5YZN7D+sB9KcgV6ncH/ZCGdCz8WdBE+EgUmt
G7QeFByPeEdsDSJzFBc22kE8yr6DLvUhRm0vsVlIekOHGnalZraI1YnoEgIRgugj
MoJdB2bXi/DmdI3+EkVDnehbY6xDSKDI0k8XrS3AXIDlqGRGQuvcJDolZRHzIymN
ZcxvYDadMOmB/B0lCxQpUJ+bD2K2+t1+J2RfDi/NGB0XGjEoiSeirBL9Me69LA6l
MFRw13Jlwmk5kPpZLc943+/pvor3nrSSkzwzhgV4vJaI2mq0ZS0SNdx7kuLxhwt6
hPftbmM0INTJcc8LiW3IA70sMQqEmlghAutA5hBqjaOYR8knGBKs++hRUF+cuhuF
6ud1+GCK7LOPXhM18aMLpo68p6T8NPCyjSHI08BtZ3WIK7IFgf6bDnhtpMtpUo43
Wg29JfILcS6Iqo8y2vTUZVLKXY+F9QRIqZeK2Z7F3F+nBP6iUyPVtzo2AWVfHFyY
Chi8b9S0wwQgWp3AnZkKBTbye2wW12XJMaNJIoLK/a+5js/ihxSKw96yHdCNYEHl
UUTwHB8RP9uO7s3oZpQ7pzLhcUDYnx2yz2g4k0JvP5cpkI9toJfEq4ZYDNUIncDG
M2svRB7pIjbBpcvwAnDhvmKtJO3ihDxMsREiJtqL2BzaMCQ4gNYGT0yGY6rjbmlF
4wb/+LTNaSIhk5AC7rT7aBvUyet0GfKrMb3HzXODELCVnP1War4b0YApQr3a/W/u
YayofXz1CjPQHbShlUXVas9pCIvPR3wCVjtfcOOSREt85Eu4IwmNjEHQuIR6HCUR
u9StRojKh+LDp/6lcGpuYSIU3Q0npVdoQiB1E/V5TyslYlOsPn4/+AAPLhgQLRON
UEdCNidITYOeusnRjFXZ2zIAiwqptUf1v3HVRsX4rgsXVDC6yKbs9v9YKGMgtSKN
pXECjuqTxRJXFBnWgwV96x7hYrKiw0Hs6CAN9zF8pyYsXQ44FC+VOKsimfBGke9C
pFWOK+kxsLxdNau+CQKMDCbUJ5zQ4TI0NdzY3y9IbDmWiGOR8oVOwCrFqBYuqGNT
03NnIgtHsj/EoIo1wQA9iW5zTxhfj8VHuv2X4jnMCOJTaFi6FG94h45GZaGjq44T
1D2107OUFcRFB8I2UjMbuX5Xa7fNlswiOtCdlAI5A0twjMshWijmwZRwYUidWinV
/VeJbFGQqCN0X9l261Q+9Jhaj8lmfhVo+/aCAZWYK7VLuv3p26rDh6rafKVtjop8
XAQ2Ya2RKhjo7IxTAQS4j35EP4Wyf2rYtERWzVBtmfAAW193sIoWt4HbyC8EKqGT
b8+ZWXSZZipoK7W6nePf2s0sVCN/hdSijxWGahubRp4717pik9pvu/Dm98LAfrZD
KdtP09PM5Cf2CcqntHi0+PUvw0932tVKhGN8CfwNtg1tph5jpeZsbDszBuzHJnQg
pbp7248oXQ92Y1F/ylgUZBGokw6W774lQInOdyo5NVXj715xUUoLhYD2pEEpkMlr
Xt/EYIO9Swrl/n2rdNnmaTyynZZE8BkgZnqbmu2945AWB8v3HL+43ZyjiZGuvXdZ
OzaOMYvoUPMksQXNYjvp8fCwgMnQCBZwZT6hxu1GWev88QrsLY0j9obnyIduArGS
/NJPrBo6jIyNaWLWk7c5wmKUGZofd1ua2OfOrFjSMU3lJagj6fDgjMSK9M8zE9hT
VOOa0MjyazWAPKOwVgwxlU4wKwGfkUyyvWTo6Lrmqo6MGb0jClnywHX+u/5/spvk
DIZVuz/raZHVr4nSmzEupPI9dvpnVy4o9cM4/fvD60UzKcBnxur0IaIY+ZO4Txs2
gwrGPKU70C7ZbStZ8xeY6f4oM596BWDPDYqKKtkEi1Qv+Grkf3P8NrKvL4rDuF/k
oV8bLr7ysDgwhJx/DjMdh4IxGoLqawjW9QHEKKfOUO3GopbxCf6IOtlih7d7vnpI
BqgMuOzlWYiUcLKNpKSjV6UFTVV1M67ubsiJJ2uDyLaXW100LqZI19UWpeesUP5B
FnwH3uAeT8jUDGqgzk0wXus0XM1tDpNnbBLDO1oSTBr7oaGkPCmDYTTdLdkE1wV5
xtsD5eBtUNbXsqlgVMzwxi69NHoAYKatHH44/NsaXgCVa2SNHtCGpfTlwo58FQRG
0yHV7xaHi8We0OUkiyC7wUSCDsmbX5XGXiR3vtZuJvK7IjKc8oLwscje4oM56Quo
0lnUExfCWYW7S6pI5E/2yek529tGchTFggcuPsfdgmU4t/l/LvOfFpklDfRdmpLl
FL46p1LYe8KHBeb9YUt2EFWc83PTp/LWbHYXKGa/0rSM4YGNOXDywuG8I6wHKfN8
sxXjc8sWlO6CvIJa0HYKayX5UmK4PgU/Ccf3kllAm/l8fgDxWACSYVucwlxyw6gG
MOfNIWCpZV3pViGh658umyiIpqXf/F8FB539c2vXoA6jrS/01/yVCjcRMBj2VRfC
ATvr8P/5DX3u4At7zI/T5FCekrSChsBivZPW41idzGBeOtnozSkXNIwzFcnfnP+u
qsY5949Wna/LXratxV8eQWJguVo8dwtinWFKa+TOg28DlETCg/D7GXnt1OUQC3jB
DwWShwJrQOXONIIfuxvFiDaeL9pXcFwvocaGeCymIXJm/8Oy3YJEGFxcJrTEoFrF
WlFzFpqR95B2fRnGnwZ9TT0P4TVailWqSfp7AdcZx0HcrJczzTYm6C/yuU8ob4K0
bRY0rHOHl0ROa1zlKjgSs7Sa+zZ6wYtok5gsTURpfW58Ws14hhCUevljIMzdYkgR
Ea3jMRL/FnekpJN1EMzqB8bEGgmQh5agYrg1XUM0+lYNw1bKdZSI5z2JlFSBF3kv
IJMVqfO7xcKFdpnmoaqjkXkQWe/xKQPlCD/+6zS46pV5wSIPIMoW16o0JasklSzS
WAnarJwRVyiMWPb3mNtmlgwgVK2MOLE2FTIo79Ho4GoNHZ6lJWpUdVoPxNB3tqkR
/FLSOn6ToA84s+wQF9aXu5HSZkxKTFzgQs6ON4oplRxOlj4+FyAH/YuSV6ze7QeR
cHK4xYdVROdmVv9uRxwTgiFxxxha5SPh2ch10djc0cIPDpUaOA9p8n2xn6kyZql3
jvezxTzkIbKsfBSTJVfocdj0fhqpvoQF3toAPm9jkZsclcHM+20M46V2s1cap5Cb
rRB2KlDXO40rhJIygPGQH8axppIFbc+gu/YAM236W82D1Yp8f8fCRYc/u56BSDd/
pFka3GOzgCmWpu0PFdW6dGOkOyfFaJBfJtbJtCP8yiRFQWuSHA63Cizmy7YCl1OA
zMWkwjuIOmNqPxkrYXR8vCAPhNu4Ob+JLO0QmTxfgkPljdK7FolB9tEFcNPZSK9u
/CZ5jGkRQsRsrs0Z0zTEe+xOzauuQtympGKSyLk4Q4zBZ+fFtItHyPXEsiyyUIq7
n3iOWDJeG8Gd8asbY7kjnh7R6pCgdU2NXfjHf2P4LqIOX1e6nSjkYW1WqQgOm7/W
g8v+WCb9hin8qe0+BzzumFzLq8FX+iXxIYgDhEzvXduIvldxV9RA2sJsffzAsSbz
p+yo4w8KVnCe6RTZpUnAymhfNOlcQmbe3DcCoawlm4+N2CxXRW7p8lhoVGdAKacu
wX5PftoDjwXMT4uJSqhpc03lUnUNG6GVrkfsSEg9LDOnDmmgHL7r2Wc5G5mUStK+
7n/4PiO90N1mgPCGzxGxOzTF5v1rdWRGKmLpezd3tkpYem0lbZujoecaMX1FDXzL
pfjN95N9t7F4CIZIGsTewNGrPrAkn9CR1uczcYghXBN1oksP6oP0Rcp+v5y41JrJ
OEw/FxW0S4yXJZB1GiXZLAIveu8a5dOYYohIXCa5s5ovK1aU3KIaKDdX4PR8czHx
OfBrE8nXcp9vicNQ0vG49N/Fib5ZzMbAgkvg4/TXEcHJ8zdJzs7Bdm7ezNVuqT6m
YHMQ5t3j8QxdVGL7SIvxypSbEewqZ3hC0rCi/B6gDnhxeVEhcs7Dt23KsjJ4hriV
iEgcBks9HG2BBKBxPMKIspCWRP906gQVn03y6liHE19K8/cno9lUoQQUfiho/+nY
n4VBP8buYznOITS+QODY2AJqpV133L82V0NbVzdUh3GV13tTVFfV/brcJCtDetht
LuOG2ky0H6OCo/4YMayfa+a+CzP92pB0mbYj+5Fw7szaM7yz2Wud/dVb6g0oKtxS
m1fTSb6im0A8PkI0PYzBsVBna3abfgnZhWFEm8tzpaNYNCXO9EJuk6uv1DBBArWj
U9FIZQ7RU3dniKixXP/zIk/hCpSdyMYYJ/WqDRYrJy/obc9MgBwH+xv+M3KB6OxN
/KRavy9pNv3E6/xhQBpyPPA5Gush189YjedBDYVpRnQ7lzFT+3NsS7Aq1i4PnaSu
NMN9SwRmGRUMZDN2XCEmwWQX0PEaoRaGn9h19BUOwX8H6wXU5PmToIfpkR668hPS
Q7RmG/a0NFwzZkHduXu8ZqDX3Pv0dNUNqlHqf/jJeaD/nBGPhS2C0AF2O5r85olD
tD71RH01kgzBfiRX9p0xGc1QOxkQjxOb7EwwCAP4avKzNjSAH8iC8ZOQSbRcqrpy
PHT5+5MCPQwDGgUtJtYmaT6+584wghiYrRjGmqg+5ksEyKjMGfincnu8nOtOOTfn
29Vw/sZ8YLS9oYCFcgtjVvFftBbQJlRvaAU26vno2euwajteAUUuUkkhD+I9hQaL
6DDqfwd/HNXFv0xYnAdY+dSRLDa2TzTrpOUrX7WzuN61TCrZEXjs11GcUQS1Wowu
UN5kHAuUVNNlKcn6TiWUr2AWLqJqp68jT5um3CAG0Dl8ihql+bX7SznMGyflBmMn
ZDnCDscvnkL568JzW9BT5HEZMc7nWVdZaGdj0Y1zBDo56pocU7FIUlpzzYDMXwds
rbP3Eae35WQ+bji0kQBZJNcjilpqkyAOVfrbrMh2/vfIA5sCwwG7+q1MOqzDiTsT
2G64heqkMNkAYTSxgp8k764InUHEmkTaKbuO0PGtjEw61pIRuEnoNX+h7sWEwU44
kVcTIC56xENo6GpwHw255dpJzRdtLO9c5jq78/dX5QRfXej0xnGosFcLQs9v/rsW
XEiyeNNUHfEl3uwAJEQhJO8ehH3oAf61ZPPpMNdnCYldBZH/ywiP20x84jJz8oxf
8dnaX8GcqWthhes4kCWIzdcgBwJuYfaXj1B+1cPztVezv6oPt90nq+FRH7sdd8jJ
2APIG8M+Icaok2aR+xcvmpbX6U2QJTvAGxbalq11U5+gm+5b2YbRyjEHTJY++Jny
cN8ddjVJO0+h0KdvcMM8lju9OV67O/JuPb2EqSt60LJC+U5V4v6CxrFvDh8/Ka+t
AFOF6QdC6tKBNvykoi8fgCTt4jss9YjAFS6PQsbIlJPD0XT24i64OpGV0NEMV1Qi
sUXyDqdAV4DAWGDabD+ytAbAt9lSlXiv+grajPA+lvTE1UiVGt76loAf2YLR0Rjm
YdqSATGSgt/C4FLRcNNmrxIH9UDxnFtOz2Yqs30gUdYJI9a99qaCBaFGc1gGH7Ha
BIPvjKNbH4Y0XRzAgjOQlEzPgNCDe9OMn3LEFuDBP8WTt7IoivorPXl2F8gJcaFp
p91zb/NMfd5S4qpf/I/A/MOitSB+Q2VAoLD+duVef1zwIhMxypPlm3UX24GxTlHZ
FlJEFdV0WDONRENPD/ngCx195BgXzMvFeCzNUghtBbZ5GFmKQe31p2fwQf6WNSfp
X9rCl97Ftq8VhxSHSgnngmFq8Wn6XZROKtbLPlFr70RvIlLkLvjuD+9Y4rfPJQIc
1spE/XyhejfgGq1JEOW7jGgn213+1dJKQuL/TV2id2FysO7cpn99w0BTXEe2wy5F
CBKgSXBKRSh5nwgqGhC9tDrNhHVWkguCqYV/WPAz08Xhkz09TLYkeWrDmEnLcEhE
tLzBPPT50oQMniTRYbwJiu7ivbGSYcVFyJZetQmkLy4YMFybtLwEELXFSdddZC5C
1isqBvPRr7LWoaQcvgW74p5mjAH7xfQ8CJJoYt3gSEd6LrJ9tMCN8Vb6bBE8Yd3W
I3gMeQxJhUsVV6shWnLZFRe2Y8UuowDAqpbPUHISQXrt/OqT3eXU9R88d9JkJWLz
kmKClr/sJcr5P9Jst8VVATkoL1Yazode8JiGY+GRKNBhH4yE5h2Qx8Ci673lQcZV
h2hegXLAGRZ0TWAcqCv+GWraAKCegwicYmRuNq/ah0OsuEnyppwd9P3GlAaTBmwF
bYUjo5atunBZUHRWJl0q4gc/r+sT7irFoeqmN6WFv1bYAUYVNDZ1jC4c5hBP66wL
tojJnV8FRVcJObl5DLh9dJA4G70uNq8QaVwjKQ7p2QCLmaOb8qiTkEkBeUKZXSST
nip1vtb/dct+L7MNmQchAK9Xvl5Ci5U9TMFSupCNkGtvCS2dJxKXooX6x76sYVrz
90eBGttD4UiaGHxE/R8KbZPn4vf1HRtfEEOmeTtthyWdoztCTYdkjDMBED8YRus5
O2w4eoBCgnOpBQtENy1zbRuMWFeZha//ORrBGWtHihtxawG/Wv40eN71/BS68pPQ
NLNg5ZbXpdfpg7AzkPVYJPPgzJBpydvIako8WiCUC8qVkan48IVTDM1uZgjfu4vX
2RpoalrVcZP8KgTzi7h4k0hXGACtyUgAl6QkOObaxVjvkDX0tvs3rFCN93U807+W
VDlI2xCfohUGgqNFyEaDeGzTM05s/lnRn/EAqRKGLE+/r4G5cW2N5z7fBEZfDTpn
vOfTn1jNH8glG+VbSaomfRFJy2GmONZYrAq15jjZp1wPOb2cBRxslP3efc9WgKH+
tNU3rqLYhMM0xtGJt0bJESki5VdpjqFI3ZczO0IWLFApuawGhRiJ7nc/FnbWFzNV
mT118alUz63UPJvNGAJIYUmF6Cty6tDy6aqogy3pMHM66ZRfDwZ7g2OLpuoWyIIs
p16LOi7zPXbkTJxhBCjoA1nc5U/xUKX0x9F49t6UkMU34KaQHFS6KlpTSzINiM2o
ZYJa/Yk2SV8howPAmgSOU+X0t5LOEIi6ZuJ1NeuMqy3A+ZJMWJ6qiESReYydUr2W
2viMy6JnvILCfOjne4it6NYttYlyalXbX8OwRO/A9LMc+JGb2AZmkhSvjDu7c3TG
a52BZSM6/cCmE7C79Hsldtxe5X1xwp4FEj/cPwUBlRRIECD5HohVZdtREfOqn2/8
B5W/ljZ1mffr1PtKloHQbwqtYGwrub8wNDgnoHvGMpsMBt2wWBVifrE8q82kEcQf
jnMiqq3BcDI7Bv4jMAqjGrH1dInHq1PnhRun2gy8/qIifMA9MOFOzhOD9UwzTCkK
32/71ODYB+IGxAmnzAIVL/RnH4gqP1krY5wSwjDtisoYY1lnX5rOxF9AlL6HRVmK
cUAkORXf2L4beGZb2uV/XcliHgCPgV7zuklQdmatDlSwbIPRMAd0EF8apL01D8LV
b2OCy+zN9H3XjCNc7NHUiyNLPHODH10xK8mA2KqalXxCuV3vNGRVupmU5vmWHEp3
ZQMRoWwU6CqVYDodZuBYFIw7J3NrPkXPEHzIs3d3e8q2rrQZsjwQUk/bssoG7WgI
+jiC42gI8zrs0z+bu0CroGVt9jymoOlxWBBgNO5U/+YaNPatlvZ5E6MeXhaKtwKL
EdJflZJ+3SB2uVb/4cqiM7gTEbdJ1WYP3Qxs6u21Wbvd4qr33HADGC9NL+oCYKW+
n5Zeyg+dP9Pd8dJNDaGpMFIkZkdJ2lNcNEB60qCnhfqnsYzuWdUVpabHtdMNchgn
7cSFhidAYvRo2G8cmmjHDliY91ASKvp0Gx0hjSkGWQnf6Xgoxs32F7Bg7JryTQPF
W649ABBga1JeoSxJOpKTYt6VLjjF9Fx5m4yw2UX3HWxMxk+qt9D12il1LI18oDfJ
BYm5wvbd/iEvMD+yfl69Z+i0x17q2ypl4Fw0p4PhE16oi8Z8YSEh8MH0sMNtWNje
QjQ0/Of0X9F2yqVsW67NiDgrMccl3WisDP1F8r/aqWOhSr1yWdvjKXRS76/hTBIf
+8vjVKKOhjvyiUeeicD+ZixUh+MdkQYbMuIXGHUmH0HNKzYdfkXjhWM5g/g3ZpPa
eVhcgEAqt+DsRvqPp+q6I72Nc7+ceG3y2+lWxpLvYl78NKhg63uLebS/iKd78Gx4
Kqpqd5QRbYHLBhEQTUK5sQj96GSPmlwKGHoa7L2Kf5uSoHUwzEg138BDogAgRiOE
NtKMTVdVxZh2Un7zB0qAlYVONGMLFQn3v+WzzeXsg0uZHtPzv+1dnTkuQ3XtfcKG
5nEOcJrwFC0LD7WVO/VNyBaY9ks7vmdLNnXByhlCtPiXQuMDL9rVtihv4eIFem+i
h4UxP3AJ0bzOAbhJ0wjYimEHNuwcX9Dd8Qq5NZ/wcwCU8oHgQom8gJ6IOxmRtbnU
RY7IGTjrQXAlMvF0p/VU7alCg5SBRshWDriCKacYc/LqLmm0w1tX5j5Q36OzN2UT
AFTeTnT+hVG0fSB9bFNsiifwQyodhFgGCFiQLCstS+lJGJx9qpPiQkmjGKUPYV6Z
uYd5nj64uSn5+YJi5w4hPH6kmXGC5L0Ml2A+V1oqvYND/NlOFmfRB+EB/G8NHFE/
mvc+yRlV/rlSfP9+nTzDKcJBIx+V8oKBwBbHEasbWWbsaoHn6FXeMKyo+yPxFxmn
ow8zl/ej+qzqeRShWI8yME69aFwS5ExtGPrZ60JmNLN4lyIbram8nBi1lWy+wvgV
x0fgduG2Sim9JwW+0THnRMFYuxo0udyrqugQqQxWgeWAEFgF9uiVu7Bxmdr+ipJW
OAN6+lU3caM4ZSAb4FoGY4luj3Ifwf+yWkd63vp00TqBPxoY301aTSRdrxRO4N3b
Mc4b0ydMUbQPkP7EZdmqcOkqC9C1VDDA94bf9SZJizDrUm54tl8u+CwUwky7xvT1
L2OlDQvpUSWHIAsjuAOrB1mHqCWf32KVNU/rGzd0omK7px12x3DGUv84cEQ7fU+e
jLNrOmVquSay82+bhdJC5pOYojKWn/deE9TJ5PK8LSDNOMG6E2PXbwS0osRxBDme
pW6ZPzh/TwHtRjK47kIxfDuDA8+ek0RVKolBxWWgwU2Hy0AHXN7f5XMSMHOA5+68
KBIEQMb+ggjg0VS6d6UkkwpOdl/ZjL/Mwq8VWkQ3kH2Y82h0RZtMBk4XvTmM9nkZ
/WU7DjZoSBLkl14M6PFnK+rjbXccbwgfWJF9tnzEbi5KUwVBpgP0QZq5fjy+3E4D
XL84taflrTU7FINbqdTbC4MmQ7FypQlLou3IYUqB8I723JkuSQUqzepxczr3TJ6n
QfhwluDJ+vGc5g3jDg3Z0XTt+dbpSPcu659pabrJYkDiRK3AbJhBzaHXeQDHKdMG
3K7cYejB9SdM4NtTK9AgmRM+iMbsNUg9f2yq7l5EPT4/a0/XJ+UE8ssieCmWuD5c
gAMueGNBD7gMh0TrDE62swsgcmcgSUDxJ/zHsBkETEtbZJGpHErrzMF5g/sMnYh9
LNn0qtWU2enAdRPuD7Af/kiBS8DgLCyA90qM6lJpF7mAfWUOufH8TGv16QO5fbtn
ieBw4ekiVZovOBxZ6o6f/py78FhD2AEcyD/f1GJskOLYklHVLrpruPZTpAXBKuHq
m0SJIg4+CWiKaDmuD7KBo98HmgynMuAt4jZxHJ88XdstSvyDn26npqyt6ee08CCc
sWobv74Rb4XK9kZRL4mFZCi7vPIcziNYEmoxxTsHo7o2sKla8xV8G+TWHH3WOpxz
Kioq7mXKqaExETwlZ59Vv6CfmQgWOX5tBNM82cM3jHKE3i6PX+Gfl5SzIXYkyruq
E8T60BoRLcV2vpEwG8KrylZ0EHPIGZAI6NKMtRcUxCnrxxvRsxMeIeeetaC6142c
QAtxwgmJMw+gm5CIphPeVyfLphVrg8t02je823zwU5kzGf5sEfnkC02l2UatvhNM
ebv+pAarqjIkFp+4wH8CRT5hg6pnipSKD1yAdnvKJtzyN+WA5gBGC+wZA0XuqA/j
17T+OAfIEkZFJgligmkiXvlCVGVY1/ZBtcWMD2TZ/875otlMtG6xHhBBoL9gYqMS
mlf2hJCd89qZxZqLWorvhyRmlQPgzNxPXG0tKjm3BsSOhSVEOJxNWTHrxvAiqbFs
Z5Cx2FnbSMKjiD2iQAwnYMDHrewadGmXGuM+7L9lqWmMBvWsLSqOd5hu0q8pl3e1
9m5qygkrkeOZfjHIgzlHfF6DhDDa9JcKSFeV9aWJh5az1UYMxSzTLnRpZUzGJWNX
R5m+2/qpL4sDMSxCvatUI7tFXNylQBU+p3X8ttTJG2VbMizFwHR8UbiPjLEGnqRL
CkJmta226OtJ2TI+4V2IueZBfVedPBGwJlC014nXBQpLzXBXOxQ1USLiimslmauc
eEL3/uWcKP+ukYy38XHbIS8cLttCuvwsTSytcDkkgQ5ih2Y+AZ3Nk4e74RTOrkjW
UBbNlPHPSxobTAJLRPmWnZs9H5P2CrBWnHbojfaK+IPMdYDUH2FwwBjNWJA3BFXb
llK+AtrF7EY2wawmkgauDG24w57zm3v6AvgUONo+O8mCSMhgOkO/DYZRcD0nRRPt
DKwpxjZmwh8IaarETHW74tUbpqJG9QbW1ZWaM2e+XObxl1lHS6QxgMO6QP6kYjOS
LsF42X63N9z0bDWH4ac3PAvWouA10//QOMtV+nWwv9s28/pKSyoCYN+S3e1rvFh6
qivDdY9PHbvb7/gW2cBAOCuwTbFFdFYPwRcRD+mwcBTYyHLsixzw4b3umB8LtsB+
/Rfhb/2kmw+IszR2omC1RSFSS/4IVyetRKR/l+TLFznfBSuVtw8q0c0iAUv8vVua
VP8Txef5VxSdTRqTtp1fQHgYFn5sZu5xCsq6YMnRj3Xse9OiY2LnChLqT+m1mF55
FG7QUFfx2kTHcqVjHLzHYj7WVc4/CGMqIk5Gy1OZIphss3jxJx+FrOEG1D9QBeVM
GELQqIbVwinDxaoWf7xE2n/H00+5Jhc/QqskMIasz0U3rLbMbY9Hw1dPSuZGZgec
pRMQIwOQ78X16A18O2KLuDJk+b5vr9PYqW/xjrU93Qwow3cx3QldE+3sBtEZvLAv
e9WygR8RY5mmrRJ7BGakNgPesbhAyk2jsYI8IJD0ZGnS/lqzufXY00FapQRfz5ki
1kDwUftkRChNWDSgJl1pJGm/JOk/SJBsCyNp744W9XEEHisjklesCrF5k4Sl4yDD
Fy9QFXj4Eyk4JMcWeQDdX34156tnZHIhKZwxSKTfis0nGtM/dyWD67HcmPNamqP/
EbxllEfTEtmNvYmtqxraOjOBVlXu45NyUbhBzVKaH2ODPUAQQipDd6AzJ8/T9QLu
Fnj+L668UAUzZ/ZTqCWXbWRPtGU3TO42XycBj0rI0z54k40Pp9pnptp0RGbYwIpC
zZEYjJDAQBcbND6r7PNAkas5v/r3/llWrzF1AOCuTayupHP5FYrZGhPFJrImA5PD
GDWhKV3VMc5Sat8QF7xlNwwIW1+XA8+mqsbz2HtW7RBPZ0sfuqPPslN5buuRiFFR
03cXQYIab5JD8LPqLolF1mNTWVp2J4f6oqVBTXgoFYyGnGZhsMqBu8762vXvyqCO
AloFyndwlO+6R0PwfkGRsirnA0j/kKnVf/Vc3w2pHO88OlDyCEwpvJYMf9PpBmL0
cHKCGDyAQppy0So8YjZIVEXzC0XHIDt3k4IbsmmmlmzvWJ3wo6JWuHySMorzy1Dv
zGUTWP+hUcIJUjqi8TlGRQzFnI54z8FTNxdeBNxWTVPONRnWP3+GFn225Mbj17Tg
vM0G/p8PX0h2vg5fomAPDhULGSsWpRJCTeeiH/HsHyp7dmBCdC0NEgv1lhu/WTGi
7WJruwf/Gg9o6xU2IQpOwaj2kHSL5m4i/8hi+flXG/BZr6Ta6S+ZmWN4eH28uvoM
pwruvnQyu2P8cRc/jugoZC78FFQoLBRHEXEhnYLFcmY2T7azS5ThsBnnxsOePF36
Rd3FDLCzSZMnaM+hBac5Z5aj9/Gc7bePKAk16bGqWyBOGP0JB0cQnvGciVAt6zIf
xQhN0YR5EcgrEfCMj+GSrJOo/8jH6H/vWo3cRBAcSV4whkIBJoPNGqofgqwVb0fz
pEsJVDjqh3xd9raNIKewBmx5edbD40VnLKY55BHdlFBFyREE68CksHkDOdHWf/o2
ZQezkpNI2V02fJi8UFjPKGZPtqV7nN3ixofSRHaIqxBZamIk402bVSCE+rZIjdlJ
Mb6WxKohSYHV7xYUAZCxSuNbCE8iZFknWUkEL4n7e1gSxCLbFWX6biE6RcnjmhE9
fG0T1/buT3Q5badOQfVpqoiJBT7rH4sad13uFvMYFRHmXY7fTZZktaIsBP0JBJB0
qL45bAjEvLWEs0WBka2YpZyQn5PhRhjmOHU8JZJa24TYNCJMfUIx02MQnfhERv5w
HNUUcKl8G/i67grb6/DcNeu53FAJHEtvFWSSge9GRE7hd9onGUROw0ulutdpSgLx
mL9b52vKNaCQtnNNV5frYllMPZcK0/MZSXQ5QqTF5qFhXDAqjOFm4AHoYGD3XxSs
NGeZfMOtOan1SByG9WqVIv/QB9mkJ1VvnGKR9lCa7CfM1DtBs0KVGFBf+8wcT8l4
KMdDEGejb/D384wAjNq/g10Qv7/SRlUBVyukfCTPDZVf+zQld7Xyndu5CKChyQa5
tsZh4zzOt+rxe21y5cCZHVi4un6kYNtJWIhBWyn2kqN4z86n/OuwxEdRHLbPVS06
1oQoJKiGM6e68bFB6ArNeiX0SC5mG3b4M0/u0o6fYbUzYP2AAXjm7sTibaooVsh9
pzQeskQg+4Q1BQoo6YW6q4xDixruWxwS4i80qT4h4coyw0RaBszPdAgvTGuM7Ik2
wWLUU7WyP4pXVdIiJhrQXCWvawcuLZ/zUPMSGOoTvh7r3ZAPZsodcnKPsAog6a7i
r4I/iwdLg8K+7AhW2pZoLT4Ve0a0zQgo/wBiccWptA02T2K0CCnzYFrkiEHXlFM7
foGK3G69sx084H6wpzNw5IRsnF3ebZMBVQd2P9xuVOkQ4sNCNxsNYRqWxyfF1Svq
PIIb+FRGf+ewpO1eg9waDNB4O2dDgKwgzcM5LUtyIC+Bqn5tAHQlJAlVnqCsBrB8
LsZZJa8cLx6CA/RnQ2JJxNAhBwZ2bQDa+3V6PfKV7mo9SI35VPYjtYJ6B2Aqyx+z
dZ1W8rI7ANF0A5cge0QSCrRqfOee7pVUdRD5E3bFgBWyGWRJA9DhM9CDtHJkfgHC
RrtcvTm4bNF7WkHxD5orv3DZkKg1ozfxqBFQ6Lz4OeXpuC3iPJEckDxiKKaIskRU
zoQDHdeRJpU4OEbA5kxfUsR3iBRzBnpQfhomS/x+AM8c8qnwv/2urGQN1K1qVTh4
xlY7DTQMlPWxsYMW/uhJ1MR8xr7Ys47C69Mj1lkrWqz2n03K2G5dd0Cevi1eB+iT
QFNa/8Ly6XDc3tIQCCO6OcatpFCDmidnx41yec92euifgI38WeOFnMAxwEUQmfIz
/vcZE9DWtGXYk5mw8eNaTAmd8zqUvpaMXU9+NyuWDUvRvOwos9YcvZhjemr4nKT7
QRiX9hg0Jgn57JBR4rVbVCo5Ts+0cXbijRNy8n/bpkSJKSzU96iYkl3TH1rCOZr5
nDERzZ3IaXY8O6TPxDuIxTLEPRs/oPnoLvCx5kBA3fZt5NgNwDbfKJJzJarrH3qM
3T4+pHRyFJZ0Y7O/xYc3HZMu1/APo+hHn9B7s1dayNqFM8qHTN8FTapYRM6WpQkX
IK+ROHPWNJf2mKNLTqgafM0JRGxzBXvdFRJaCchIbWLvDKg2sjVZt3kJEB6O5zaG
eTtSk5qun5BBZylSOjEZvyxWbWg/T9phlyi+6fiCQDvUObdwFaRPbRGwWQ380VhC
mraJL63bp9D0MGsGe8dBupS+Y7PRY9e7ryl64+MCqNMj5JRMiBDPTlflsDTh24HA
C/Fw2SonRhSsvHTa7nLzWm59bUQX3h0QmFWuvHmkgOEgS8xt6sTDE/pryZ9vBokp
VOcE4D5YfyJX6nfS7RkFAOi3GbTJjkxELO9fACooQdL2tXPVsp9eTykt45UaumyN
asOu1ufcEHa90SN7AhdqzhY1lQL5dkacjXtzdgsZ6vxzLjkkD0b7grS59Ym5iZ58
j3bFxrUhD2CPjB/a5vuucLsrrXh2HhQ1jPBM2wvE99P7+y5DxEnJlLhmMh3VcTS/
3KlpRMRApGM1X97FrW2q/n45dM3ksbMo5LcCVX9sfjXAXel8D67jaJd5pZv9d4Na
w65rt6MFWn9lnjm4Gfn1uDTtVRrJ9BX371JA9iMJtrZw2KtfH9aOQ8VM3y2/ISZa
gxpy9MnDQegxz5M42nSIoxeYRSTJw2FD0UFuazMJPTV10FzxjwQcG94WSXdiaSTa
Fn2DzuNuzYwuZZS6OIr3Qz0p20Ej7q/rbEjb1FipsX23GUaOlNfBSj10Fh30prNQ
DRwNnQ+kp+zEY07PuwbSVT/s0cKUrAt3eAxpxApchWkMzPaabsYn5vM90W2j/NOx
Wf339zL4QiNakJvihstN8Ieew9QJbuOABPmbuRpGDJsCZBdRXlmVM+gDUQ00v6b0
vZN2738/LiqCY6nyRwiI4YMWpt0gr8wxaMY4rSVek7z4cZGA7uL+/lMIXtqyd6Zm
LKO9if/9pJNgQ9sRb7S1XOV8RpUNAtg35k4S71jK/H8SfhgHvrX9btVcuf7g3GMK
IYbZ+GEZTwwCXdihVe4Mr8VHTx+t8uhEhorELV+CmCLrTvwYJS1uKvivSjwHpKw0
2Z/gsoeVjfWKnLZQql67xxZyCb5+moVFY2azgT9FDYJflrX/1CKAHcGJh/YGP4CA
Wql+BLFZ05wlLH5SJaWJp0Yc+DjiDloUSZn5N0iWw8BGA/sXZiiJ0jvurXLdlkXz
Dzy4VaxOHl3YuVaBu97DRqKrxW4ponHgHnstvjGEloR0xn+PBAF5H9sgR8DuH5iG
61hN+fP4SQgy2ReDeeanu7ewAcmWWoyegtJQcycjO719aqxwC+o6neiMMe8u757C
incrQg4OUXtDv/GO2tq0cPAdvPGQOiUVbMHI8B8WKSHxpQGB4ZuBgwEmRcMHCNIw
Ir5P4v3nuOiP1Lef9iyiHOqhGFfX4rs6RfmvurR2nYSq5Ou1p4MFtZtxn9oL/x9A
a2a3VGUhS+L8YZ936tpaPGahnzCHyRJOgt9asdIDEERaWIXgctvRVla9ajDkCdDR
Cqs9jNS4Aefu9RsY/PYStqgFdJxLnmNLsdowUg3aLFgKELLYhBTUUaLXv3SVkX+Z
tFT9W6Dg6g5HmOxBdXjJYukiZBMS8lQ32+9439Ha6AoJWciu5b2hDpiQ1g8PBnOk
Qf5aOhLMm7/QZt9Ago9Qf5cQfg3F41YcxT41VJR3TI/ZDFIIjHucrCa27qk4cDnT
8sjfYTt5iggaJ3StyTd0P4JCx4IgSJOvfrzgtR1aP9JxzvED/p3US1Gn2JSHcgim
KgBrsnMGtj//Z8lHfgOR6rHobzHGSxxONETIv7tUjHOaYNJdqdtVB77dh1JXXR+a
hmbUWrpmJBlcJ6x0cwNmnT2qKMMuFtdBVB3SYG42HR7S+Pv/BpcoCG0ggmRiCmJ2
lsYBGbLSEeW7AxX8RKxYE60XK/Qzk38R6+NYZHNMX2GRKPB4xVbD15jKnAUewu8u
cYo0NJi7nHOYcdrsWu7UcMDoioHuHUmELfixdp/mWBm5jpmJCvy9T9yIWOLnjCug
17IUrv0b/f8LAzHS3VswLF/yXIX0oGz12t+/a8c3ck1eIqA5EqxjIdSGTsm5Q3Bm
n6AhkmJBCNXwycEOc0sBgKYcYTdahip67Ju6fK78ChIAO5KOq7ZbPoAEjjIj2cS8
jrLLRqi2cdMlr0HWpenh71rr2VL/ghPVPSengVZ/ssx1CpU373k78nWFRs/gjI4a
yU07w36ZWcSCPXC9hfwyktxbp61Xzc3qyBKXXjhcKRLMUrrUKDguOWb123t4/+cq
cFlxL1bXUljhl0Ep/qF3MM1I31D+jkJt3yAoczNkFPXRSpPcosvfgk0zOpvAHwj5
naw61NARbV2x5Fe+FqxWPTdAt0c2nfAwQ4xpkoUe8mjbheydXx+Q0ncv+zEXkeeq
STqDyTKILb6VPLDOL4lfpHMehsyj8T0fV2jDHbUSg+1dEm4hiBltPUPpAARDumsh
sqhUvWg1ANxhVx7aJtb0QZHgfXVpJVCEA8N55yfJEXNIk+ygE5rk9jywRrrNMQfP
/HF4Ev+AUefC4kXzDr+UirpPAu0GGW0Bh+d/40tThBWnO61qsoBZwL8nKUCKKAfG
WcB2VPiKeAYE25HqvbkoZmK0tHJWa4P3JBHmkPxjmHReufDd0HYZX1R3vOVnUp6E
QK/xckhA3blhjJDFjxuOfZbly41btJfDBdQCv+5C5ZwrT/AyPyXCTlpZxy6d8K5M
FWU8g6LCf43GKwPxnk6r/IPwX3sI9Ce78rv7r6WkI21phXMa8wzq8n+tOf3MSFGQ
BbZm33HYfem1gWviEhgl6HBX/YRPLe+l663P4f9mZvmwGejc6nRhRtr7egXdiCa5
imhkue0ITlCurl6ZR6V5aQD9Aaj5gMhxPsY5Cze7FxRjdLwk0u2km7iIQJ/8UCdn
7/nvBMx12Uo/A1nr4pMyO88PRvrlK/7y8ULRMa5K5A4GrXt/ChKqf5TmDvuJpw6F
0Kze28QKgtkR4fmreCmdaYBAH09D4wtTa9VWyqAsZGuGkkB3IMmMx+Knhbqez5Yr
lVDfK62oLcQ8oLiy7sOOk2kHJfTOe5L5o9Bq1VXjJLh1H5gIwF/A2Dfxe/+c8xTC
m/9Bcz7heaiPLS0KwSCcLjeRSgOK1pTPimmweSgpW2B0GG6YJMpMyLnjzCB9aJyr
3HfnK6tKvLF5/l6GHqA0BuXaDe6uqzFCZKHYSM6Ly3HDeDTmLv+lOyim09isuKGw
cqDQY4yhhNJukpX1qZkD7lCzefBQ/Jm2Pu3EtD+dNuqAXngy/BOC5INeZ0SAtwEj
FO0kEjdBmI0ux9KoE+fHeqxPhpjtCVIRgXkZcYpAhL3J9l8Upg5pZUmCeDB9ICXk
3oWXnWWhIjplRP4v/9Mqyjd5QggA1CTUHG0AR/M+dZfyMRYXOtoVWRGExG9YhRtF
90B7r+UC1wcqWUzMro5jrr1EygokeFDBWiCauoHA9WhqdCeoWwJXYqyS2n4NQcP2
CffRuI7IGSVrsLMxBOPY/A6qVuZOV/jNLjZYk+8MFMr18IB8h7yGlpqQfBoH9ZUK
Lna2sFxxT8VaQyKZS48HxNT6MwKlDGqXRFIfjvVcetTnY7DCJKYfGvRsLj+Qcv0s
LdaMWxbF821Erj5Ofur/G7/Fu/9PuMfJXX+u/3QjzSBic7J6P0MISZ7Zlb/IMhnZ
F/fRfByBPn3rXhHVtAD3nltdW7e9KOCgjEelRpo1RNa3/N0pPSVEZgTZo9lPHN7Y
Aj6Pm23bWhdFg9NbsPygFrhDaw4C4JR6VIlDLHFSJJdnMOKIhAuS3FYFHES/dEuK
8wVYuCwaB8zCMbJZ1vsPKqoQ+pbf7yTntWIk8stUatm6ASgETAbGX7TWH/N4GTKA
mOWqoBt38eNZIbO4loX1H9Mu4ARxZWX3VYkLLJP90PqIVJXY2jA+8rGJ0mw3Lzzk
RA5UMNp+lcKFDNTGpjjvQAvH8unDpHwslep7Z6CHX0KqG7rlaiXkz6/Ga6laM8ln
EGAILAzHrkqOpo94buDgqUaIUYiXYKkbg89mwljN1aOqbRYk/QPSdnCOIjMotoS0
RAimGUID3OMsd8M6+HgC7jGK1O5T4Qkes/focaqg3B0m+adhNnBfgEKH1GpwAHVe
E7p46cmOND6bVozFH6J1tlknSSRjGftDYDOVoOy9mdRLCx7Iop/QNWfyW6l7+7tp
p7hPfNzRYE22Ko/DwU5R7iP3zT3HxgScdv6rTllAial4TtLKixkoOZf3p2/n7etu
OPGuqcz5m2MTFR65QmFJDHShZRfo8IWviYdYYmHM2DfU3dZE6lkASRz9fAiRtuJm
Y34Hvnpg8S36Q5KKTDK+eDxHiUlRP84NnXxj+vwpa+xxL+J7lP23gY3kapdBi7cv
sTu1AhEjA9oIRwehNJ1VPNf+0E9a2mS+ZZZuA8wEednaXiv+vRRnIJ0kGKKATZ7z
336sJngV4VTmLYLBFkjURDA1O7wvM4SgyyUU0aXY9zhqLr86QJ2vCuyS3IyLhCl7
Voa7JUsLiKegtUJrzbIOWwCOtUexkRfwV/WsCUzg90pDEP7fMgGULArLoOOKvs3a
VI+E+zPdTBwMT35y2ijBrrOGfc5fopewoJsGQjfuPjFbyrRKPEFTb4FbflMVtz8T
wcdK+eLUJLjq3Cinn5K5jLqox1+tF0wgJw0mKh7fVUPL1f/ywt00im0Ba7SdbpBP
XAQfchPBxR8iPVuzuZWPwd2jZnt3SrwzZ4+kJWegoYy/v3l9qz2xDOlmQiDZuQAS
oaF5tw5REr36BfFMksbpmwcCD58QL6bn5SxSKjpWLqNUPaMD913+ulgjlZvHqsgJ
kZeohGWm3XnPtNojN4d9Lvadm2Gq4cfBPCKV8usChYhDkF5rYDU5rARETqv6Lly2
ocvE6c8lMdjsEVXSnxbOap9+INW07Rtw4oZ6QBRBWfhjRlj02E4LKs/VgdQjW9o0
CdaFQyPb4UDwX0D3gTxG+HTvv0eTcpuXv0hFa7UBvj0N+41u1k39VC3/M2S9xmP0
BXGhG3JyGZ4eQ735CahWS2fv7gluam6jdoL3B564ufFho3vCgals13LbDqVsGTVa
NcO63SKfhLHfNWcNDjusCDrdyBF89ilAdasFCkP/Jts7teDTBSGCXOxp0hZdpkWB
dZRMik5QVzvHIF+KjyWahnbTEdYgGwb9hJ2V6f9qk76fpadutbl81W27kfe2V0sW
ZzEtGU/AlBUVSYhwEI5RvRV69RTAlAXF2P88lx5ujPPAGck3N8Jf4MyfRzph15t0
OiIK9raW09IEVC/Mc0BHUd52E+OpaYDdds3bhxmO7kxDt98lzeM/MwmR/D23I1T7
7j/QwMr0RZCQdHjTTCrN7/BNuWe6kYLsItnoOrsrb45BT9V8CNbPy5b4NM/oo3SQ
qTOaMPDbpi9Et9XogzVO4NEUJDhm3jq5Upmgnw58C2+aAvrE/xsM6oMqGupXdydJ
Abenvhzhje2aGlLOWjwqs/H1mCSz+hlrsxHPzSwesul+lMtAjV/bhyk5UAVw6NSS
nH+xHzrwH2bLlUSUzipNhGZtUgS8YzMX8wy6BbjAe5n7hSkOnJpQQxri7LLWZOaL
gJzzRWQlfQBBDD+ngK7wjIkYHu+WvxV/b4NgZeAEJ16zAMpWtzjqTtayrs0BKFvB
4B6Coxn1V6IiKAryp9rnXEjhKxdtJ9o2wsTxdin5R2fQ2dhxuSThBNRT5prk8xN2
hjEAy+WSV8VZLfgIp3kkMfg2lo2435zhROO8Eu9TJieFi4GPeA6mGRjERisNjHKi
3puSy+3bUF8mZFY1V3h2dj1XIu5ZOXrnFs/5vxjSzgIHISkwdDms5RDR5ZKL+blw
kwYRs/skjnFj8YlNhuTuhsfeijnWg/M/MLAKaxgVZs+bt6OqmDNlFZrFFkdlqxyw
Q+Q2g31Bw5scsgKyj1/z5o+0Gi9sadEUGy7py3Oi+q48ikGrXkhr5olpdZFP79Ef
gPBKqJXyXnSm7nyCP1iiSJBpkeUapW4yOd0K6az/koer5M6lS+Xu4vUfGtL+667v
JQt6rs3tXbP+V9/ecrZCSMse7uWZF6zC+cBPdZBmR4w2IC6hfZN+xJFmi3l6EL+T
MgrhCWSWrz/IiW+IU000D7W1WKy/w5QUE7F4RY2tVjyCQqTce8PmDgexO0aCgsJs
NFe1Pek3mhz0W2inX1oxEr3td5pajw6DpRfyg0Za/o4457bvL+d4t9P5olYwoPOO
DMy0FJ968+j/wPMFDijwyzhR2NAcNq+rp5xGCdDpmYdMVSIb5BGwwQQUyO2ZWN1a
57UHiXt46gXQy8AHZABS7VRxP+r5q+P2dzN45c5EhxsS5z+Udv11yYvh501E5ud7
kbFlIVdxgKEZAd0ms+RFnuBP9tTNDexj1Eq1Y1XEWmMlwW8Ts9JcePGZwkAVg5Oz
oWYBBru2mySBtWYixCG+/LhlaFh4xhikRxKFaSlqpN6RHvLM2/3N490uHnQutzN/
DgK6QOBdvfdqIdih/U3HiTOTSn4zzqceAZ5Br56KZ9GeN8XCxwWQDHyTzZuRirM0
4QIJdERTxRDyB/dTLnByRCkUlcMIy1W0BzCYNyAfAHuqFjNCmHMGal6vOOdzF/XF
/I2YMW44p71NGUVDBju8NtUzzwFFFLrjfUpmRo92VTCJIB6Ui+CwzkncMdRCEZu+
Q9LEmF0yNUeJycS/0Dhd3FqR5LRIQsamOV83ytnRNfu5M0ouPttois0i7PORr/tk
Abg4SC6mizfP+oAixEQ+LCwJqRS4oPfu6hpRRWVb9VcVyqsXbt/nISMqB8YdSZyZ
r+5euFfr09VJa02xKa5uM0K/XQK8Pqs0ypJa+trSYo1Gkrv0iTmFGEYr/hW+1Gr2
bYD9Ia4y9rJpNaBxnpstI0hLILaWLftChEb5E+HpPG36K0E/k1wjrntL9XXd8SqJ
OzZs+OJ8xuw1TXbPWPoSp5ngcDwpDaAFp3AUFTkFUKyB/4cDqc2bwdnJE3GbCtjJ
Fp/PKtbMPiy/XCPHjejv2b43qiyRSsdEgcKd3j2SfyXuCTtiO8kpkSSrFXqCAQrD
v6oMrhMdlBhWTdiHhZ+1FkPJGRvt4VrEaKKW0VIMvNRINp8xwG6fDXizviCazM7P
yc9/YaNNR+cIxaAtp5JfefJExNceJH0Deuv3FShDAlSMAaiKk9SM9/jTlh5ekrVc
DBjpXcFUUQJ+bUjG2ZI/DKPEoJPWRI7lYVX0PTDiAO+3PmT3YXeqXQE6B+0OEODN
TF7rfZ9kuu5UrVa+Fkia8NTVH7/IQQ89hfTUVzYy1rjvf17OeONh5jWopqb+MPh0
CfJ2zCAhmsjRmrlz495foZgNrS45MPIeNTkZMZzDf8x0UJtdCiVEEJZiezqxxKG/
JPRhh27HmQ1zdb02LHqgs/DRIawQUOkgMD2BPuyg1L0tzPkp2DJ2vIUeT3guf6Aw
hlhOYOt6eoJpRIJMkoeVRGFG4DYrA/tjkcpYcZgfkfDpu/m1ROERXurI0ergalk5
TnpyscKUT8tn1aRcCsW1czyGVe+ZCmrWEVyfNJBvrljoWKPLcOJCtXdip9f7CWm9
T5qB44N1neKUZBHkPs6z+2bwCr35CMiA3GIJaxKUhOfBjTi/N/hEVAAPw0dAazio
3Skz/8lvo4fzACTseDk1p51Md8XCOH2VXqJXa4/+E9XNrdRH5h81oS7gsdgi5XGY
6Wtb5EZdHJH0eG/StvKQ7AFdAT401oUrvXtxNjoKfYnLO7SNO2bgymbpNX7D58MH
j/PZWs834133DAXII/YQaw8VX5eEzECCeH1X2wc7Zb9S/tRmsAU5B+Xif5M+6fFc
4Qv1RiNb4dG2cKHBtKSIRto8zNgMRvEfQrHUJKwol3Iv2FYYV/5GAApK4/ZK74a7
uZ0UZsnnJIRcXGYINfs7P6tzMLbPlxLhG7SUqeeA/C89exsVIEhLiJIjwESsD6af
O81CIJcuZ3JGYHgEBaOljwXm+tWKi/Krr08vwvKvIDLys1K57tczFIQBbc+MIh2a
glGAf92ADjcnXoN0qZpB85S0K6+7Ef2YgylSPFB57E+yt9EStzBnpI8+AcaBMbWt
0qoJtYZS8ZyEKGLPGqIwEtPGLYlcIpStr5dz/qB3i6D7GwhZPGGXeDzSHtslDX4i
Maf6sjtAK+eGULtGYuYl2NmuNHuzI+yoJqegNsghY5OmykjdViGY8Eo6J5KmbHXl
2wZw2O7B7FJ3NBGw0Y6p0/ags7mtVSo0gwLphOFt/67RwuQTETKfyXxep/7l/kLj
dMKlpZnb5RuUAbVQ+PhnFzDrcopIw7z9LEsm1p37UbjzvyBC9H4BIKdNEZL/oJpt
54Pe2i9w8zsO0QO5vJWyc4K+AGcqh/aMc8Sj1blG6SXum8/1uaywPAbWA6hkMzVO
74UT3a6n8s6eh1fzdQtjWVghL6x9oCkNxssRmdJv7Xw+FH4g7P95f1z+bFXHC/yg
3u4DFbaM3y0BGXMn6UBXkiTt8zPaCOfaCs/1xmofqpqxTSNOeUxRMFCWsJBD7/y+
7BQZEUZLlyUrTNWDUnpxJPV7SjAfyKRGdBB+wTlazkQXyaziPJMM00kVTjB6o/F8
pOvBKAVH6NG3sYPk6xwFtw7cZ9atvaGg65cq7v1n0bJz09DhHCcCM4QApZcG4P84
s6rznnDnOVUADa37ZR0aJHDmnrZFSd/WlAHRgMyrxrxpomxdzbGwhYwikmsXTB6Z
LRk1ZhT7CCO2uzGf1wQbJsdj4rsx0wlwJAfxBH0JHyRJ08kG0Af5/z2z0ikVEh4z
URnOXARCqsD22bmY/HuAmW5cNVUEDYA3hkG0jf9SJVvhvoTkN+3BaXCJyHo2OAdU
mj87OWvweD7Jg+rD6Z+9YMLzlFJ2Z6hkX8OLxIWEqqCTK2TgcMj1mF8IkT97d8HA
vdeAwcm1hKI7u1fG49RzrD22QonXF9+ZgpENO2u2mLRC/7d5dafv+LAYEjhLi+f5
pEIlVhXd11pl2w38hFwDa1q5FRuF91gMMJNgqulTtj+QuiuEoXL3ogWpxld6U6nQ
tWLiY8tjDXKLkG5PbmdWfYzvsWAVYOfyEOHg9VOm8DcK0Hq3jkxB30mfvlVdgj8l
FCfzM8RlQWnvA6xYd/PYekW85CUxa1kSndwBCOKzRIld3K5xQvwPP3pXbYPTmSnO
YnYXRpKDNBjylXV8uvXW1NSrG+ppp/b/IddwY0BMVhil9wbSSN5MdQtsswLHiCte
PcytrTBD0mdKuY7kDkX2hNGFxVyCPgiL+iAEwV1OwJk6GGbnubz2Ibaw3yw1MdNO
6W/B0IePzoe+Z93bZM6+eLDszxOuBkLyon9K9Ait0WpMZUdkda0Oqm9tt5EYrEYh
XmkfG/44cZHQgQC7LJfNsl14NzRvyXHQl9eyCoCtjzRdKwajM6ZkovnuKzJwjTI+
rvDMLhlrww2MtueJDzl2Wwc5EIuTKLvru84h1H9FVhFeAdVULTa/KcM5+JmVBtht
Jn8IcyXd1d0uOW4nbOrL0GQ5wrK6xPmG1OXCd7zyzNAUfwbA8gANWsu/t63DT6JC
1JNzslXZk0StS/yK+7V5j6IiFtLJxBUdvEvBMXz+gXxfZhQLHi7Py8q8oGjGIcu2
JmgElmDS9ODt9q0ZXkrPiLd38W7+u0nKHRdlvfK/bwAEa8XdaDzE+Kqkw/tkjixI
dtkHJZtkfd6qiuSiW8SvCY4NnIcCxbnBbTGbxzMGml1zR3waOAlfJ2ftBr4NiIPc
zZzIjDd3EkLm5Q4I6AQqzWY0W4GzmDwUOYBa01fAUm3mshsCNW5QBKGFFEhpgkEv
CbQcxfNC7gKG5mohZAtGtbQ03ekMgh2oYzP2hCwlUfD8jLLrJC1NCQFQ3LhYA05u
wPbgI2R7GbZOvtgT1d4aFdekyq2YICgn/S4x9usU1k0BcbFABPIUTONMLg0yPKyC
fxvR2vEqOWvJuD3Bwwn7k4bz9QMoasjHnwaM+9n7kJMurWem7QNW+oti2YBIwCZ8
G3l5N5bXIRTNHAhZMfY8ihUqWhn2+XA8F6LnZpZKVYgwdnc5HFZ1Hn02ixucVnm0
rvgM/LyqX49gZdTFBvTi/IBqexiKYkA5EWv32CUKVbYQtuQdjHyvP3BSvBJiIW1e
tpzTFqwiQrq3AFeeadyPQlMWtocqtrWgkmY3fYxZPp3GT2HUzrjkosaHE9R2b8V0
SCrUXFUWxVu7GMfaAqgYACz0e/N/uZBFsx096H6Pd0ahmwh4gvckOXsDbkTjOnvT
SkWx/+TTSSrEmH2bhtkb6Vly9FIZ7tIdjtvKYbl3YsZQjaB+Vv55Vu7gTm7GzX6n
NbaIijjosCc8ECgT90Aq38lkV0txvg5OWQiu/zFwAwjb+0R12MAjym/OrmOAvqjs
85bjTvMWHEgUoN0feeViSW04NkcWih/7VxN0x+EaLlsHSj108QsoTHzgsWGdVm4Q
3wJ9vGPRB5dZG9fWMx182YWNxCHU8GaxK+xtXWYWQe8Rv+r6ugj8uoQ19k84oTff
8ZAFZVUi9pGtfCInm5HJpwovIjoCdHNy18zj4DeMMkyLyE96SkV9PW4MOD93ffEP
ITAvfPxuLOa+JrhwYe1y1m+/o84zwVKcHZZDEOto14Y51Vvp7pdH82kOJkLYQVws
fA5iURKhAZDyxgX8TL8lAqbGYYJ9Nfe6925vOOgT6skxBO3+A9x1uEEHyKG/fzdN
W6BhSP1x8VBHFg10FowU+rsu6SkNHReyIglzHIQCUFw561dqGI0kJLKsCbqnWC8X
7aXNUuX6/QOgspQIisB0aOwW7dksURENx6/HA1LrW/nlfQqlzLB0PINj4UhGHXXN
koKKlwGqrsRATz6dSYwi2pSROOfrPwIIo/KLstrIlEWuGajqmwof1zZdYxbsUpD9
93CHclIugQngRqXUJzXtfBT/k2XZtM3DGjUikBgti98+EE6A+oCGWm7nrX3KrZhT
PF0yWTRnzv8RqmpdQQE+Gjq3pVnX4B8A/5MWdbPwh15D5NC0oJhQry6ZIEDQXjfe
GVa9ht1slg35nGoWgCVCnlFCscFvqKPd30N4DAuAT27DrpPChAK7hRW92waDzl6g
LtVkjCS5ggQFQTEBiBnmsuJkKkE9TmC6pHpD95UXPdiy/AGbPSgMDFrI6IzdMBkJ
oUCI40YY8RxoYEPdJKtXMFhnd8J2YAq6K29uuCrBr8c6qIw4faC1n1bIhFP0c69j
1AuGUd6NIkMNqbbkdn1k3tfwqbkloRmnm2qe9Qait9OUqoY5klh8PXVJtUdPCDrb
hJUV8gOWXJs4hFJieGDSb+ss4v2CAltJ1Fb6EWQrbY53z8LaVgBGE/xOngCFi1py
zxPo1XQym439LleZxHlidG4pqQJgkWhg14wq9T2yMq95CVN7HOoXbgmanEPWcz+L
fcIfCyskpi6+hbNXuXIn81MINDMxRZDlO2T/V40NMnW6Mh3E40nkTGAKNgp1Nppi
kKw4Ve2HJxzYo+YBq6lt3TJYzMDDhLN5GLTH4F5dTst1JgqAhUucvGe+JcJKZ0rj
VT8o0Ee1YNat80ZIh61qmtwkSxLdbBYfLIDBkjFd2jj2AIxWdNdcAyHRPBuQSIl9
Y2EbiTBDf8EJF+Ijn/tM9RYfrfPkrbmJehZJctbsH3NPBPRus8/dgeZq5FOGX9sJ
99Ymkk3e9LdE8ug1XIpSDyay8mSI3S9wAA/gjbtsoCWCveCHQRv58QYvekYFpXra
GdVj2PrOdkyaQlMvKgxJjRVukT3kOOyTcgw6pZV+98uKtn5GXgqjjQh3omdg0QuZ
s2Y6ZYma+L/5BjuqKIvBtCmVkr0jy9y/so9O628HtSjoq+x6gBVHv1v8BmaRy5e1
vMwb1UjnMP4Jv5fmvDaDJaqj8yHNqjknbddEk7Gt3zPtS1/3ZTMW9noX6Hmt+6Sg
XkfQt1frOP4NWZpNRb7Gg3rGWsKK/q90pDbcE+JLE4dS5RS059mHaohReg428V49
bXPLabwSkOJYkDVh9xS9ur+ki/bgO5psbiQrnvmWjr5+OJ3mOYqEfMk1wrpALlFi
7QN5D9lP/gW7KeA4zWQlzf7pxGmVBwGhzIdjRSVy6QtWQl8Opxw7//YT9OTrAWzb
IYp48nqTTM5gh18Xu0zRT2n0nvQAQnznjkOdZfKeQCu4l5d0EsoCnLoiW9/UbFjc
6yR8IsXtpBNaPdWPceGsV5sg6s72fdqJc0GUNv0Oo7qrcOQkhSAhaD87fFyPyF0D
DNDR5iUskjn5m6CwMJFpB0FozvZpRSer8tpEYkHrkstFdLBFrm5JQNd35kpp2ajn
FGy9MmOXmD7BCHwOXV4iZ3Rw73on2Je/jHO+YqcEqeD+pHNursl2jl0Z8LHgPtyB
t5a9oSm0BK6GIUxDb4dP488pWEnFEbAptX1RqzJ1MKutvuuLHJIJW4F3MFCSqZ1y
eHKcHoEawnrcYBUHqDqZ/8yndrW0dcqjEaTDEdRGZ41EI+FjR4sRYFBG/gwSPGM8
216v+UnNBBOt3BWTJcv1T7zgmj29Gi4tOO0oKOOWGNDej1HNjAlhfpCDrx/CJdez
4zo74ENSD3t5ams/nTgQgrk4bNVjUGYY+5BnjHnavhUC4ly4crnALJhap7UtgdpG
Hn1nyA1vqIjF5HTlbUnSeYSLq12RmWbeDaJpileRGrNJ0gC/gWXG3cPt92WHtkS8
B+sKEKpmJN6sM43VlVfsYe3cX2v08DTQ21FmwtZf6aa0zrgQCP9gW+IOD7eKep3a
3XtL3GYIR4Qi/rhWOa+Nn7qAe0qa84m1mW254P3S1+ijNCS/l7akwCpop9F/zbT/
2O8jS9qjbgtmY1chQjq2+E8igh1QFMGwj1daDYInr9K4K9ZcOQBJ/K1pAy5zd+O3
e8erzaBdgKNDdoAJLMWRkD9bmDMnMCbf/qFYXUwNcK8Y4b/7EaF0NfnKH8c4SxGm
quGhufg7Gct9WLDwDjhwgzpSYYKSF/6b0onb0zuZv8uxssfPPwJTmwWYzJXSllTY
VdxTiZvqKfquPMvJD4J6HpSpyLzItpI1aNro2hr3hdgrrx21Sxe4Cl+jbB9B+BdL
tbM/NZToLVjTGFt3aUHnHTR6E+GKYulhaFb4VCAraXG+LWkgUtVsOl49D7a2ETOF
iCVyQDwEK7CKfYSWZOL+sGPMHBObfRp61bvn0ughqsqVLTKbCpoabJckCWLf2SAp
E+Egd/NP5xb9wSZjeyciAn7Lp8a232UbgAcjpa22rE1hYTrIV0WASR5TX8ka6Pkr
k9tGR4eqdcppIr2bH4w6c9MCPekPUIzXW8BulvywKA+QAdeow5X9SF9fbz2DiP0i
sR/UzDE3fe9gNX/4LcQ1DNKdqbHG3Ishy6UOD01T2NjtkanxZW0QiaZIMTh8GraB
nN9tm0WynRo7fRyoiKGpJXI98uXhfcVtfXI5VM2Kn0Vg/1QtW59QOu6nZVcX2BBJ
t6VKMGLr9EH7n+VvyUKME8FMwZ88zosbqlhylheXOmZlLM6/miCgLbqagDowb4ti
aUzual7X+XvTO+HpK97U6n7BWDD6q69C+XSUb83cP9qlur8YLMDfxwsSVvG0DXLy
VJxkQZLcJBGIO+oPu2kUKKTLAe0NpuAEc9pWbRp27Mqsy9oRdeioqUkr+0MnUOdI
t7/cozQ56qfvbmCNx0SL09eAD24lFyCatApLaXGVmdhUapORFQarupfPJGLJXNZm
Do9ql8nSQVh1PTKMPFtluevPJa79oiFjqDGVZ0MwAOPMC8S4kKY7HugFzpsOPBoq
bmm27+AZpo5rVOcjtYJaw3TAP6Oe30T9cu82SYXMGP5abSxfhGzIXOywaREIPVv+
3tq5kCE4Z78lpQY1g18/epml0CZfYwwudYDHN0rk/CT/4nHpDhzBNesKORoZIlBA
Fxa1klOT2MA3DhuPgWCRz5qusKd6hcjRgRF23NTBzuNWxqdWsb5HGKer+x7FHhWy
0nlH0uX/tThRdwEw7XNyx1w6Y2p6dgA7MmCz4OIel9aJ6UkIvjUlGzMA/wxnFgqC
xHwT2a/h0BNcsFuVAlBQz66RADKQWaBS6dItkYDykCqWuifh6a3mtXftodSZxNCY
okGNKBz7TwDtBZSfsmXexNpdZGegem1tHTnb7XBILktWwZ537tKblYS9XeiLW3Z+
s0HoYZOjzYyM8ehF+q8GRJ/U+nsKAUm+RTIlH4RSiXyL2KCZfp0F4xYJ0CX9/A17
sdIQTKhc+lOwoBTwPDqPfuP/k6CQKYn+ef+zvq6u3qDe+AfVVanaIp0Da9zIcgM1
TXMJEbYj26EtzRm+rmY/kS1rRiNh3KzUN39iMbnHgwLvDrxEXL+v5blaqFS/KoBS
iDQQXKnQxsbNw8EVtc1w5yupTdVbWSHXGAHSrBqru2MXkx9Ev3ijuI7IzDTZksbD
jywU/4AMK4ziGbw2w3/Ye6IHkjFWSEzibOavqwNT7xYkNOnDlRTsLpTW5ykN9dFs
zm/5H+js7MK81CCMlGTYEXOMu2+UXqFD7HBvJvqVPKxY53XuhFWYB/9SwAX/qQ0V
R4cMpQVcCxs9pR36aVjmDfr9fW99WMgAb3m3thLaA5ESEXzN3gqKDKe4GChtmqUs
9ki4KOsgTUKfu5Ge8b0DIuFo45XU99me0MLeLKqQrBCehB78T1k1eeHjYZBXCn+9
7rH9BHZuodIdIRMP65MrGkHO7+43MY7wy4x6xOoykySBsxhnNw5x39Mp3b3UWO/E
yTJUAANS/uf6vQXnGzz8WxJc0YrID5adsdCux0/cWcmansq4UcIWgLfAJ8pCnxFa
dOPGOsBAqLAkN1NZhav3gzYs8IQgf1r4mBgPCvQzRtmQ4eBZM0U7/zGQn2o8iZe/
hTmbv9MiX9Hq91yo421BEsP/qPtoNEmSxbuhwQ8ldwHxT0O7HIvjBXfPzyXzkGLR
WIrhaVCtbsNdsD8lLD63eX1DeZuC61haaElSpwxsv8Z0SkrOQXSDIcFvCheETydm
XaK7Ywb5+OLI8NPGwuoa6wwQwzrihwc4Tes7K6nTtatQDpKMmj7sQsU9TtuOFICi
yQ3IkcHSuvbU11z728fiESDPqoGUZe5OGk8tghA4VZCWKTNiVF47SgQpSdC10sR8
7CbMgRLj3lPuHAZ6N4Sj3uoxZTEShfKHuLLIjszTh1fuVaQ5a3V+70iwLVbs65sw
ZZEpomPNFlxkNDI8Kz2Kyaxein6uPW4aUfECMAcxJqrbY7/nOXosszEwXRnP/3r1
jXA/Pd5UbKbipStQwHIBYn0fuG/t54W6V3UErcD29guJExl9Caxkkp2YZxa04b21
BfKRhxC8g7wFSKG9B8N50MmMIKpXVDyfyq/HZlUB1W+ZNt8cuD3dImnVQ0RMdNz9
N1XUbeIz+UGE4v8wzPQwRy4WBDCR9GAXqkx4Msj6XncdsHlRHRXbuD1PyVm6TBfM
hSTWM6lufSkmnS/0kAmL2zEB50m0HMBdg6D+OyoXqtzkcXrf1n4NUvG74yLXnndp
4gUL4uNzZ5KWBZqePQZE6xKy+f0iaqyhjyFnsqrEmN3kjaNdYB6Oo4AlXiyUR13v
LI4ruJhBoubhL4PeoSZJ9Jonk6khh8Tk8YNZ5FHERxXXNzwpdzg3L+m33bJM3k0H
oCaJ0CU0fou+R63p7FZhjEPCZ3llMN2I/mfhISTyruZ24HI6s0u918V4JUYtV3ym
o7FfVzV8Q/uULTf5RCGDPP76/uQ3gD7LINcugSAGndVMz7z6tnBWYIAvpH16X/mn
UUmLQ6Sd6Kp0h3KZ+Jl1TSm+SjGS63OEhDdPmHCnxedd7fPbZBhmF4JE1KWwFyQs
AnNxIFdK6Hsicft3KzWDdNcHgDFN6uhhYYmDUAM4jmhBO6hQnz7BFKfw7ZoDGV41
prMdxx+Jep0T9LvbgZGETlX80GhTmUC7ViQN66udP/As0ojfN114KAx7s9kLNIG7
S77zjcfdxu4FWtKF2xP6/03kdMbakH4+9Ti8VeAHvCI6lg8M0Io8PVhuRU9YnKC6
x+lsXT3sk0mlpOP5JG7PDLKHAKhEBpaxhv1ZfUvMOpxpVbnQcd5h18IAGU/udD5Z
hZn3zwjH47gt2oE1C+nD0QZvwevjvlVyz3d5+Lpfvdy2omy1Htwa+ZnEue/hs/pi
EsVVRn+8s5pNo4tqzp3urOgZLVUba38o/Dyb4gM2PDat12C0PiFoxtX9Lef57cuT
MaTZx53vLhboYWDuTG9xNSI7Llr8fcB749lJ+nSA7rfo1dh+ZMYVehDnAuCKWbRs
K2MKuOBnkOwxDh5HCB6hBMEWDyubdhWzdFMGznljIxJ4YJh1dFjjrbYEHus09+Iw
QeLrA5Nd5BrzBIikKF5dBifssh2F3WYaSIeQLn9J0OGkUHqCeH2IYhEQzrGZlfM9
GayY+mVmcSm0jnrRegFfb8PsT1eys8eaAi51bmMGLOsqJ8e3YE5J3sFRp38v20ac
sF+Aa/5DpGJ+EBA4JUkG/tFK6LSJvVVDum8cKBlheKoZYh4x1Tz3IdLWk9whi8Fg
o9pfApOyVw/HOxaz81xGnFLmndsArR2fTDf95u6kBtNX/O2DvrS7PzVxYI/wh2tG
4ikghz2iW9kurcz5ZzLl63KK3aWk62itHyHvJYYS71cZ1LtVINU5uhcu1iXpWe3I
wKSRkrruZ05oCq8JKidoYZbio62uJ1h5P02GTZrfPm6Q36I1mVnqkVrM7zjkm16B
7IzyFAXIbm171+ovsMRoeNkMtVAY93e0dKUs6cNGEzI9xJ5KlEaqj82BcxvbG/Z2
bIyu3D9NhBspapWpIRxUC8j1n6YhDRlmPlzRlpNh3zHeON3iil3KWCwwZtFipPq3
8/cImJOezgCqUWbfdm8/+tTcZ/8TTjeJgwnz82dkZ0dcprOL55B0Rq/J8hoWxqNc
zhjUy1fYT8sofeoqg5lh/tCilrIlYFRX1z20Ij9e2NA+x5eIQ63/5BIbzV2cntRl
2ca2Y1ei3xa7yFM26pqvt2l7ITN0bljSlHO0HdHNhSpngFDLpKRraEm7XdjIsnNT
fZuvDUr8zuyfis2G/XBzV40KySq5Yy0xFsnUwN5fTTt0IIKmHvkFCP1SXSFSztSa
hiACrIwsgWMQ8JaO6QO8lhPtNLDZY4laHBvcE0O5RqHavobKHl7n7bw1NjBYLE+l
jsoCxCYZ1Cv88oHnMCYIs9sE9DMf2xo4a/UQMlzotPYoJLjrCWjr0n9S0g3tPoTv
VFpYFtjdYPRA9BBb5ZiDUjcliPpMCpLwvZbK/BjbgQniKcCmU6hewhyBbrKunMHE
9PN8lE50cPdSBrBWPPS37WoOa/lkin2UyFXHIM99pTyIg1A4VUkZ/BooD2elj9iv
O4d8K08UZ94iIuUankWyZbLQYc7ohk2tILfogtCA3hUtFHZaisi+K/jhw7/ndJ8q
WiaNGJZ5BjoSxEjwJVDsJ7RX2nn8eNAeLFg6AC9Qwe2UHyjdsw4gKUlaByEN77Nx
F5IKrcSYPRaEATZlFHjMg9rQkG3h3sF5o0K6kRTtwNV1Iz9OUf/JSzzqIijE4Nlp
qrkBLen8wjbC3Q0xbbFJbqjvVQQ1CHMIZ2QfdliqreVeTeh3t3S0ZjLSut0637F2
Hmd1SlMmNVrmRvC4AAZ1EK5m8b1hxBgy/3VFAROOQnW+Q9WVim7pI0hvHAnVmBb8
98e7QZrwOqR1VpaxC03x5Zuj+Th4kzJ/JRDMw2m34nKBpdR8k7oMpMD6qjlp4BTo
LteTRJlefXDbUcckM1RH2D2HKaiSv7K0cguwc2x2xLL61TgIecbWpesC19X9Px9F
KmUv2G285/qwzs9PO08A2EmXg3awVytsx524qN0gZ0M2EDk/u0lC4JIV3JR5mczP
lWxEPO+ar/xxqZ3KjCNk7f4LrH5Hxh0kRlRMxw69+1m/MBQsPQdwTRk4qLv9NpZ1
XI6EQYlf1NVmGT1kysfFf+7IEMR92pbobLrvU0+IwBZu9M5wdZm954IJVaVQd923
z6b7ncrAxVLKE2VdJa9CaGVThlp/RYN2jyoWF7V/BOl3RMXqRGkpgdq/4PGfH44c
QOE2gpvafh/hLMsnR6hx8IFNNLBcXzzlG6D1bPzR3F0SqQoe3543rfHr1nZ2+XLE
JhYpgmN2TUyAN4//C5ixW4GW+MQ3CB5kvHZtn3zyYRNR/hRGurt2qtVrDx/g95hh
0HBZMsGkSoghgBkVuvmtk4pW8RAeMz0wm3PqO3TTLpRHnoPGe3kiL5VoFxGdL8Hb
1+MkjnXF+XcaSOd0F7+MgReVEcUKGrFXUl1xjurWECmJI+Ip8xDuqFS3HLq490ZV
CpdopFovMs62uslPYOlv3qI/FAuJDl/7+4/qUyLv3kTyWmMJ8vbfbROzi7AV1aVc
qnHhWD7IzsHYBdhxaYs30+ytwNNjygnwbWimiBTLDp1ADT78FvFQoVsZGFHpGCqy
NzBnkIEKfj4Spo6wdlYlNCdTmjDMoiEG5Ls7OfnFBrv8GVDaBNSQ6WhwTnsZ/CEs
Qhew+3GU9gGGVjetV1B1WfNVKZfJi2peqxMjT6dmFkvU3d9FRaA2mfwAX53jUHC/
GMc+V+TzZO19+IFwyQaBBZ9Mb+iahYT6KI+WFZwc+bdpmelAs9TPRrKBTxvTGC8v
q/ZsmGJlhNBgkPhjuMPVmmWq8BZGhjzlOXoNxnxefK3nDpEhFcX+obgZjH24t1aY
YvYovsORFSLezANEWakbOUzRv+wTrRYNfdsqZKofiiuacrhEEiOfLUPjkLeCvcMs
YQcJTiNXWYb9YQbfl3aTssbmp9CUytdtjJpQr50pLQySn7kBPriZX8dzZkT6zcu/
kTTf5XlI7uIByNiYJIkPvzoKgZK9TNGw6G2Ei/YBH4nQHH+CPvM9/ge+nPbKJOGv
x+ggKuO4gdFcwX/rB4yfJAIPkx0D6MDcaN5Wfy18i0O2gsaaW8/9KqPVqhtZAj59
9kdny+EeouUliCPlhdrNqWtXHl2JD31panywhOGpALhslcSRQfAhjXJ2Y2lXg4Ei
G6aS2+aCOMqUFu+gunR7sEIQ1QQXKDF+y7Xf+KR+RlDNP8+ppI4JWjaTcQY00ISR
rNDaef/7boo7V/DiG8Hqc0ih+VkvE5NiSARGSv/dvBRjKg68zNebccey5Sl6QzZi
u/S8yO72ozW3lb8wCWQNev3bwEllUP9SSsEFw+Ue4vHPpy7Kh5XDGzcjhF2jooJv
eqOw0CbRfvYoDYxFxASMypm+HnPifAdrXR63TrCJdMibRArkKG4BGc2ffd7y8mbH
yvmELFdoKSthZSAIzioP0NIx7aEIH/28qWH74ZoHOhYNJiZtSHBIl1gSeeOqiZ2w
G921kUCDaYHqtIKlV3RJudCfBrxFcmw9BKDq6KlDDzPVnu+4k1ChE5d9ToY+ayE1
wxbdjOfZZWRrtPgrRu+qJXosY55k9YP7TDlSZUubALsalONfq/MZnfoYM5Mja6sw
cQo3byyjMvxwiBHsn+bmqxoNTG1hLvzNCpbiWjgEULciHc/MY0WwTsFyDYFTSfgd
VJvKQrcZGkzkzIM2bOlX1zRNw3zQUnYI+fSoOiAw8AZaBQaGPsNs1qy1AQxBLtBK
+eOFskosmQcwdz/Gw/S/DxdYvTBln8osZFLOL6SzKAS2gYQG/HNx60SaKhTtaZwP
jKE3CsIfpV7bQ2W+CgSoGKOdEiJ+3vzNUlrornARTucC4Y1s/h9eIybP09pEea7q
GCFJvFiIedp4oBtZuuylV9Lm1wsqe8ie3QykfyA9cU8ZS6NofIedxXGs4YZ7bLEG
qbPgTipKqfHjo6xlU2SJv1h5FOR8gHqWay3Va8ZS3GnOZWn0A1rtC0/oM+kg3kex
pAczVyZTdzSjIvuwBdQyFHbXn3s8TO9BpLcmQqLCbaIKuw9pa3M2RczpUHv3rxtU
39SfvQ+uDHuSvejexjGY4G3QTtUL7ejz7leJGoRGB+G65qM31Xn9jOxPVtt3S6Uz
m7khK/RMrNsdMPlbBANqZ1ACY+qJwRlXyklRuCITVje4zQdSZ0IBuHlEAGwlTvJb
OByy1646h+HZaLTIk141OaWMsLrSBjJwIHa35s1xPLDWQHcVwjTf8XHcyM0NQFH6
BPyHFeUCkH+m9qrnusKHoU0ug0oRZzQxSRNjnoKSekyH0XQqc75nbAzuxhI8Yhkn
pQ+LgmVYOH6GqJ7yJF7Fwft/5eACoU3s6DfAWxJMnTHfr64g4hwTLVaJDLBX8/pe
bKKWA8kqZmTXHiaKiuzKsVd6Y5H+vRja5K0Yh+e6MuufkYnGxUdmV5wYA9E92J3O
2EQwihxCveeNjsV8uPhO7qM7rKWh1BbtOe5vs2de59czWM76x984IK3zB4n5LIYW
nIdM6Vv4Fz5+cjAZeLWeiXcalkFhawhNLbmTQP16krMAP7xnEX0v6XTdz/8KW4BZ
mPyF4fSCNBypjXoqO6HbUabw/fxub44xJ50qZ75eflnr2MoLgAJfCMEsvurW1cVm
aMJY5B3e3laPT1xibRaxZUUfvs7mQ7XP5Ol5JCh7z1YxSpOum2m3/7iAKiJ3WbRX
RrppCIGQ1lJsfzrYdPI0Z9fN3nfp6UodK8P+0vdnIqyq+p0dozyH6SMiVVYxRCs2
qNZox2KaxYXlzmUBaWlxoA3Ru1k3TXuBvnvH9glr7eliuFMxEa6a4CTDdY0CxJpU
FLjRUIIsuiqgWkRY3OBqJ3Rw92AjmX6hXO1xKE2f9vBSKZnvO2RGVretbHkU8K63
lNtuog3FNvgEUcMW2DutpneCqlzzisdYFGsp/h4qJkXf1LISfaHLL6IFUhE9ifUi
zFUPrmVxf2IGf0d0dqz2mnjDEhfICxCRMsn1R9qiHQ88bYmPubXGFjOxC0ngPASx
Xyi2Ov36Z3CCxwsKtul36GF/x0d3FVrPVfZ70v/9CKreFqnqQQ73pv0Ddv2Lf4Ov
2SpaBrsL68P8NxYNjZAq7d0qliWjOgVSE+OTBpilVh7u81/ttHDFbf7pRx+Uo7ep
4tWv0hZXuIJJtRBYK2LNwT3txJ6WozeKZXH1UXCooqNqH/bssRGc0JbSEu0MwtAB
edOoKZkPCXnsicrA5/elMPuSuapWCbIMgG9eAy04/6tdTRMJSq38wS+akJEJvj8v
yqjotuEO1vBITDtG32X/Tl0NXt8tCfAsnDHfytcP4BjHxsQJ8/ya7JoAdjlHTRRg
+5TFshoru2csotqv702ZAH/aBYUcmUobDy80WMECp/HdunFTnVP2+IsUCPkkG56a
xJ8Nm7WYKV1Xdz9WKsNLYaGZQiOTUU1x0HgO0Q0MB+sx87vim+iV5NxKs//+fJX4
YPQNmefdDxCzc+x8vRjiq23nyYbgj0l8P6W9oFDU3h6xYUY1F07U14PRAmHGJ+nK
9ullZ60XR7HPMNdewd5cYBrbSdUaVH8qAdIpGeh8cDYPNMDqGbzbnboVX8gYjfjF
hJbFy+9Fe0EjjYnwIt5t1bsEzZwe92T+6Hic+zHPzihsxAz/yXJwyyqUqCEXzXLC
ENurnZVwvnPkLTmdEVrL+wzwO9LKH16sInOm7tujCxsThEVFVm3db8axNNqtZr3y
VJw+4cvtHzRzOx6ToiE8rQalDI/p6vqWmNRccBxjqgu8LR2UKbDzdlNQ3psCy/zA
/38oXtOY0dBEoJAF5TwRPqhq52hKYdk86RBhXqwkYebQ/B/8WMf6LIuKz4PsAcmM
in2ouQJ0mUTBFtU/3i1FdFrsUe2Cvnm2wiFvKN+bS17HxQYgNvhbPVw3d9WUsaHU
yuVxxxrYOWyQ76D/WELyUS1BUDzrsl1k6VOp4FZMJv3zuJ8im74Aw24GiDk6sbQx
suKBbw0ISvCtyKD9LX/cEPbDGb0M9M7WPCQSlgjmr0LxDECfDuwsd6IGyZzyWNPf
Inf6bd58XfdOceO0+fQIGlPwjYA5tSDYInxkb6HE5YJ72VHx8r3Prb37ORJttyjl
YuL6tBH0BEY4CdtwbI5mDs37SHBpTaNpmM6ba7SqiuYU3m4Rm7eQXL2X3gWhaRbA
c18CbQRpgQzl/7q6pfJFTmJqKfqMgN9Rx/5uhuncmV0P7l1Xs9Xr1GC2NIdapmvj
CNtIddj67gr8bD3tAll0oXDivhGm/bqstT/M4c9zLfjyL9vTtSShIaNZkMy2CT3c
KclwOi40Q+x73DvDmMKrInATD6koToyNnKsbL1n+e3IKvpRy9dnXqMuRaKd7DXVG
e7N2xVeIQHAu0G0FvGAufBO2TD8ljAZUkEk2ls0n3ftPcWjYWT/KP+kf+gJa+2gt
KIEfEBXnSY6EyFZgnYxSWl4ErhXCLvCOdItTGkyt9CFaBRtgDpUCynbd2f+rfYWq
ThBADL/s98IrcF8DOq4C78goqAvyOGlgOwt+9KXnk4y3Su81ECxsKhsqVUjHClyn
Ik6yrKEoo5LzwdxQ3ImHSbIYqgCXfpo3FIcdiAR/Dc+f9ogBE8Slu8HZhlBedeVQ
BEofHCLDEAxdgKzIL2aUwTUAX2wp4mWJTmD3xFROc0/FLNyZpxOlvl6yU8MPcZSY
4wbkROrHs7s8HVGncZsl15B/xtvv4Z9RgWO/CmIX3TuWXmoEs+lzykWt+kxE97dY
o6MR65O2u1ZKQATTdQ83+O54z3UkwQT4G2jrK9RBwVOsFyx80D/JCNls9ewNyGgf
3aAEMIaNlDy58TiyuCYdwgw3Vml9eKdw2HM+MwZNp+skAq4AdwTSwkLfgCBy0HNE
FlhTrh7qeSWjsvzLNSk40LWAEoa5vHa+xJbwSHWvfeB2KVm4tFzJNEtY4HIBIWdG
0FOvWO4QRbrDzZpdWYSq0NdjYJpOtQPKuj61HqhXTODklBlBBpWomxsIrj8UAzek
JreunlemI91Qo10iH5XNJc7jvbrezydalqofAzPgIHxdlTL8NFALhrlRt9Pdf2Q6
1VftXiaG1ZtwJOYVxx9VEZztjY8YJwIyimBGzZ0Xpql41tk3Ls2gyt8RBldOVp4M
/D06Kgj88H7ffcYhlzeL3djfQXR1XdfmJPpLqNm5kRgiyungFFTpapJ+P9NYVypr
4os5xNher3706YmiYkQg6l63n03vRUXXIhA19bgXzMtnGDHQYQgbHdxK8THzXVWV
fUsdArVhwwRED2udwAmEfKmhk2Cy4ly0frN13KXb/1sEu4uonHGccwClXnnRbyNj
mJU3jrz+QB+LLN6Q5kJM7sceqdjhH1lzllT0IXQjv6EOt/JzTU4i9ZAfNltuoaFR
a8FR5Nbvoqunov9xQSytX8yE4hEB18XWyxuQX4IyBVqpU4iloS8HF2SZHrNSTlVC
NXPC7//9hiF39/4fQmM4eD60/XNDL/ah00Z2p7x3GjVCG856s8a8JKfYzcPS342S
3jYOfzfqczQqe6lPhvub013BtzUBNJYuC+ZtkvYrSmrV9yIz3oNMfseDwFWKbPFP
61tlSgT4fGK8ZuoTv4+yfnJjg7OD9adHsm4Ya4ZCuiKI/Kt0nAMaBZxTIcSPjkQV
wDhzM2LUiKv51ahr2+nUQZdhLVlYsMb6RaBLyToKiCgAEqsv0K6q5M/xKZKg+0a1
tNHSngJQgNVeo+z6TRVqZPmTcZWxQYUje7AKJ+O08DNuo1UF28yNiCYxCWv4FA/1
8MF35lukQMrYRpASUhNUFb4A4SITOy+lA8VMvaVcYy1h+/8BPGfm4+TIXJAryGWV
7V+PEEaa6rdu4p7KI8La22P9um29SM/GJc0GvKW3TxpRQr+Xz2TO7jd6/JHYRV+P
CW3jJnaHn12/56w56OsKe5IH1S2KVIGaIKHRlifGG6rxZZdPAbvWQViWTrE0yQ6/
wtzQJ0y3pnYJv1oCqE39pFNx5HjSzJOc7Uwb/D9gKFjtjfLqTdlknf4/M7zvB28c
rwQ1V0iFOkFg+HMM+Najiu5MyhEMYnNGtSd8LiOIAoXtAJ952vDNTkNE0mwn8Jfq
sKoXJEO7BRvH0zeOpKBdCDKS7U8WVwqJ6st3jVR847Pmg0Mb018wQ0PBORZpl0qC
yVArCk8Wuem/DWzA3d3U71lFjinctyVxVsQ5bojpipkXorCCgF4oJtkJBizHBxgK
4QqLTHVkAA9WxkqP2ZcLiMYbcO2dv3IXJq84aiplX6ZiW5WUOteumHmA1Fg0ya9o
62zBu/y1uc8mWsk7LNaO50sZzrnzTieDl1Kk2EEYW47jj85jx1RvLra30zSL70LD
tOMWL3/15Tn1mwl+EebOVKitTicKJkXPkh/E83nayxJ2UBUwUqKL7I00RxQcQBUG
MxP3WNi85r85T94rpTsHuG2H60lcHXPOz+zL/Fw+SPb7a0xkDd90FnLMpNvEYvgf
jqHE7Bd9fHj0UadPqDu5k1glAIqNPAdTbxokopcSGvPYySP2ZtHXB+OrBwHU8gmL
ANHdiG/kdbmFs2Y6y7rYWYH+PA+WWpFT6FUapc7Pa9zI8xtfUTkiCxddoeFYchFm
PdlqhiVZ1BqfzJaAkktGsIAIMyyZQeeej+5t8T4Q4XFM59G7B6UjzduyxbTmU+Tp
is5OrQl+sfGjEwA6nhu7s6+GKlUbtJAU+Qm4S61m/h0DEnAhxPWjkA9j/tNnqPqB
t5EgNI2zQ39RqOC0NGSiDaEJCGqv2Ve7ABdM06SM5Tr+nbgBf+MBVH734yB9lph9
KqilCFGtrz6HdXKYusML1pBk2E3iCinnQFsmmUqsg/o8CTzcUB4819u3gPySz4GM
mSkR38F8rHrBzTMlaEF+889H3DrbXRwmwPmFIIoTHnIcjH5YH+ylXNOWMAlhgLTm
O3031uvQBmJ9I0bHHUWW9exLcW+4e+TEtNN8JkUkGz/YriSy2vx3pA61zrRerryo
OSzrSotziZHhPQpQS2eAuVjjaHAR88OE5zIY03uHPWFBYrgNpkuQFAZ9HuqGXYIn
6EVe2y3lC6Ix4xU/+L6AtotZu8GuH5IGDj0mB/OefpzjE+A1ujnaWTnU9S5aXHt2
2+9vTIrFFhzTXW6UL36FYEM/NHMm61tywUdJY+TEARmvjuR09EMuZTkrFoqqAjaf
YAr+QRl1uEf6kOGJ2Z1FIY3+8stISlH+3K+CM6rredwDjMSqhUU/pbVcE8B5OQ1G
TxCtuJo13WflF2sax5E66PLyE/5umS7vGOYkHtEORFywqVISCzEr0Gj8Qunt4RjI
geIPTRgNDj39p/q+tAZ70jWCoNq6grd/5VuU7xAQoVqhkC88Pkh6GVd5G4M/CAX3
+eNtTIPhrA8583QuG4nyHjoPU5Zcc9iwVv3LuX1H7mNSojCElualtsXohdrIptga
suK1MNqbE51C5GfHkpQMqCQgnviT2TZVQGYvDwW2yh8T0qXEI6W1lINwvYZb87rh
QmRYjAIJ97zAWkh4/+j65EvbCQvMPeQJj6IJXz8ZJ0ViN6XE5/BSd7Yftmr8fOoc
Ou2gx89LLMVhevHco85rVuuMBPpS2rsfFpUdCNddrDU3VE9TdsN5tBMcB8t5KTJR
AVXaYpzoLH8SYiTdKDe6VMnXmF423pi1J51fOM1WPq0+EWiv5zXtt82xzyrgtHtQ
uGaVE+9WpWRSyoIusns3KtA6G5RYT5SpzbM+Mnf+eF15vBtcrqTLktmQ2zAXrc2f
ZJHHfsARnR0mWVREqpZYTzmsXEr+pWvsmkxsky2xCrhjoRuure/Bau3xYGjj/lWY
aPn+fanbqeaLG70n+mR8675XI0NeV5JYo1hhtjYoqCl0+3yll2yTtT/5oCaA1NHf
+StZZOYNcRDskFSyEamFNcXugM2+PCwqHzTv0ZCJnfPPrybKK7NNZNAA6IjOIf2A
fmpbqGToVjQWGOV1MygSiZCDzkBpNzYsgOHV5gyAseun6Qor+TAL2lDuTeF9tn6L
OsJmAVS2i2/bWARMevDbQ8xssORh3XiV+Scwfm5ErZ/ZfdajqbraPg/o4df49JK2
aQvk06y7Np5ozMt7FiblPZS/bl/VtbRivhYooh3j5YPr4w0HpPf2Kr5Ei4IlDu50
xk8u2LuPFonzdwxJKfCMywwoAHvH42IC7DUdjjgWdZh19j64Pl3ldFjfiLdVb1xW
cjJZw3bswORNflW10W4Utv/yUxuRafGpraFfT58SfxBU3RsN5N/aAjg8K65vQKpF
8F27BoMkIY9B+5l5aP2dKoDjF8ajKDnOO1NI2/V5JozN8jf/yJiUYMfnLR8MlRYy
RohmuHNvm2lnN1geE1dRcdNcN5v/f7wLqr0uVGGUoGYctXITbp1Js2sBtLAsCZ3E
xVML2cn1JHRdL9HABDtJwf+jAjnig4lXo4ag6BtxXqWnRVdOEE6lpBKwRDwXPu5G
gid12eGDwH8fJQlaNBoB6MrO/td4JfIzC5F9GVQrYkI/VvCs/lKLsKqJ/vSOsCkX
ayDUwrsyHL9Yd2zS41CCd9nkl5SLVqP0FekxQZDQV0SQvtI5C6ZQWt7le4XPUiDl
dWjVFv+Sq42nX7iRY5+/JRfpARZMe62qt6qDUConKY/IWENg6ioFU23SqID9QA9Z
n2lpNag2iE6Cst4Ijqre3iY1QXTFGx2lj5Q3WvrEENq0tq35yelu5Ee7JfQ5S81q
x4o1Dltq7KmwC7bsTt6IpNjkOn7Y09hfXDcoojayb7j04MQ8naJlzOAk//pUTacn
2QPUZkS13cMjrKhciOyv1MnJ2TawInm7v8I7mX5R9bgEz4jBmMqhqjCPh6U8p323
DF8pQINsb9s28sOpedbIgl+H/nV14YRhiRwdxrghqIsabREE3MQC6nKYEmOgc5QR
dPQVH1Wq3PI8A0Ywzw38rWdU1k5AXiYwePcBTK+AhGW4wsoLok2FpGov8RILUFGJ
oxyK0mu98c1A7S1jsUOnNIY08Yfuzodl/qZIuxidyIlXNMCJqH7c2V59DJQniglI
NtFKuxVoQfp4Ib+JgJ/9Llppnl7tnzdugjf3vw8vdhGnjuCpuzfsXaoxEId+gepx
i3bEWzjvLJNpm+5lD26mrNeF94ul7w1cuIE6FppBYlBbVJau6Nr231JK6Ns4dzyH
N2R4Kh/qfITklrUG/awmBNC99gvz/ewGeJ0Oy5Gqmy8jz3ypvTCJq+jZbsc+TDhO
ZLyOWzqK0I4WXiwjY1B31nuuWmn3K491ECNABD3cikv11Ggr7meLfCUodwLsdEMR
II6veq5WLA37QP9EQUWuByU6Rvy+Q3k6fDXm0DHf3K00IqejJczfKMFSHcpo6SCJ
7biDdGE2wn10+bl+tGvCi5dnkdlP/kVBPVFWTkV+Vubdu4ZwXCI5JjnixMceVVTy
io3mdgWOUUQyiCQJ8AkiaWKNyIAzxoEOQwM5y/uinCVjEC5Q25nin9t3GQ52Z2X/
H85ORp4WVujf90rCQH3n92D/GPW2uYWF/WzHfmdpR40x6XX5soi+4Ld01juVPf8N
0S1ORu3D+bx77gQLXkVSdL6o9kBy9QHvAOVFxrSHs0L7CqtmSF5FpH677xFjAY7z
sjj7tIScgd46QTnm4FHWBPZKBGH03ubX8x3OXbGBfRewzDI0d83bnK4kZH0gMU8+
xs84OY6raLaTmZNTdSg4uWhbo6a1Kxc7Gz+LHWJiqlYvv9pNEcezUwix6axYfTGI
XxSuBIhJT4g0HpKkEGKlqr6hgoCviI2Gm5tqEoOeTELZnhled2R48I0TWVVccMiR
EemxZySFSO2qN2yida+fLUKmPK+ajJdJlm0nUDRITXgz7TNmPz2xZOlSyCKCMuID
Sb/Dzx7B820De/b2DUfg5zecPqqKB9BJ1ms0kN0KDzwAOmPT081sjCiBEsoi1E7h
+C/Bl5s73nCTcjhoRi5EcFu5GTCG3a3++OAOwbcv6ZUEMUFxcnZvTCK0DcA7mhts
EIz/nBjfMJ1lKRsawRBpjKH3ETaJcfM64UTjRFcKAlMrTj23SWpqZ/4TYWrRmpRW
1IU7WHEo2/MoAxGjzhKaW3hEdgczDlfM6EWLPjtysITAn4RIiOKk+5TkcQv0Td7D
mUNmxgobnwFTlSSxCon9UZoScrR1f3N9HcGxIF4p1QIml8Qo1HBASDMTcKr3PUUa
sK92MZfjK0LWtx+omavP9MN6KCqEWdQ82uN49fuWn5f8kqCLm1eEsUprZ4v+CZoK
mKefERJG7Wgl/o6dobCb+4tR2TXVZQb02jxAXOW9R+uXKzJ/RRkT/C+NlTDG2fc9
FTigqn1kTllSpU6wX1wGgAYhVNj6tC8IqRYUHGugVFWSbTLNL1W99XMTJh77ZEiE
GJ4pAQGaE+m7zXELW4SyxOVWQbVN495BKvM0tQMbPMbc8gLJVG+NLKF3gtRLvXuj
8E1A0wZbodhN8DLGX+0H9BJzemHqWloR0x67Zqy3zMm3+IW+vi/L5QY9Aw2PXopH
2LptCwHEHVZlCETzZ4R6DqD+UowEDSs+AwNvmdkN30u5ymz4UReXmgm1+Dp01wS0
lSCWbF/92MBY1dlWRclUzdM0I+bhXkmjgfgi4MwxCh0ctZRhp/A4TscWEbswYPEW
zdDgO4HgjGxuPTNADCJxcI5B09c2SJz0tdQoq9mvSITQ0LgT9hIID4R1n4XkcPQR
LrprTlb5r+E+v0QD9XmdUoYXb6s9mjgMC1efxfUbPih+pWpqfA6yJOeFEk/rhxjm
mN89LA4HgAvLzwzpc3M/O9M2QC+GG7jFHL2/vk3SiS7/OePP+uYl6A5WsT/Q+e5s
O59a74UGzcw7zmPSnhvu+p/WGGz8JsfXYogaEEiFPVB3wk1I1tPSpMKJ7512P8uG
4wTp/tAV/vITbjZL1qjg8t2bcr+SMEdy0PbblaoVG9Hw3juz6nwhK0YG5/Edv6P6
mQqTbV5MlE4wYgrj408oR+7m2UjsevFVXy61NSP8DU5BGmUgNXAk/8p3FP6/mkt5
IZpAXJv1ONaU5F+jcsYFoqGBfAmwfc9c2WhwqXzT8qZJfIrVO65ltFSALI+EkdAu
YTnYChShFGwxr3LGKbOo4NUhEKUM4oTYYQMg9BmfzXDNfk0wHdeOAK2ejySDJHp4
pPFTfpaiOFZhKv8IgRjv8uRjplnNQd3BU7r9oH6bdqgZSvH6dnR/7JzB7gc+vmUB
hRv6DDlEWsg7s9LK4glFFXhpTwtHxre0JsNrjj30NnT1wGl96HNUJQEAqSo+VHrk
qnEcdmGty8IUwrRpTnbD14NPQsjdBID1cxf3oVRRZJld0t3eAlGWW2EBHVn04SH0
HWo9qa9iG6oNPNAb/y8EyBLS/3yNYs76dcp21hlLDeLakTnDHgAxW5DHxZcla0jD
n161VtM1ls/2HHpDOK4CPJ7dT8nkL17lS13XAaCaUKTSzyUkKkNmvEViF7rDPwiZ
nTWh78ovsPnPJZJHy6OdPM5G9BIgZiyQ7Hc1gYcuZlz7R4tigGB8aRiiiF2JRXiZ
u/EXMSb4NyWdcHXagMlLa8baIEnE0Bi4JwZ2CT6ZzK89LdaSVaoH4iKLJMubXC0m
siHQCUfYGd4Px6+Txj6V0HVjecdGZ0l+zCncZIA46SEjl4GIdkHkIz21PlttmoZB
hl7gGHdgxQrA/EgLfHX80YdF62I+PLaAtyeNwhU08mX9jMMNjzfvu8p4P17n2mOy
B05JDQ6+la8SAHgqjwW3bS4UGTGk6Hz4XuvXOtX3BDtEBKhnGdVmYl1wErkU5akk
1edWH/B3MbeCdBxdqbS3l3HM+eITWCu56FdHNojbA9P0nGtwaFNwHdWhM6gM3Mf3
rf1Dnu1Rd4WGn9Dnd3T/cX0kZPd/gkVTVjy59vxurs9jbYqYdfO0gSJk1J94/WMZ
GESFgYqfxHdKabooCq0H7MYFPxp8w5YlI1FNeUJ0Elzzi6b5GvsM+NG9+MIXwoF1
nJCphjAiQ6UXjOrE0vsY8LUplsBZU1i3dTIRUUWTeEVFyXVVPeyPr2LldN0vaipi
dKEqgA0aYIVyd7gGzsml8XGNsWQCw+B+QpCKhErgQDcq1wkHBGVQ8QKCRhJQ1g4Q
w59Jy0wMh1ZQ4mjpc5JD1TuOEMnNea1cKLWDFvjF2lCspR5mT6wRDLrkso8ovQcB
O9U1ezjOIyzOmpHYAoHZFNtB6bSWLQYw7ubaXqbVbqSzmUPxX+cIk84qdN8Gxexq
bc+j9mb7P72K55C4M1DkJLScQxXhlUl1Bv6wj78gYc5UsKbr3pWEVI84TPPKcwd0
q44HnrGMxf+fIzslMsEIOoEPMC9VaiHDr8XWh1p+Q9wAO3RrE/393rFodkiSR9wp
JaxJK6yGK6m2bhqZxD1RH+XRwWjlXDKGcUwRmo+uVbeueC9K3nsXnIboOxQPi4bd
5QKp8mLoPZFGekcmggmXa6zHGIfgXGZONPu6SoS7YXbVr588hka77vgrh1N7kc40
tKtA+TdofOQXd79Kb4O4u0M/mQdka/uC/C/lTfq9vQLLIwKO5WaHzZyCs0H0YdVy
FxljJ6MSExECG/gTUV4kCn7VRNuVOjPqa9oma2oudfjel6We2c7coJ/Y8GU0t+i0
Rh3d9YFXY1v2fm6AFFizTNnZUrZItuq7KDQXk2Vezs4JK8CD3y7rO981Em+peJQw
HO4pAuRshdA5mfsBFIBhqMwbyPwCKPkv0izCuxOV8RVJs/XxxLp+a5a+26PuRS4x
ohlszzrcKjKWxIdfX/gnmIpuYdgXzqSOJiNfxT36Rzs873yejtmUOMWlXNGU494y
2JT8BuJSTS7rNEdkkEKA/PrXgw4M7bxo5A9gq6dzJSCrR5wTsCpXglJH8JxEZdoG
CI0R1g8tVcAtwzjFoMkx9jujBG4XXhDxOr8KvtmFNf95v6MuG+/xHJsmye7JWw0E
YrHVsrCJPxtqnSeeY6Mh1MxAIRShcd4IdStKlj66JClE+TZ+xnjHwmUGjgudWUwt
4KmX9aWkTGLHzTUjqw4elbvWXItGRkbgQpYh/mYlfmw6R6xAbhjX8g5GPwUt7A5B
DwPzmEaqtl878QEDFPX+9byU0AdiBHeVhPbzDwc4E1mIiWsEb/3KNWxa8pv3ZHSe
9uZ552bFN1hXBXyW3vglGBXXs9HKcDOaW8Gqe8D2CXa9mf11vbOJdHpwTlfexb7Y
D01mMphx8H/nITxxixzCipW56FYWuT8pXQBXoISwLsBRIA+daU/HqIGtM79ayzy5
7uyuh42sx4kj9tpJL5K2qS5uRVIOYjDyVVr9QyO/DfLLQjbYDKHDmWqq7l3w9Dr1
hvBYB/r2liZpVOKnci/a05Xz3lJQWjx4EKn2OMysXkLJ4O6TLHQlb3NZHdPoMCrr
XsKxoijlYrCyDnpCF39MQBVbrhIdunopj1XzXu9+T8Gi13SzVOq0qhXsdiPvjc1u
eSiF2xfFL/6ZzH0Kcs1j2eizG287wRDoDn/mplKy4iDcSUGi5VuepmN14KL1hgHx
10uVQZX0WYRgS8+5aLswy7jhgXaPlpKXishB3Pww9//E0mNBqtF4fypjj8xnBsuZ
endYbOiPBxie23r2igWLdqvI3Gnuh7A1osR5QwO3xtYJv5lmrEpbVQ8KiK8mCQeH
VqmJhw/rJAcXMqh8lvqNyp2Z2rPbjJlH5v/UHZSz0jCB6V63KOw7KfVKh8sNNDsa
3yHwjTKoAOtvIzqQE5I/p9SHUjnUZq3bq0kCP4D4Q+Q46yxNi0zfyonhfa4DGzSl
0qV0WlVU4OIMecSYe1OKuvULkJIgjE9T3YHYSZ1w4zfD4uyfPtsaAfMQHWzKDJNC
gVua0mHgVR/J1PK9cSzKaso7lffqNuL4B5soqrzMe942i9GWJLIHy/qzXXS/1wJH
F4YjWxfUCN8oE6XAp0RC2ce4NMqjpL03+bqg7UpXbc4RR9PqZ3rZ3VQ3lCiJxOHt
9F8FKk23rFDcA+mj+X/wwOqXXK+bFHqZqk186ohL8c9Nwkp1YBzxJ7fdZ2WiVBEx
yqiAYrWeodUI7YQXSgJX9Bk1nczlLvheZhe/2r8SgP1CVFHXeTP8YGcseGnGoWaz
phl9r+FUOkz5/L8I2dnRZHi9P9VtWI3sYFGghfU0R8jYESEdZ0DCn4p0GtOZZkIA
shjjNr98Lblpo8LyTYZ2L0CAZHiRVLgRn9hXgN605keaGBpGLtLD75V+aV+0MHra
VcDBxG0YziTjhbzIwoHFRNjR5fDh/V0CG1WfpDfG59qGVASyoSFC+nOr8VSC3Mo9
gMS1WCO30QkeGM2QqS8diRNd1a9F0ZvTG3sWCTzI1ApaIhzPFsEsMVqjLLuAVkI7
nL/92MjkhjNjjtR2MgDnUulT3UQ9zgyycUoSYgLXbZCGWKmp8de0zemg3kXY9Isn
XWTThway92FeeOtgvp0hjK1S+/Sj+dlZX29kyALYub1WkNINej/z/ydGyqPCAmef
LGi7sherJKXIcng+mKnuS8Lc1XcspaOWCP+XC+azS/YMyWRq51XelfzB74+Xz8sU
scYUTsGiT5vM2234Lnv7zQn9aMCmZHpoUUVrSiAvucRwJ/GvvRIU6FbtGRBtTbVc
QcKhxZeS4+daSWPK4vgFhFh2hUx1JAIuUJAezCYbWESQIvd1yeapW8lnXoCtVVB2
K5gPhNmz0d/g2gDRSkxUXbTpyACDnZJSwAyQ4qwD1iNKqvyw9k+BYIXf8G/ADhTG
H6z297TRmrpNXqPoE4n/FSZ8UhlmXrdVSHFqf+RCqwBRaDkS44AMYpv226sUnSUa
mP2D0wREcDOlPY5u/JhCyqEtEmNHqOf7b13YmxVJ8RlvblobRiBp5ycHNCS1QaqM
YhfAlg7Ik0qHg2Atcss5FIUvvSd4UZcKvxX4qerEWwVpIm/ivuHj1Gq0HCY5d8+2
yboCv2apwUT7sZkX2MHjO6FsgqU4TlZ3xvBqBVj/vHgBkBJfODVjrU4PJrAcoJLo
jsPehH0+J2+D+nsxwUHzCqvLYkREvn42iIN0Cono3LHvG8bBR+NqHvWFSA7/KSO3
+THP3wqRlWcDbFJ8j9dWCSzvxiIvLs+CrIBht8/8FUNwb7ZdBWz+Z9kW1a3qqATn
aG8sEQQdMeNHvPJUYec43Z2s7EiTtpGQtSiX5b3YX0gNRJrwtyUSpct01EiVsaKh
ZPLDmIcZvJh5c/n9HKP42BFrpIpZSYGfTboTDE6ctzPqTNxPypF018PeXr0FDjvq
Y6IVvvwIQREhclgfa2hNjODDmS20+/v9YMo2vmmC8A2B8IsoN+5rRJaC0+FikR7u
PJkK3NXqIAUkivC6LMzIHlNAccOGEW299/4+YiyDfm/ZPl2ew2xbsUt0M59OlhEJ
zNCkT5qcC1KJXWTLNTC/uEAlitygrZ/i+4QN95V5DRdDYRcdYEI3xOIZXZkJT+7d
AYyKc0h52g5f6e6JIedbjTF5Jk57M11Qr2ctEVjF2J8qan3fFA3NbFsbWdkdbIy1
ULa6Y6jhqSZonKqy7J6okM0MySSUyaduEjyD+bbd64b64SqrcDfDJeuNtfh8y52S
AfDN5qdGiLg4YtqBnOhXnjrwnEtbjNaROr+rISOcG14NxjfaveZnXZeghAWFppzc
wC8VgGJl3oI8xu3i3FD4bBQexO9gBgsjPxwdc3UK/iZdcoXzecc6cTN3xRYzOKMd
sBeXHi2/ThBZyfqyjvmdcuhgnUv5kxF4KvPWwOA+nZ5/14PaHB2k/3Ag/Pm/IiV0
XaTkjqRbncP2qKaQlvRpJgk6+gArQuDjj6I1TEP9aXCGQ0x4pYZB88bKcqXklsd0
4KdWNl7aljEqkfLv7ZrJSpURiM66zckD34asVNaYfp/yf1cSR05nfhhgHE4e33rG
qN/QkHOGXWCBvB/tAUkWlMPrkvvqPwXdoWGxlXsPX7Kj3TpRH0Nk7aRQaqGrN/pM
+XrCsHsstFjBHkIVT0sTi7fB/KRB+gX2yrL318Aqi6Hx8DCVjGlS/MzgJq4Bi/TW
TNQ7rFot0NITVo3NfTQHKNG0+vb8Kmci5OZYIgcywQC3XQo15/7JvE+hIgM1LMX9
gpN0PPNFGWxA/OGJfKX3+MRaQ47Ugvcsin7/UawpOGdb4bAFT8fV9JKytkuWVpRu
Aen+tHD8ZbCpA84nV5NG3DQky5bGlL51AC0+9irln8SlxkPn5aVeg9764eSONu/t
2DHYa00errbRRpBZCRuFitEmYn1qYniD95jGgjQCOeadUeurMhqVnzb9hBjsW9cq
0PNwQSd44ZlCYszgzM0XC7Dzc2CUMPuZK4IaXpRGZkfSPpHTW/P4jXB2GHkfT8Gu
PA8G1PP73WHOJGTL2gTpbSgR2qHe7YgsTBPPw2Teyfbix1btTsMGtm+/7rx8XCH3
KLk8ykyORTeWvrE8xMYC+8TeTNdgzob2maxtIZsJ7UhQfxo7UM9oH9EUBY6WUCAZ
TAidPQUAliHMGJOoHYxZfyOwglp90HGF/uZ3cdgkIVMdQy2BJ7BSp3ATai3yG8rG
TK5exeQhQR4Ut0hNwgpM2uollWLcwdiOem5kmZEjHM8JXLZNeoCgB79a2ZrlmFKl
1OKqIhxt6FyeGsguCi+A1QSvPusIV8Q7818A/Ia3zh/oPBVSa/Flkf93f5bYPFBP
u2a5cy6DRaU0kYNTDayY5eghIgrRv1Ml+6nwCenTcBTXegArms+/0zA3QE4sukWw
J9wPnhQppY9TlqJ6NbAaO+5cWQdKLgSmsCwLh3P4uj3/GEZ14+d+ahr6OELmVQkW
votFiTmTzj6nmjcDIpKUMezpLyr17ucGnnZcbNiEQXZs8rhCCdx3BF3c4EPK8KuY
Y2H0d67DdNxChBY3jo9/gEcjY90it1vBxPSQ37l+CzTS1B8ZEkBknhwJxgPZCQ/X
5973t0ChhZtdYw9UdpCL6+LffFdQCpL18oNbGIhRyg183h1Y1vTZ7xa3+MyCJpr7
km+0E/dgjdhDsr8XhYkNUT28/mM9dUh0w/MYb4oG9GfCeZzyj9IijlC9HwAdvToo
L+Pvg7lLtjmxY8JC6GgMz1ANlmlknkvmp6R5me4WXFsZBjF+7OXI2d+ywyz3aodo
BjepT+mEsPf1xeA7K7m50lMW8mW0bvCc5vfXKk6Kmb8G1o6tVan2VTr5d31FBATI
JvnC3wFotNyUA4eFhKV1puYC+jIGISjZClnRqDBhnsDGrCwJg2lx5nW38ZDDLNpf
SptUmDCdW6rtXP4PIxGvQwVUSmjILxi5PLSaX4D73aRbqgft9pemhkrr+uuOI1s9
GUrCJk1qJYN35hDN6rHL3r10pcz8AHpFv8fMjTOHy2vnNKj8WeM3SQcwg4v2M/IC
kcLGOtdThwJo4pvZ2RGykOT7tiwWV00wyhfeoKjUYky7rpvoiqOLc7U/P/lBiBh4
NolZfFHfMrbqfDyw9NMGZbeA0IWGMzRsbDABS0cX4XQ5eieBmLaq1TarhEU4uYX8
twgkMOeNjKuo+iiLh8e7BWmjEQ0tdr4xkQShqwk/vXKJLrHFliUQ9A4cydQ9D/2H
aBthZb969QSL34fGag7WRPIt3Q/vjRRLdiR/UEJJ+OIgu8MGUCQF7sG9NScwp/6z
ie927z7oKcCBscUU+PUJTyZ4ZPxRwOQNbsOgt1uQ/mG88rtJYpmif4JEtDfzrATH
y3ufSIf4rdQrbDRlZ4HHZrR70a7mSBzNXAaMGYaMznifph2sKHBslE9pvJ8iZxqP
m9WR3GQ1WMNQKIc0pthg1h9N0sj1R2xOqNbYGGYodYHsgHCBzlgXDbZrg9cLMV9Q
4s6lbK4CteeBY7Yd5yc3wciNgZCMTApfmbR2z5Sp+Ck8BVUJR0/mw8e9QTJ3UqiW
1sRBT/71Ck95TZ1c656poRkhx4OVTyogt+eqKXHROaIqT/LPcZSVe7yALz6/Zw1O
TRL9VtR+I16VP5pTd0FpLdvpjSra3x1ZIFwTE6Oq0JGNHlXQB7FvCPjDWIBZWgkm
AoDj4q+vXEiyl6ADd1PB9KQQxywxIRJXNuwd5ZJEs63aSLttwOOl82ZZ1jOVXw6K
OOBhAn+JJsXJdLm92aVeIpl0dJMxkIMCI5UgGqlDjEVU7RfHiGvhmdbtVCu5kCs6
bwFZk9cTOh2fhzBVnNEwbnqN3goQUhNJSzzcIcebGW+VOjcl0wCjS9RwWjtHOJQx
cb6uIs3vXxY8c83BFzhv3VBYLhjEjgVFHypHhFLhjVvQ5j4I6w+oDHa5liXY7eSb
ID+Q1Kf73nH0nQctP76ynDRXqrF1j7J5uKJIdjVuKkeGEW6VdKMfWg8zPL/MEB1w
V3DMwehEHzG3SDRYab86nUHIpLuswXjuDEZgIcNJE5wqCXOlzjROUOVXJSV7UPtM
RTcjIbJtDRYdkxiA3DrWAsCxmWiMR60v6AcltPOHX/Bigj4cD6/hSWzQR5vu7uEv
wT5u3ziSboPy7LTnp07cBa4nG63/YQAsj8hzrkpCFi2Il0xOZ+jFhH3ZNrTb5NAM
PPyppFt+qH3ZHwc0HhJKHIqGT9U2/uQZXyv9UXQnR/YdX1ruz7ZdBbFVx8wc5E47
GR1D4XrLH0AFFoYoCgZ16QZi92c7assoelW30i1kA6oJxRc1upW50V7YGJLLku6w
sO2n8ggIESW/+cmYg8ryvfK58Qspyp8tIwc4XIFF+9w27l608e0PGIANzC2sSTqi
de75YKSkj8YQL1cdqVcRJBxKeGA4z0Cqg15W7V0RiPbV8wMXsHKge0BDXhmFfPzQ
Vp/DxkoPOlexKhQ9iFSjJoPzmfQ8Of2XGA19kc08DydWQIHVetZKBLWmChcG+E2S
E6u17tqDhpAyqP5gLougXZOPESs7gGYAYShxZQ+SLyWQPPGQha47Ai0PVfu32vmW
ZohsoE6iY6+LESkCw7Pv/fR+GdIgv4bBGgk+1N+n2Fl3YnpdLpyAmZEAShujAHD+
QHGZOCBuiL5jSqcPcTPSbDnu3QcYFIlXHtoNhexjd9kiUCqvbGxZLWBZMP6BlXdT
WteZijndFJ2VQG3snEEZHrAkuDNq02u3NvsvBVJWZGZ+RWwRSUMZsXBYJx/U0qsM
urDA+tHp2RuG+EGq3xKt2T1vXymXJi6wZR7UJ1WUHOF0tUKbiTLoipG4LFG1eQiI
wieXEuS0eVzKuNqwrF/Imd6JjFg4fRsbqxvFUNQPp9UCgTHd4+DXYyBVqvW/ddf1
1Ab8gLpfi08flBPl3x9uCyEB7EIDGQl/+DBczuW6hMgNLKJzvzaCSEDotoTxEVuP
f2TyB8dvTYBepvdqt3KCE7KCHs7SjEN7jegQweGqH+Pes6Y80jOAlTVNzOEsXwYn
eRh9HHvCfVaqwpP5wM/6CPfOBasiaCkX9vXuQ6wn7pFhTNQVaxfoQLzi5s3qdlZ/
oa0gRtj0ooWhom3R+Ub8YG9kc2fCzHn9qhuz5bxRqGn5ioqTz5zLnCxBWvsUUFHL
EHkjtjU/pEoVH8WVX1m7EPOddcsLMbUop59U5xYcmvqF20qDrdnPiSTN7pWf/qCe
yDCX07HF//rVh3UtZKwE1Wi0VjTZ+IjLFIASBawMvxvK1hV+HXC3PhZBX/ySdj4K
P/R5pwDx1qj6HXIc0MglwfrYbyPJThZv3+aq+HND7KVHb22H4oW4xbwt7fdZgElO
Qdxwl1t8BWE7r/RrXFRW8taXd/wIz5Pu4mhzl0tZ4p8LlKxl124eSHT4fTDENqHb
X0HMUgy4H3ecaw/6VC8OOUsr1G8te/bs8BeMwdMWPspyrHmQeDKR3RT4A0vf/0Oo
UO9u1KWFU6+seawL7uIV4itSCZTQnvebJF+4owGCrP3psQ/f0TR3XwKuEHaem4pJ
/A6MT1ejMix/BJYLszVh55AetBDs+kwDvsS+hvagp0mJh8zbEJVTPh6hpY7PKSRz
NloGmt1Jq6K+KbdDQ6a+S/gkOLcqSyF54ehOQCc6rOdh//9uHSRw4z4gCRPtPxY6
3NBwgmsE19Grn1IvWsI0RkPJ+sq1oWo22twPxbzu62fx6niApa6AcBs0xNf1fi3q
Nmw+P+1Id9p7S1e2dHcaHkM9Zzjj/k1GMg5pcG80J0DTgIBvRxqNpOxZHG21pBL8
ZOY+9j7QW5cx8Qfsd7MMCKQ8BsxOmqhHtWFFHeF2oyEboUUSQSOCDxKzKrf25cPc
apXNseDnFk60u7VRE9RQ1hcm5KFNM46ek8coi0FUL6aehyENF+c6JVT6xWEcfxe9
3d+PHuzaRgezxBfEGXxDNR0bF1yihpNs/RLejtG3C3PnookkZ94bGtPNbqvrL5mC
xoVIDmvxfW5JE8ToZ/hSO81Y0DWzFuJX1rUVmt220MYPBCTQm+gAXBFpfimX2YnN
LldhZxOCCNJEvl+nLDjJIBTnvIib8Tw0B+lpVsC6axu/4k1lrf9XOc3D9ByqZ3YF
MYHmEfddomZu1p/seGvWk9Naz2CmZGVau8CUE1x2CepQf7qU0D7cSbXaxiTes76q
Ri9C4S8ZUsgd3sdARUS7b1gr4qsMra+tz7d8oSXOmumqDj75e8JkQbEKIcMGghHt
nBNrr0gkPHNgTv2tvytM+4zqzdLdbZy/7NCin/wErtk9+8xcWtbxfoCHjIF7McQI
/or39qstq5ATvhvvnttx/w45ZwrzUU85Ifjv6i1ftJkYEcp4PgR7ABEqz9XCzcc3
UntrCKAZ3TaRRG+hYFOZh4nnzlt6fBxZcJ2OxFndGm8jvqo7/F+J5hIWgAs0CrmC
kg1CJYOIHELxMNvXZ+eHZqYnyz7ovVrBbFCT9Op8Vp2k+jzw5v7VNmrCWicaSUYn
O0ODVV52j4XIN/sxoKak16t2JQtlcLWmqH3qHi1rjGsFsLa8fYXZRRq3SacGvbFK
f14cj6JWHF+iUJpeAP/MOTW1SkMOkSg0POGPNYqI/gW4+JnUg4Mbj6R9xCvjwsww
vhJxcQEpnfr2fFfqaEYK1k/OogBGj9stOlh8QA8Vvveq+8rRV78nzThPOjHUmVdJ
Q3QQPstQC6g8xf/X+PUevTrd+UE1VWSK0EFXBpCZdWMgUhX15ycKHjaU/sXzB+H8
F4mxnJVRqng0qy9hGbrSF5kUsDI89JR/7vGOEltOdYPEAEw14K/q0ZaHQLP3k3vG
hQbobL6WGg0HL9N8CYeZJ+EQtd0E+LixCbhkoAYSUUHckkrarDPKAK9i4RRtLwbq
X6RD+4HVOsAiX9ZW3x8luZhpBqncYBbg6uJiR9SPqjOcvtZG4eSQXB+EMFNMT95i
EK3DspK3xm6U36AwHAxToKl1hfUqLY8Fdt/JfhW6Lwx/6wq4Ihdq0gxk0Snabi/o
fRHueSBJzoyhgykohEhs5roW/kqve0Vx+x6gmrBBmmu7BMKdhPgSJczrEU/eQJaO
qfK4YC+BNZU8KssG/GnOBl9UBRh/dgHclTSmm+z7oKudbUvMuiABpsg/OUdzCzj+
fIU/01jJUdE9boqX23SFKHy4pe3vE8JXHblmj2S6DMtspsltr2gYEXkUTltnB7oX
wzXUtkFSRKJ9K7+LATghzD9TrdJHdf+LgzNTpFu3JirS6d3B9aAG+AJWpKQrBo8d
pZt8oYdOEDTbc6uCixQOPdIKd/X/0NuemZJzcpOtjnD0RRXj8IHmLZ7l156PLyID
h6WoNbhBE46Uhx7n6tuRWFLUFUwNSllaXBolm/ADy7OLps/icu62L11YJjyPo4/L
eRMx7lufEeU5OzzfRlmlIhvqd2CN9+/jsXjhB8RdA2DPkux4YFFeyhqBSX6ESjyc
GKeUOW3KIwa/7eOdtn+6AQXpXU95E3Zl30osGEPIY8G0FLmZ5OVQI8CE7qGMQJOr
XIGs2o9C1Hax29q6z7hOn98Sqhv6/a8+u7iNJD2vRELJ3Y5r/OpLjoK0UBSVfvXS
H4WP4+NeqVDTavusxBEEYrTuPeacWiqcsBy4ZhJGqDsuyIgyuTN5b99nMnFC/s9H
YfkQOt2nIKFXINNLOua7IYA9TKaQ0w+Rjj9s5AQky3b+qsQAaM74mmdC1HDWDPRL
jFMExZE7WZMYSUfjFWlrN+YNjATZIsBN+PxccAOy5dYvBVnANMts9K3QrQBu9ADQ
eS8Ygfom7jHBSNsBXqdHlvmHXUrBeC1XsIk7cvUhtq4pz9lxCBSZPSVs6ktrAeK4
NPHaGBAhpw9xoVtgb9nhhW5AwyG2tAkZfwrvJL5ka4X8RDUV10tARTsoI+35p3TX
NUG6siGNXRMTLhRTS5mP5oqkuiuyhIlZpUnWgVPGlb1YO0U4iR++QaxPgbgivHKD
Bu87TJ+KLhQjA0ZmhNKBdr7JgjFS9kqxT64iB+Q3SiBSwjWj0udfFiHUtvxuty8x
UJ+fBwi/wN1rR7aUwTlUnUwIKqhdqpyFgQep/EDW6DTEyPkrPbgc1EYAWb8prxuc
iAeQtO68xh+qhKKunBcGzD+QE827MN1AYAijoEAUxN4BS1DOqJgRYsIOJfUv0SvB
VFB68Z0ACobM4UnDFLWRAxZFdeZC5VvxRMlPFcoHkUF5wqBReopA53Pi93MuzsAF
kswByIGZ5HSFlEYBYhLYvR+Q8EoBS672sP4LZRCBFW/ZLdXDPuhEdMABdWuvhm2O
Ugf+3Dz5ga5fthzflcP9ttrRIIXim0rhulhI1LjSxBk2Yp6yjhP5VvQ6yOJyoRIe
nck4th4gCePZZMkoiZmiJPdFBJMrJqYpcJdmB/R2AQmmZHTA1lMPlS3U+xOo6Lky
HL9AL0Bjl6mUHeDR+nlLDdoBlyRladjLOV2XNj2k23rJAojDtt3jIQizE2e0e61x
1qwnEuGBnwRidx7Rs5FnxA8wAJdqT8u8aehVKdQ7Hqx9LD2WbQpRq0S3tnMzsyAv
MLKuVu2OBp9WqgpKYWH5KxnsXyOl5+amxzobbaRTp8eXQ0ZOqMLBJc5u0P6Dsz7S
ALk5Algll9rNBGcGBfxZot8VnYqCudt1zmZX9GcnwtOU3Gl4iAhTYPzYWg3tZHFl
hGCvlZjCYtHdziYB0YMxxoTYhhIXFl+oS9+7XSQZOWCqiIYRNt/lzyM/oykN19Kq
E6SFi6g5l68kwFLoMWg2J5pvqpqPdevlbm2LbSNzxG48QZYPaxT5DBP6xvUx+7XG
JVcm3WHGkJAbFiTJj732VA9MVK0CTzaqbX6LS5ifAKo+BVtijgWh7sRf3LR3yBEK
SY5EyCFRpP8Df2hrHBquB8zrrP9NlO1GsmhfkOLXLfXHCbljvD24ESdYywS1cyox
z3M+13y8i0VyNslJQJwZ1/I9NK54VIaOYqKihdQ5Ceipwmw1pA/NzBWEdwM7vPYv
drxDOiweTOYOM8i2RS6/2nkkNfDGxkuDOL9TObYcaBuH2tBCTW8oELXGUN8/TTRL
MB6rtDhIKAPL2uszwLg7VIVEKVamYp42wNoorBqBRSd5sDSjnxz/0W16ozgrZqNZ
0zoVG/zDELWMzbiiUdPOJaHpbDSW0GFKOGdewfW7MqGfdC6VowZNXRzlsRul8UwF
ep9qw2txZKV8iCKdTDPANzk1aR/DhzNIzNLUAt4eKQVR8wrg5gSVVn2Gp6EHHBnq
v5IhRb0X6dZjMnTP+uyAMxn9Ps+ex+omR5qWxOICCkLz/rbN+2Uemelto6Brsa7J
rYEIELS7yDnvxScKMzXzei5rw0AulPOFtINiAIkH/E4ZJyVTngr4yg+NruZCyzq+
f/FY4YQYgcjvvoPQ3rRNB0O3x8hVGpF/QTWfBhSchfe98OUi4a95ngBMeYUHLhVj
M5OXHCyOIbAZ4FPKXxkFtt2rNZY8N6CEnONDLi5Swxw2cFb4I+QLX3wd4xpDtzPt
Py7tc9//Wg3VZSQTbp74bCKrU6Rs4LbGFvfgLW5HgrrmUDQzroEKhmlKiBIyco1r
bi3dfXyBtTYoNluKpX5WscxBl/MidJrBiBc6t0tInR9+VSrITtDD0kKyIqfX7NcU
o+VNUZMYAFSedCCgALZmiHVb+Qn5ZRFk4VOWFU+lsFcUZWAuRHsZ9CJGmfqZtQHG
+18tjox44da6j+JvdI17inAjC2KUHVbWwhvLCYvgqbjJg+rsDZ6Wv11fbb4NL5/Q
JPII6nxW4FclNcaLQw5PX03a24yXyEsE9W4mG0cCFWTQggjS78U4/MxDoiCVSsO0
I81B95Re6h/aQfvhkoD2BXro9BTloUt3uShDj3OWHlCFdmMHXLlDPC3JUVoSi9Cx
jeoWzdN9RuJYLKLojt/bimmz+C78sQfEkf8euGKTP/17XSXKkig9QiUbMxOc7kDA
23hN0VxqIk+2dKNypWDXbkUAjYX/0GfjBKfBkgpvC8nZVx2dH73pJGDVy5jbhMFQ
fEDgQ1qQma8orhhp0pq9nf0VZN6FnI1x0886Sn0sRhXAcjjd52/Jlf5uPg0c1jMO
UyOVOg+RdKzYkI+3iNBmlfqYjZlkgXnfLjQQCW+30rySPg07DK5bMyyRVLUPM2N9
ikp5ZXvFozUy71PmaaHyVRvSkKUxAYPZGLzmTfPdy9V1FDXhqPooRYQYw0NC+/ho
vpmC53lDO3Wjai3kaH612iURenecQ0u/3ZILpBYFFQVv0Fzd1Kne5Ajj0UfDhTHj
ABrPqj3v7ale9J0mtWz4ulf4+5RLhHpJDcahcHdnrlHYWlBIEE1uCraFBLTImGQP
MuA4WGXyJPFDvNaryxpGMwFtfdDtcrepXInZbZaB+UBVxBkuJBY9TdKili4+hi17
x4tkL9Ccvz/NT+AsfMicW1DwXYAKIgjFyRIcRf+8m+hmSL4rcqc1kBS0/AQ0w+Vg
bxcdwRcF41q/SBdI/Ef/r1bZcZkSMuqWWgLW9d9IGC1gZfZhUKgya3s5qx5XVXny
D5AZVQp3l0fsBA1Su2+kM7F9tDMwYAbW5fgHREfIW7x4VBwzc7tAUVu56RmEKzpr
QxKqr38x8u1Ah1062umrdxQA3KoMBre/U50VjlOtyppGGziodpfdynWfyt5RoXE3
VOSbvvihPSbkYlkL354wnwuwITB6EQjc82gPLMneApnNw+1VBmDPINPQajpNQ72P
Ta0t05B0q+vNDTmYGb+nSMK1vgM0UEIsYJ6tHWNfrNaJxnm0/PxEDy9ec2nnKO1p
p6td7lJ4CRf29voCpl2+SacRdY5jjV+MhYrzDhEeIL3iwJoWmDl3oxKRCqvDIMj7
hUEZ/Kvj+cH41otR94Kjes401UM4qp+kXEOts7D1onclM1n8/HkpEXiGgImhAP/B
Ym4NBLrBJzRnEVWSVVsnY9DXOTfpPCG3jIa9t5mkuYvQjmC1qtrbw62vQGV0j8ZR
CgY2pgRtPVfvL64nEgWwRu3RvOOHJfjgwxfoCorh8RhOc7e2oFATpgZtMkIIkMmG
VbEps6/lpCefp1aouw22seoeoeXyMUIYPQk2qQGfR+3XRws8KPpdgFoxtUrSdBg4
DgRoyLaDvfnw7r2WcmfHZI1ZLJdrEuXZ2x7B8SCp3VUPjwANjNbLU5MJbme7jDHM
pcncSWxgnDsfT3pl0KOoBFvPiHa8qQWNzYjtQ2kTxIzFxgZ82KRUEElyAOpF4vN4
t0Kms7whmtWgeS6lDAe4NzgQhKsFl7xor0JAiAW8ABMJnymmv5jQbOssxph4ABc7
D0UdZnlNGpbu/Lcnu8SIUhLRddkbN1N/Xl9Y6OtLaGbcWGb+zES8gASIsEIk9XHj
DlkbWzyhxQtotQ20dXLBW/q9k1wWsg+7tLb310+AK/i1JKlSjuL1eYSUlGF0qrV+
7S2UrTNfkKcqVyanzgtFNmyf5MxQyEr77+mAm/BpFUFfnvvnspKtDhKyjYmjpmyq
AIo8F3W0p4G3Ok7Dq0XDg7+zxtMFLyCoU00jb62WA6z/0xNlIj3hyLlLDYotNKiK
8ZPKJ9VsFdt7Mkihoe+bKxNmyKm8V7yT++jd5+okTyxFu13qOjqmxxb59Uk2cRUh
I+rAaKDyR4+N6ysBerZ2ZwtQAgbgFXPDckqI0qnJeVRyI7S+FPMuySl27jJUPCvW
D0CmTEXo3FmVUf3liMCjfG5W+w7fcB3w5cf9q2bm8nk06YkD/ndNh7K9Njnrg4tI
cqGBOG73PcUt4jn4qeFxrPTc1BpoHWd+6ItIPUPyH/OIRfMiOsdG4HMYp5xRg+0t
OjTu+xhQpp1flM21wXFURK8QE1aUEIZJ3fxntLEXGlUmZrgYdPhMNcDTx+BOAtGn
ibwkjd9Ke81V4shLvS9p1Y6pdaOlhAUUozlAkV0rBM7iEUybdimoQDbIioQIi4Du
IXwJXEbrW8Y/kcK4gf6QBmclrq15DBkTCo/EU6Y01Oeuzyn+RQy/NivQccDHPZZ6
chTJCXqGp8Hdq+eh6S8LV8kKJIBFIIYoVboc9QblWPRoe+ReDJOJaf5fgnvdNzeK
kYUdKsDn/hQFeRXGF4TseRPUhPhXmsyke+Tunw/7vAP9JE8M9SiZ+SGjLN39MuWs
INGP4Sfmo5SFxCCOKwKpz54DaMEcxM7E2jBW3HOdUvBf6MsJCqCEj6cw55h5eLlN
YfZeWd3Le64qPyFmz4dMyckHJexzyoaoL3Zb7Es/B5fg0/8Kstqj4trsPTjrzEqM
t4V5xzFmbb3Zyb/LOD0M8MJnocdnkzSLcbEIsEf+g1MB+MbRF4TwNO+t8j5cR5WE
DIZWTuwMghkrng7vmiVfEQC+tqj79ASQth/fpF8rN4PPBPvxFEQAtk/Vqz6A2wxs
SaSUcJYexNryNEye+SAmUXxQ23QTpg8thQ/hjFvJPBc6I35nv1IyUNJUQGYTUEBC
ocyhFf9j/q7S718/ikkUfcszUoMGYqqO8g9Iwmb6jDQTGQ1+pLek/cOCbWrNZV7J
vwY+KjxL+BtGCteWlhcZ8Ew7nTu2S6N1uQog0VUcNLFENz7URUagjH4p0vtEPzLg
umFr381VijM+2K6OKDbprxmzNcU2OjDNKKIiMZD3gHeDpx4yc/tB9P67GKDo8269
bgPLgI53RiFdCCxuyOplBkeKwtNvDdVZ9lW3rAjDd2elzplqqFXBMqrpTnCGFsTT
hcVK30vIgAT54qcxJfbpjM4pEBiPZinneJL5cVBx+mzoFbVi7MpkTfvEAy8uyUP1
6VmdtsqILDmL4pV9IUukGZRcrtqBEf0Vs4thGS7x/vANdL7Bbv6PcF1nulMOz6l5
QVlvJrbopRuf9mxhd68jYhT43W2qknsksWXUWxH/jiI4XGhtw8jqFNQvhHfiiuZ8
QgGUB0zAGZ2bc4xXxoObKgJebwNkWLiMNIrbIIu93BkJQeBGW6j7juVFviSvChJA
aeS07Xk47r0gzD1zl2GR4w1HZ0Q32fk8Pk9qlSiyIaYOhcYt4FdnNi/2dp26zgil
jl5qQsJQtWUnuPEHtpY0P6BO6bm+oapWRdz6DTXGajRK/afznkf/+3qqrnyGfs3s
G93fnvymuYF+G39vr5QubMoZfkugshI4pAQ7cjW3AU4VHEByWF/CgVGf1FywIbyF
IVJTsA4N/qyGehd/RPVXYVZAN2NFD0UrgUdVBY281bjOaqcAxgLLQfBC7nks9pIF
SKUEhTo7YKB+dDuQgW4QncNjvnwOcBpSvI8hPcu9DOVkd+v0DFFA76XmA9jDiYc0
spWFwYhMpH6n87aSoQk7wa+GnHZuy/2KmrlOlB/CuRGrd2xi3I8tNGIngIP2DGcQ
IJc+FYeZNqz0qbgvGUMENAEuI9qwDexObgk8k15SqicZsbXOT2DEEctT9yFSTohb
eZttYadZIX9Xs7NIlKyFex+EAfv4mEYCHT+69NeU/nEBsxe4gob7ePE7TxeBdK6d
5i2rWbQl2CBQCtbijFGuLMRmfreEsUicHCO4MwcK+LcdhqqZSCgwpQdwS2OHJHPr
pac14fXcScamMzubZzmRuTbFOQ2X3V3KyzNlIOb0iwf67DQfukpPSXXnwuTYuIyb
z28Vdc+66LMfUq0aBiwRepSwr/rTrREWo/ynyklue/jea12zpw9NMt+KSrJY0WNb
rRbIgo/N5pbCry4M6YKGemuFXsdg8YMT0hl4OpfuQJX6zQUCy8Xd3OSyDQca41tr
ySu7u4CGtG+mqYbrXpph6sPl4blPIOQnlvSbdLipjC/IlnjJtHA7EaLVICrlu33U
BhzkcX1Dyuu7+cz+S77iVAfNHRJx1WdTgRquTAK3b15X2flc6vbwt7Mr/DXn1tl0
fUL50xby4hd2GqswvTfLareWdhy7aFtoLQXFNDypdaejBaQ6aTsmdZQPq70ZxJus
D7k28lRs03Udbp6S/q89Tk/nVkrKCZGkgUCK4Sv92jOV0TU+TsqY21atdsf0k1O5
Vk5zMZAfd4Zr2fBYH69BCqRU0Dc2spEs/PKUkuTLfMdX41u4Yo8pRMsEZLnm5YPD
0F73GUTztA0Uwwe++c3VzBmGFMlYjhNKmKDDzDYah67/DOizI3Y6F0FkuZqdTXil
REzcTGcivsZ7dHFJoGP8BlyXrQfgF88jEZAxihYu2rQ4hz88IDmyuYS2f2My0iKF
vycxGsZxI7iP8ntWsa/pOs6HqltHnT/XFyg3RB5S0LtC0KApyAMVXx0/eHAjZp4u
KmVrTd4c3cF0YnCHVbo/T+rP2sEBJwF77+Rbtr67hluRe4Hd27In+B0ZhOVCtz8e
0fXIzw6vYNVnjz2OxlLf46k53TCyzBMMjMUXBIGYwNsDlPjwEJZ6OUdAU2wuGX8o
86TMfby4xH611aHE1zZKXM4Zoml82rpBczR0Dl1J25LkRr4NJ3zzHtegIH/SNuL/
RSVCZ1JgclaJ/dAflIiRz+S+PdJisnG5eN0gu0+LoiyHaMvZNW07ryy2cCU119qM
lbpjda7sIENKCeClkUnTj2TvX/SO2BslUco1FN4QfimLIowXn3ZLdp9g3Knvs61y
T+t6cTShPe52JiZX7ujQgkaOzxXkiGjQ6J/VvX7hmIT7ShCfk1Nl3bd3o2nKyaMB
Bfh11fcAax81fUz0oRwFbTbzmrV7OTDhc0nN25hzqLcKpYV/UTaU0z2miWT486NB
qJPgrIWug5HxkuUYb4LNY4btzUQoqkvTHUl0exUCY92mjfHG5K9jGevU5hs+nSxr
bBu8TOhNCkZeNhgW+Q2TbqCldJcStRnkpiyzCYwIjqkQg1WybFpJJvuDs25LH/tS
QmLCyVH/QxrapFX/P5M4kSDS8yo0RtLYwNtXHnK4YHGhSiOVtit1TH8PpSawVdRZ
nlr6JkZZUXjMqf1ni5y3ZIN9ktWBfBjgkrLMe1ZbeWcvCJRyDMm9fC095FhB/zSt
9Y8pBgvpEHoAmcpl6qHVFsPXIa9lHN2sYAGTHspdhNElWI/i6XJKURn6VUFvyGsw
7tpOGsl5kNo+Bds8wAgYzg01irkyROaRO+e6QWuUvIVclSqYQJJ9ZhmsO30iAbeU
NxrkdCw2OOqZM+TuFPgIiWPpbjOeL5D2AwL/io6hMEGH8ikHPdhqXocq15FokowU
eVxR8y1D8ACB/Yz+IvxAow3LFRQ6ydfI4RcS2mQZ5BqslOmSlO4bFTRBpYCB6aet
tuY6lYnoBitKfdSJJ8mnF1j5zuGh5cuhXqFFm3XRW24VLidWI8S+52i4SVaqapAy
KbNc/rHNMB3De8kYY6JQ7MXX39ChUf4N8h1pegoZgih4ql/f572K8SuUxkXZ4ws5
grV7EKwmOzT7ULuRCdaf4ftIsTMhJSlhMcsCHesKHeDu9iXdvKbo0AO02gDbzmop
fO7tk7vvZFhu+qrmOapz9d0TwMNKEaWaft7Iy5k+I7S7M/pEe7c98/ot1AdJqy0k
VreIW7nfEMsEwUvXUG/aoHDVifZkep1ekYwWcEpppVUNvhohcf8YL4rdOE1Q+eHr
zOp4ERnOP39McF0063LIXxle75bET/rwHCT2m2JZteQKme6U/LWA55fnsRUGr/h3
9bZCxMSsq/Nm55SsSYnDQgF4v5VyHb+nsLO5dRh49VGscr3SdJukjajWuDxQYody
QDDNwpfN5/GOsUgwoXXfRrPRJ7Sd/UjDqqcTD3hWxmb/xFOU3Tid63lh89UjBh3O
byxJPaGw3D++tV7ETf76lGWR1zkae7NBflvd8SJxU7kzG/OYI3NUxTf71mA5okGN
vsossLzp6iw1uXJjBhmLHLLdQZetAj1gT7jHnoKRx8SeVNJscd1/1FtIsd3xYjcw
i7iBSsnvHiZJ3S0jFzgOxQMXKZU5t+DlR1XHy25ZfQdwuVkxyQrIIIbGNMJrSYrb
LCJ/dwhK/Hd/nIxsr74OQ3ltSAypzMI3l8U1Vo2QEkim/yNGtWNpufcdJ2jRgOoS
q40UlEo1oJKX065JOe4m++i0SslXxkd5G1YvzUdZZpPDa+XgN+huWDJYL92S2MD9
EcsvZcXYebYQf2zNxkB14Q8NM+MrA7PxW5EpZu5sM8+rEtTnEq7lnFXXif1Dnu3d
opUsA9mzrJmp2kwafExh/UN8DvsDiYGZaP3OIhIvz6tzW21JuRi/YJP+AKFW9v6l
KiNrHe3vIQfk0NCTq8Z8FTP+ePZkmZPh71qx4bBFZgqkoPoAfaQMs5kzxI0wRZxO
IEKx7iN5/BXBsKmOJLP3/savYK3KRlbFDILtP3w6wGmgmmARQUoLfOtRc3laOl8o
KV7ueCT49aTke2r8P7uoxVwm5fxOgfKSuJe4k23BBlxs/K8nswN6/k6QWaPs0Pdx
O3YM95WYAkakcDDxK8WskiyNzTHFolG3cFiLEXXpLxpmepN+X5XXaFvVzpfRdYVG
sG5tW/ECEW3+btKzFCWUcac5xExJzdDQ1I9ZmEXu0mTs0aM1CVGJQKfQER7n77iK
SSN11Rrna+559BxUoA8kGoj7mRv49wkRyOmV0ONvngE6xs/EkouuMpdpgqAYoekY
FxKtgUNuRZtTEQlhSFG1WPIYW5HLF1SIVvdOtpDx0VqlTBbxrkRRNnufiozttB6n
yLszwqHC1gXeSSX2jn3Is021S9uwDh4s1WE3aVzeIBhE2Nr9mb8YWq95mcnLtQyv
5/CdjF0gqNsZEzZNHJ9RPm/2UhoZGSBys09XxeDtzwo6CqrY+5X92AWKZGw26wbk
Om2RhNHMcDYdoijoBAqZbpY1Y37ss/DOxgknaXvVuywKYsgCanwwdxGytyd2yGqd
+Asf9sGzW2Uz0m4WF3TAAkJtWelwxW7jH7geKG3+z/2CjDFIFWaFvzc+1gBP8+2H
lq3e3dxo9TayZhJsNKqcj5yjq0Y9YW9jn0Ir8+cz8XOJSO+flqdw2HDGTc1YGXCX
GwoXFU5LygRYxXnbm8dMFUvZWBur7zkQviWsB1r24U1I8dNWidZ4SQN47b3Rt/Aj
QgdNTKbTm3F6/Lw/XSaJAMkBIBAnK+UnpLAPVhKzNhjAtsQV0KsSwpZ+ParL5poz
2GcLMEcVOPMb9XgJppgsQKDq6+gXDNMkAxDKooEm2Q761U1GrqUh8SPt3r1a1wj4
GmWY3en0xyz8A3BixbdbSAck83yZO0HY6XejdKgDoLfwFA+a4PoytCjGI+tqPQ7O
tT7A8hWNqR9lKELTi6XZgXcK0MzKTVmtwrI2vZJgnfKOaec+zZbJvGrdv8CCPDn9
EhfU1xWxD0DWSg0pS2qkwIYbm5XGNNqwUcvbIRxRjHV7fDsfagt/onLFmmoQWScR
Iom97rmDraPSRaflew418S4j0JDXm4ca5UkYeRdqePjgqD0U3LJHptKqv7Z5Ftxh
M5IUyo8vVZM/FrV6OZUe53nFLL/IskbphftQq+NRJgfm3somb0lakpjr0q37rwFR
A2pOero4LqKSKQeaY+0q8NcUb0HF68WR60hA082FoLT0/JKMeqqIZbmqID1eMtun
I+dyJ/paMlkqAWLAY3cym0GFwqe8DwbSmyK0V2YAB3eDdMM9CjWLqnhop2EylOm8
sSvDz173KZ0JaRW6iXjVk4GRTYpxA9U1wBDt4WxrNX8xoy1iHP8Qa87pysLsRQig
Tz8Ix+yJeSlU+Hl6zMfCxKbphMxTzVoCFmGsclDZQfSlsQQdfdIgDEYBaDDn7BVN
K1LhU5rU6H1zbb5dVj1el609fSC6cbu38xP+l8/UFssfq2HNu+stAeI0MMgHYvcX
bsOpzs3JgiPYh41tzVAfDXN/JFcAJWQmOSwMZ5Fp8OP0hh5USaUMaL/D82mrHBuB
vLabtg6rvbSUkmTjCdIvp8KC8axophzZXeUzz1XwcVo1IBFUDX3O2U/+Hbaa0Jw7
cK9X5eXUXlciWe7WE7DGxR/2TIkoxkNQ7rjh5s8f23KMzMpkUHKTwJREacFBeWCu
UKgugHhHSogK4u1N4O19mDNyZfBJvVRDPshTMPQdZ2auWWWjWKkGFP1Lb3weMmcd
R03rI4b35fD0dB24io81wgTuB08GAlUwR659mpmqOnQEHt7OsLWXcUtKnPqbUXUu
Tx2w2v0QRKvLsOyE5ycWm1EGhlLL0qzJqo+M/lewLmex8ZgvlFyh5/BMmcs53a28
1HCgxDSqTUWE3LQGkyb2IwgMKpWM0CHYERcbM8fPzbTP+WuFNmGOy/PiwoY1uR86
cbD6/w+rlGMZSxe/Y0ROWzbFG46lwyXdHTduv2l4TvzQLW4Jg4zwk5Vyj/FFCQGh
JfAitOiqbRbfzlkUMu0LIPRrs4ksLmrcXoZgy2kc/GQe6XqK06Bc2URbIJAXSTEQ
xwNaEIjro1oJxNX6hM/4Z7G6AX5og9oZBXN/KCJhBTBfELNCubTmAcvjFmSDSFMF
jSPq4sNIITgxRUmAHqiMUpiUR3n6YTw+q7dzv5wLg8g4seZLVYzGIDKu06zlq8PF
ggq0uzZ+A863qVNPlxj4rZTlYB6/N86MC6NTcfdkEV2bOKNlXQoi2AFB4tgty75Q
is+n7qQ3IrKAzaVwo/DdJKye8mOFm0RETXRHEVzPcZJQZ/5fjwlmIxNIMsuNZGSU
nB0p98z5UOiM/8qCIt7oas+qGYe6+6ecFcMpPQevdJA00mOqncisUcEgBguYiG43
n9vuEeWuzMBzvb/TPy9ejXRsBN4KYS+3R2OJZiQnGOBbO4bCkkn/Thy0oklKyuw3
0rO78PaBFAxYZcsUUWOxhAUVFcJMQHHecB01zwa0LxGzbRmP8xQ7ubpyEMwSroMs
nw3crzSsstqNdeoThTT7U8APeHyKa8ZM9TXgNzg0ofp70YlNysaV+eYNQaXP4N6+
dHPvsnJoLoj5m156RDD4c0DtVWbmL7/SajEDsdAUIx0hPMpdau0pnnoow3A1RulV
kHiDLOIFwffrrIRUFiN2v5jxwZ80UypdjAFDl8006VElhf9ybhzxcSE3sIq2a8dQ
aVykxmBrnrpwKx+NcO9MjAPsJOdhVDKK9CugCGP2AnMwq7b+ZaRN7c4omcvQBj13
N2tmd7qvwdPETN+62XWN1mSibK8iTUOpuLJqdeWAEjbWmyDriNAXU4V5FWMX0pZd
A1iXXYrqfEZaiLEoioM6Jf3UhvS9ZpKcGF9C3+0zlnCqt16blnFqpc0Ocpuafdu5
IFqiyjdu+zMIOmCt2w2I8ipmuqUbWd6Df2RPklyWDI4oBtBH0u3Jwptt8DQFIxWN
yEYcxCMWlTmNiTBzctP9+1q/uUHJcDaLhZYQqEADsiXTGnMHKEJxo0IdPPUtjEhU
SsMBbhAXicJO1thGNDKqGfTB+fUY7i+horAVcSskOpCxzHajJjZtIRx1MIouwqgp
jfBIwhX/F2QUqkdDLEyFgYlK/FMkYWpPchFrLDDOg4cEXcdPA7ZfWXMbdnO49xyZ
8BVL1Tf91T/0zz3Centgu/fGcyCHV1/Oc9vY8Qylk9v9F7y3eHo3RNiqbbmWjkf6
Fb2fkdbI6MPpuVtgkDzmkdnb4sxCBQpFH2YkgflskIpTu9J69pUUbWUedlabUSmF
sWVneEH4bnZ9Pv1FWtbDglUJRmee6kaqptsDf4ckyZr2uANx/q+DeGVYDjHQDOAH
Zof1fGS+b+FLjBJ3nJfGALW10fSo73dokp7OvEnaiXJgCNvCoMl9G2EfSu/dGNzV
cQFeKrlsB5kvxG/bPUbAE++shjz/xOaavBjerxe4TUylNZq8mNixrLl/oSV2Y4nD
5O/s0QmA4z2Ru8xfbXUH1MUPheu8TJncag7AkCBNaPMenGYUNZqCTadLhiTDP8/7
jxEo84DAyNMTH55m6YNgQOcziC1qfma8HfDH3mV5ooT+bgKBEVwKwWWTLHHMpKEZ
fpKhK1B0KFyU97acin9ay/KFWQ/t7K5bdOXtvpgbrw3mQs/ttt4KNbDkxJmBuBX9
XJaRkJ0rAwZmqqkLkfFQq0AYPOy/PVRkOVWsXgVVX7st1fqZyQtEFjYtoW+pgrUK
q9E8o9icrIIC3pWY4TF4ugnQ8rBfqo7BTKnF3bUbJWmVTstbhp6qbvY1f4Vc/R3L
I+LqPcU4Wky68ZKsLp9oiRD62OO/aKxU+muQ46cyWVTz0btzp95CSzEL2ze22xfU
Kik5UQJTLUkg74RjmN+DO17y9zVdlelwHV9GTOoNwsZZ/LeK3Q6VTwnom43UIHmZ
6xqRil7uXUJGPp44hsmBCSksfJbjlBHIr3FhDUe48snl+NZ+BtcL60z1qnp63DBM
O9249RAHcKgJc3FfTFpdwZY04yPzheNHA35vzc9fe+XrHLUX79dWf3YyA72jcvPa
xJB5R+g8e2A/6T9i9LpzioPqG5gpweEY9LB1Yaaa5h81RSLgtBnhOH//HhXJEnpD
uPMPhAB2kO9lNDL6BOGHD3LjFtZO+WKE1C8QTtuNVBHxQfZFzUHkK8ETMOhltvAc
LqSrcScrb0DKOxrHcxG2xqa9Dv9DuGa9gtixhGEpTCHl2Knq86RWdfSJbAldzcpx
Z6Cbo3KiBCb8xjfp3on0ptLZK1C8+1ocWWh7Cco+j1yLDycQARhFFbv1GZNeo0jr
519xduYI5ZZOVSK42hU6L/cUAKd5+Ee1dQ51RqAO+9vOWtJU4ZAIh7c8EaUGgdiW
Uv0N1jh1DsIcgoGcHC5gL1l9hkZn6cxODGaAbpuHdt9/8cfs4FjEZRWOZ15IgVeO
Pk/+SdU1PBuxPq0wqL4H8BTwG4scx470DVj/zJG1yD8PJIFUeUlJcYegqBIn5KfG
w6v4WldCDpg/VBsFw0NnDhD7LnjOc3ahkWOucBteGOWaQtdk0tOkM7Wc2/OXAKf4
0bd6JXpmvf0MLQyhtHjMd+6JHEa4OPpvM+PV17+UaVNV5Gc+jI487myT39c2+5bx
v8ah5LWIRcuNhAUIcb6L0BZIHMIMNYf/2L2JiZ+fKSVYOkZ2Zvkx8KmOEpwI01Pi
6Eta8Y9y5PN63sP/RGyWrt6oxB0yR4AvjXERtWouixJOhP7B6qmQEkKGLFdhdnTq
u+gx9KGA8CZwPgKiUuOE6cuqJm+5MSgyoGxJnbeunhn+X0JZjPwy0D/jm6hoXpY6
J6GnPQE7GqoXh0iYtpvFtkMvl8AwhukWtBhbFoCVpx6CEbRhe7ahPiHCUqYiWMmA
9RStipYlKl9p6UHiJcdX60n90VuxpXIklZv+xhxAC4YYIvYKTxMNoiGnfCmz8x0v
SmNcea0mz65BN1rK+HEte4cTR1mFbcpaNv8uQ/XuoHbzi36Lj4xY8RLY39uVvb0K
dIgTlKyvjEo2/a04U4DGlEdLeE1MdkfxPMkiy6L5hLjianUCa93q9L8Enz1sjaM2
K+8tC42EnL0aX7I3ifcegKh4/T8AjQ0d4J5ja+SswOhxSATPGfE2iMDXsa6xyAhs
PKBJSf3FSFu6K7ggRRYfqmfJRayPxkN2F17l9R66Cy6MkyVG7M7tzWi/Hx+tFxpS
f0PPMESnV85Bj/zZ1UqZfa50cTDoIrtGGl82gIO5Zd7WXxv2kvu/upHz3+7hqP2O
aqIVQsSyL2GbQhaHqhbh0E77H4FDMSC7rsuxf9So6HAthnLC6+gfRD4dLrgGwxrq
Wh/CKzx29RLu7OTUxwjAVYrY20Op7nUYoNqvvPT9DzZFfXs83OSLFy+n81nmNihB
K9lyddOfDazqKhlht8zWWmvgFNx2DGSIkt6gNUCO5MwwnRUpwOqxXUERvW4TYesM
7tJ6CN1hfMocyZYefiumDKa92IH3farJOgvSJ3HM3c+bLC1RXTm5gOORktZQhznm
8dLfiX/i2XkFFtZctOFK//XhPJryKP70VQ7HvZEuyBXVSnxjtiA9tENyZtoliXiN
BtESgM9W8vpf5YARUiCwOMRB7dmaEFrR2hhZ/iMmdPh40LIS18BogRYgK8z3NJOr
4U2UARkfMti69xdpyWEOZEoOlH4wxQW7cm8sXTIHyc0n8I48lSltrK/FTysv0xI8
5OPv3A/0tf+7dNtWYIyfs/1FLUuEYK1R/rjm6AMKmqgWe+xaVP74D1MqgBQAINpu
+j5Y3qUWZAXmN8+TCL7crzmjZqyppGxLPR4ZKbuWMJgDGQhvkJQUNLpdNgZsZjRx
6pgq3Z16mWaQcbWoRcWtyrQY46PuLl6S4UWqSuXO5Jl2aYb+5jywCCfDipoCIiN+
75nvXDViG3wNdB/7z67gJ1225dwV+3BWKpm6O8sf/dagzkXaaQDTN5DDzblnI4d3
QqAtaPxs7Mx4KJVsYcFKKkYwpEp0W32pv/FsBi9jfBSPXZjO8m9EBpggE5fIv65x
1PzeBXLP7ss7pTdwKJ+bF9SKLdAIHUxshbeCeK2uBds8nx//RXf+8dpVK26afQ2E
CQLRYAJS+jV9f7STFYoRP2Rk86z5TtY3PCSBg5sFzlDelBArGEeNUtqk8b4rwxU7
Hg+dT1J98xxHtYiBMyjqyWquNfXocqWsUwrnLbSn5VxWlZd2+8aDjJAb9Ptf6fQo
RdsOiBDwUcCXT+eBhivSc+pZ5h4y04BPoDGxxsARAji1AigwuXXsHXCFSEu9lIa4
/N/vxy4Nn6iUMeYwOoaq1O2/9boQSxGEv86eEFcILW/rWefYnJ/nFQYk4DISj4xn
UblxVRhO2YEBHjhG9+dARni9X3Jagp5Rwux99LzVX2uNFtlj7njipK4uYLW8Sa8f
PDhfMIA2SP4Gy2B7SvIstDdVxP3fVkE/iPWdzdHAZvl7h3f6iShKVU7gbQaPIU+L
wlWBKM1NZ+IuMHPTyl6QLFgRXrZZNHj266uUmGlgTbHlQcqCtRrsKXGVgE7tWetN
vUF/xXF1RpjKIRwlH4fDp/3ieS7HGEK2tEmJ0ZD59MURn+RD+wweJA03ZhA+RqHJ
Ek2GqXLCXndTI+ADRZzBVE0C2nNQ0RTMtb0OxyxOQSNhkIX4Rea3GKYN9HdwGgJL
T6pENDcFUpDtbKU9AEExwdU6SrNPkhnmxVZH5qVs77EjPjRnOl6FTBD2VtxXceE7
F6K2dD9SwZAC6vc3DXfwU4mzvcg2uHorI0kGcrpsoMTsLNUKOqzYOpcbShUsBox8
h3cJrXIIYqvUB05KD668lLjTFgu+iCuN6zRoq83AWVoLXgcoQIfQ+5pGmrjkvU4W
LP5Q9iPExDZPuKVBsI6NbZrcWUTQoaErF8u7LPV9Uc2GNcLWUsMhI+t3joqbWH51
cb9ATjhVWx3OtKLk+s/mGshoH5WUkb6pJ8B4B7vCmKBEDnN9+cSi1Z4eTLe5984/
BQ76iCLKfsxvD7g8NfPk6cwYqxyD8d1rWy/2WzmMK7imB8WY8iTcP/eobmXBQr5U
rnmUYDbRoGAxjoL3M9ilBsohlzqM6G/iy6qTVF0b03V8VK5P/rtLNDyOAUqzj2cn
nmwtwseRpI/mc7uRDiQSW+91D9WP1J2g5+mDjkYk6aHKkNRBBhZGnFG2yFG7Nb+I
t1Nna5wkPIV5mew6wM1rKwn1qCxBiK9yAE/8YjLJck7prq+gIkRhvO7YZki1tlAq
0Dgd7Fqa/874vFB9CcsOK8On3dUNtWwvSMG5qDvR/XTgN1tJNHRL/IPscs6/MbUd
90LmYVvLB7PE0tZRabmmpUuAvYlFnD5yKW8xQoNvp8OitgC4HudxLCjXgTDyLT3d
KX4Kgzc4aGEJk+400Hj1tn6rONiwmr4QJ+9DhH+y1zE5jrjpKrXIIeQchtxwzYdS
DfcRGDdDG+aQFz5GJE6OTxLwVKDlFXFHhlW/qatiTzt0tkRVkyJ4nf6RzMER9Oys
mMuY6kUtHiYaW41mjp8ccXYfI66sNywbyYfz2V6UiFT+aU0+TUCLSXvkkJCWFAAm
VHDMNMgitScKZRrJSBGryKH9cksNQ30pLu7N6Coxa2JOjY/aQTmDvnUkQYkU3ZaJ
9liQwHCoSSKLouJX0WsBPjchF878+4n9OFkNQRfAsAktv/n1XRbVXKGjtoBcBCfk
UL4AoZm+Jkrqj9u1/s6rfLGbBkALf6/f7imJXWRbex1lamX9Z596m6GgFcL78lMr
gTMxt2zZhZnhjrRoP5EIf+XfmtEsUfWTEpa1P+8Hlpk2EDRPsKSwA6tw1PtS6oLZ
RrVI6eOydr+zFdWnUuXF2BjVd5Qe7C4OeOrKtNg0e9SC6eliF3Ucttk/as3uqYN5
vzhIDhnoHgDoXT+TbttgPktbgvZD7wQbQRefEz25/Z5JH9VreBECSDPCV+kTR1kf
Qdcrv4RXFs7d3PwZOkOfXSLtj+H/2zLhTgEJSSu5a4ht6aa8TmRYplOs+JOod8cX
i1gmyHMJUrLBaOaQW2oEz4eGLEX+5mMe9zf+fS319ZmBbQrrFL7hh58IOOz2rwYR
vCHAPMXKrQMmy/P7tHdFA47nA3IKUZYny3Klhi8JE8YdZi98tigwI2+yGQPa5ihr
+8rabyA6sN+CYGXMEC3/8qtuvBx3hWaiJh8PuytZiFU47OqfAtVdWqeu97r8ElVG
lxkx0HiNC/uO2waZpm/+V8dc5W/cMSxO7VeJ3JMpJHQ/wOdKqbVEA9HAW9NcKePe
cao7i+ZyGDcZzBmUFF4Nc4QAFAGcTiC3d47ppctSUNw4BGYYXyuU+WlRQtfowAIS
h746p+KdD/t3Fv3uzYmZULenchfp8wh6OeeTsy7q0CP+CS3sh2CoVMz82jIk0Acq
wtA/dhhugqdxG3k/IZvCNxBNr3zgBLEyNY24tOAOu1mVUwadRyll1oSb50XUKVEv
CjdZHZxuVofojlWtHq/2NFT5dnnPiGDnljhl3FAxkrjo1FnvebZ60EL+vpSD2Zca
tWTo5AW7J2cTdjnLqbE/N2vmA+mk0K40VCDS4gb+l+6XDWRa+ZpCrtrNEYRzSPN6
Smq3atLAYbixrR6ywabHlnzs0ijALzHGKWfY1XvryDHCea3OG2a9hIdjpQRWyoRN
LV6ezjl256oMLa1K9lBDe82Y3o6Y5xHpUBhrtMZrRAACoCDU2Qmd3w+ubpqTi6CJ
2Q5Mul2F1K8ccHztBYugEIHivFVsocsqOmIQAc8790CDb3iimZ9ZCoMgqCt8PeLF
+GgEcd9Q2xGcemsSfCy9d5/K1+OrsGlOvgWmq/qulwFtQ9wD/fXGjALWHzOO45Cq
D0/7LDVOa72cDKppouX+cSo9Tc9ElFl984PuxYVXKC9jr0d0mWXSNYCa17GSFKnG
NEbiX2Y+e+cFWlioH12LPK6sklAfTPc7HZY98/Ab5WjClw3YPei+HDp/36TU6br3
eU6FWQzWNLAu29n57qTx9XTYpMEqZNRfk/dG8WzI4sxvWd6rJ1n06PCD4hJJ4bbN
VEOFT66bzLFJGA8E0JNDh0ybvhiPyB3gLSowcSKWFyCkH5Wfy4WG8ilNAhSBZFXr
+Cg1S6qC1bNkqLAP3WPuz52ySqwEc1T/qKDruzTtW6nQD5dSga4d220RE7J9x5Q6
RvPO3OxBMepv9azvSd955SCzC93mXUa77ddLG4lPbrcNLe/60WZ1PpDF8EqCiKlN
fj136ux7P4CrCdYGCttc4nPAu5dwPHceBBkX4IHnDm2FRKU8+0tJ6D+XOaUN/4Ks
DR/SOTH0yMWm1z1qXe+wOaPJqsYM4lAxdao/BRNA7gO53nzWfP2kWJDIBF4ZRCb3
JBbeHeX1GxzuyWjjK1qpTGa/NmNM37NOL8zSKrRnaH/ltAJgYbsaVs4sEqUUSsMl
tEyHSY5n8LwXMBklRd5vX8nP4RW6UKlbhsGU785krSkXMXeNp1iGGZ5eDrcTF8z2
xig/RyjzJg4XD/e00rswYKUyALUnYCox7t2SKViOFaVjfYy/1gTyl1ApmeGVLKAJ
aTzKf2EPV3LDwSX2SSS79UDn0VE0SEfbbS5HGdg44VatNYFMdN1VbsVLTPWyysmu
Cz3GMa+rKqgJISiW/3Ed80VcLUxPIvQbBBDtVISswtNp/txDxjnOk86LBR6O9u6q
jwbNffrTQ4uJlZKt8FKZjyunQQWyCFrL+lx36x8zG8zSz08ZIBPFkD7//nIaqis6
brMlFHWTbC8hWRn2gEy0qoIr0VsvyR0s2C0EJuJNKR+KRMVwq1RL1MRg48dmWmeZ
344fN3oZjIH0wa8cH+cP+uZoyojHKMSactJaJ2Vp810ruzr2wy3UF7I2RoDmMzqk
1AuOLx1if48usfPC80+Tv1DSrl8+5b+63/UIcoeOfQka1T/wfZIMWL90Beww8hf1
9ihPOeU3Lj1BRf9H/wiVYlei1/HKGVO6VDdTop9dJjeDbSBdJ7tH92PxGCuUvqi6
88uPk8wFdepMXxuh/oiNvtpQaxy3an1+n67iSVlT8L+nqfki7eEleFL6gABicEu7
mqpeV4IFYsSmB9WcJTc8kpkHuaSs1JKTbOU9s6UH7Uh/WsS6Kgj7etPCdNSJp3Se
QXcNMvGocnfUEh6ZaBYohpIr1jxq8kIqFn38yjBoEkM89xuTE3QFR3J3p4u7ARGN
OfSRXU4qmnJHa8rw15HcRz5o6yHAFKRJAQeOMXxFXlrXNmMwc5/htSbIBuR/t6XW
JHqQCAwDPe7AEDw45K7HSFq1F8m8RM726yYgrDO/xi8Pzsf3gSaYIZ/lu2vQxB9w
t44jDvr4tI4u7JbS2kduZ1Fi0AkmaSqFB1qyAiAwUP752/MfvB7I05rp9lvuxrvi
2HyIPQmGcvsz+LksMi9LY5wfrpaEQl63UbCKWVMZ1/cRF2m8ehno6GUcZlgVDBvH
JCYZ9xqfOLxJgFtClkNUjpZC118SFwSDYObKxPCuCprliinFCtlCLYPe1MGohoad
mxpPc+wRRLELti31REmPXNcZtmbNluGAVlIakp0I3FdRnz0CoCmfE8PQC5Lbj0F6
BBghEa1+cz4wAdbTNl0trT3nYPu4oOXj2vNRxu13g8kK1ViQDEJl6xBlo7sC941I
523Rwr2TcczyOE91UuZr1GSeEQ2qjn4iDsf0BTwNG5fUSkjPsKHavR3AwbXOuA/5
LjZhOtdQB7VBzZdkIlynoXptlAmtYYKhQnAQAnF44EiAjU/DEvMVrAZuBnWpVBQp
4sVekYCRFLwwve9QA45FOQfZlIRG5Q4BJ3rI+esl3LOBUhIUrVqNkU0/9xj5B/QO
WQiB+7DP8FhphTGH2ifbr7Ftzn8eURb8YyMg7kz7PMO2J6TcpwIhdsj/AojCjJW7
J+heV4ccdvrahAsWCp6QKQVoVyJBU76fR6ntEytmq8kL+JrDC+2njDtaCIzIBZnB
tJKNAFjaE1CnBpqqdMmIIt+Ci+t8QLcYXd6j0nVwj6AUiI3JcLyiCysgH85se7eP
GBOqtfSQqoTLC37te3LS2rjuUwApliCYX80s9zvT7p87eOnJPy9Swh5GojyfPnxz
1yinQbaP4Sa1gzQIDeaym7OZsPd6R31Wjd6e5p+3+LlLfXIOH8rFATv9E7JIvfcl
1kaUFZfS8s1vOt9E3c/l/7g+eoMgPCxdD0aGcay0xwAHpoI2NoHZA7IfHrkBA0up
Ta24FRD2yTIDKIcjUo9Qq3E9NccdIm3pRiXFj9C3FVHYf42m/qwLPmQCTYtOryno
joJXhuLYBDuJCG1pYxOFmW5hlPjF6XnpYSfSnYF1RsPkhcoHAzemfoGqcYAVasH1
6D+6VZepPDw0sSJuEtt9huUD4W11PEebci8t5nOHB93hVG8q6eIDwwxHeNKlyL99
oK7UWQqfS0iMyKqv7DOWHF2vwIkR6YZs4TakSbwTjHD4bYcsFejOqHXi3yyGCxCF
ZsSQ7nGU0/KgrCn+8gBmgWZZl3LlzO+f3tnjrCRuhLgNd/eXP3hDCn6sf44UZFuJ
JN2kpQr8C6Bb/PB3BMZo/Vt6l4u+RERxvbSiDf7VQ1jnBcX4IKLig9OdlbmxemFF
/Fvl/Z8Gmh2pYmT1cduazD6apTWnoWkLu+OC1yO6siOIMIWidt9SX4IcLZ5/LIP2
BmF2D/4lJng2qvwgxLz+xqpMXqXClPRnr5qHH12QFWxdPO8FMZ/wCwBaY/Luhvnr
V57bL54WUYf/dbMG2EbcBYnFhcRCFlBAaC0c9JarXObUtYsZLUwHjqzhd8am3HKV
npOS2KIvwh15rVp+EV0Y8fnoFeiSbohzd/at3/aKWro7wf4oF4/l3AR1iVzBgKer
wJB87jsW7H/6t5BiPudSDXWdU/xLPSqPCF5q5A69YLQ6UPYIUhfK1oXFRnUnoJW6
+nM+oJTItYD9g3AK2LlC0D0dozra6CtG7NivlXSyQYuHbGY/E29Y3QwSEJw7oy0t
TdPJFK10x88VTmjZDztnbHUQYUECW3MeRGarHXryKo5ZRNgc/QVGJxGTD3qp0x8D
qO5+FJX6vIdaer2qUU19mu1+lRU+/hVAhmWnBAkoMLoe59sYZXIc9jKMLuHE/ySk
kHvesfBxVEOyL4CF/idC0iYtQ/3ypRkXQ7BpNFlPwewkgz6LqcIRHCUhqlGhXWwe
afdjkH5zy3yxJqjYE9RMgftB5QO/SUGIDu3REdvfmdByyMzOZFSkORO/bsAYwIR5
G39p5eZOKBmxSsSPbT0HfIUuyTZn269QzDCzKeBMy20YvaIxiZy2mSIbwGE+1INo
czsE3J8fZWybIGujkeBoEdHIcZUT9Ix+EGdTD+OUcb5fLClx5Td/3gxDpjzRjJV9
4hxIYrMRjX1gBYvwjFE90yXcDY6AuhhwBoVMQVw9CUnKLhKa26X+L5TRt1qncBEB
525TXMIrySzkxtclI+r0D0r7on0w14Z+NC/Im+HoCaxIziXdSQyMbhzORrWLHi9c
wm0Ea3OgxI9Vg2PmIl7f6KpaiyidlQ8/UfylsYiEQXqL6K//RNqQlqD6Sc+ZKB5x
UTaGmlykPGkTeWl9Tmk16Keo5R6Ujs1znxBgaCjMNzTCIxBMfXpQ1+ln6mirm0E7
Fdm0RqJOi27pK7LLuPcU7QoJA3jSO+vJjngPBj+ooLDMQt8JbwQs8D4icXsjBw4E
B4KfDmpAF+vf4lr42kGJzR+AZZtLYK28H3tbKWepojcLykeQK/sAz0W+qWymva1Y
1DDQn6jOHkQdioFxLlhQi6s+k137rxGyzIYT5E1NvIdPOizbE4S/QoMFQt0s0BCB
7krPauvNrof0cXTzmAnzINa5euvsAm4YAy9Wx0Kvixy+hTbn7nW/6upMLF8CLNVW
sdZTxG97E+t3ehSxjGpKw45iHKKNECQN5vE3/CNMEYDboUFfqoPbDdKTxOmlXEtO
7kyWTl1msFVpqVlWa+nSAbTkeS8ZzBWAt6lrE13Wgw81Uj9JCy9TFFias/g1DA8q
g7P56PbVbtIbpw1AE07QBJesg3dbm3sBf+BxBOJQ0OV6L9TSFW3wa3glOUqGp/Ph
qJxpOAgrPcXR7WDy16PaWm8ceOBCw8+9SENZb981E+0bnNrq7lcGCCbi6GtX0uUf
+6wbtFCpmpomHMelooOwLmevieVXwpJQffXG5PhXyQ8molm2Ryd9nxegwCdukS1F
tczvcE8Uhnnhrh4FDuJSph/KG0pl3gU8VuvT38nmope7rKpdvTVzEXt5hd4NoaWW
u4T1qzAr8tnieStLlrXmuaCdBAIzMLeAlNc/9vqG66C8JavAPA8MqUNwoJl836VY
KPxzUGy2wOxhYnfbKr/Rb0n5mBYxkD7bpPX9mWuYEa8BvKh7Zz89+ls3emrJVG0F
3muwZ0of4A/INx0UIalT1ZNI1aVOH9l+DSxRRHoTwdqncElG+veX0Qv0RWoRUu4G
yQNjcvxChQ30R+nJpyQ6pExSWIT1cVuwk4ORsG+5aYPvlF4Lwnt066jl70M+6CwB
7ra0WNdHwAjIxvxVlycqzvJO9e8NVEZT7I9cukx6gzXSFz4dbkxjqjbSLZ+Fm+w6
5GXmzj0/dzq+Q1b34sOT0KBFx9L+cIwucNhd7VutdU/Qfa1bMPuRf/arg7ZnpasR
eofkor3RZ6JAs9jTZgYPdizPWJy1oIHtLRH2SsrMDFYN10V1IPZ9mVgI7/ubT8xI
pKxxOXOQZnFuHMRLK/Fctpkdr+ar3EA7jY66q3aMFN/Cnb5Khfc5+KWZPEGL0+hK
v8SMdjkvL1dd5QBuOGNfKW4oFS4bBNnRWGpLfjyofGcaKe/or04i0wxyHeUXy1/X
OZJoiaq7eCFMnx2hQ0B1s89inSURsFnF/iAGNuNAyU86GmJaxSDlXUwya14nuAih
PR2qYDZ7Hfx8EGD0K6PgHFo7Lz6pxFIZ8/OUHVCeWB0W0Ejd03zax5Khag3yjKoY
/v/CLmxjZqcsEJAgQwojT0CxlqSd+gtuKsWvzJyQABL91OtWPDzFAlHsBvbiJX/1
X9qekNNxHZcWB/iLZcm84cXvsOXEPlqNNCCPDBONcRwImmOOPBwso4EwTPg+e27k
8xJ1YTrncCrVxC7cEHnZrGXiBJwVBlbcTwgNGGRvP/LEU9aCbX49gK7+h5ppI9HS
E32qUcUY/dw3O49zAgMKXbhQrbDjrw5C5jz1ClMno5xMsaRmjGPLArqpR362H3uU
DNVru8CebBowgDPgHnpKMMU/mQKX4N/SS158Ca0P/jV7NJf/h5uV/qcF7o7pepNb
KgMiZ9zmEfE+gn7HJKIJe7mivP2l2KBzISpMRdFuPSZVcPWVtHc3L1RC9QkfzQZ4
A2ZlFP7LSSpkJdwYV+ne+L42ReBJySHJ63QB75lK8lIBfJ66KVBsAy5Or/4wcgJO
VIIHE4Dd8upEfyQEM8KALFhcvETJbo3XuqjnA8qOhDTwqIML7Swg287K1HAZOZdt
nDyD2ykVxuGaKq66/juDplnI0jpZg/8YFM3f4HWErGRPir/zubJh17oxj4Ih0Gml
avGcl3e7JDH4jF9NWUlr86Ntb/v/SsDEV97nzMbpCzwc+paReevrLkP98ajd2o4q
Lu3QLI9Afuc+6rPmDd9dIO0KkhcHkRm7RkxXYa7d7PVAKhihSOOdyV1QqnkZZ6RS
8FjpgfDCU3FJyZl8bLXp1lkbwjzuIPVv8jK5zDOUzNDsUG6BmR7LeWhReKXvlOYL
9AMyLG0paKMQ1roAIMlLpBg1a1lKgYACGAU/wTXC3sJgkL8qSYesIx1sIvy/nCNb
Mgz+J+OwwNs9CaluLU7nputLo0T7mNvez0V/tqrLxhXdJjQeotFs9KGHOuZp4tbh
7yho4PmQcZR4h3FGqWdt9WGSFtkddqnOeTNGMbTUb0yzXOXud5xO55Oa4SwSeKd2
nlfXWDznwVY9Nm8brCNVZ8Xw9SgbfAbfWGoIryF7ozSbaGFzI1t2xhNWAgeC3Ic2
WkstFS2j3hnLrjUFjjb6Qa4FOXhBy1ye+IwnmGZSMxxqPZOvoMkEH/H949ZIZ5gn
r5aEyp2K58Lpmt16BBs9ZINWpcIQLfOGIRf5WSjWtEUKl5AJR2/vZCTq/KzA6sxo
W6MlFrCMe/M+7P/OESM7ujTXTSWuA8eshy9uA6ImWx+YdtKbhYcWbE+ua4N05Cbm
la4ZM64xNaDBsc5wi5Q0GnIEUnss8eGvw6u/gFJxtdMq81ZhLogbb4FwHlkR9vMg
MsjG2NvRbpdKgugrPz5l+5/nobh47rxcZcU7aMuDGXK7NhPPJrRYotLbyykFjhuN
HzfobnDvEHePIwQjuA0Vr3c5mkZNRsSCdlRjocpwiUzd0WT3RBejBySc4x3GFSK5
cdetDG6DWnkuzGr3tVcNLc5cVrNkzTsUn/YKM4aTtipewTGfdn6fcegEbnrhHRdh
aGkKMSPzpzxnhYXzF2efiV3XehEoYPW9aaZ77Yh7RwzoacbJPbhNLOLk5dpztrs+
y4nDI2X8I4nGzfP+rXhF1xrGV7Xtr1dAwEn4tZpX3gzxbBmFEQedULFd1Kzg5cS2
pDUxbbmR/PfRoTAbRSiaLkFxIf7aoEM0ZDBDyzI8p3p9nQC+F7d5h0X7eezKGahr
zJojVb8p+1tY4Rs6xeYy1VRLV1HicAAlVc7kP6C8BWAo8m3wTY8MiBjfNwiVrzcO
qLfgYOH7kmwIefq5m5tWdofe/IpaxmLYvjulMRGMpqg+UpcKNL6PwPvK6IMIQXhc
JV0ezkpI8nLlwRq1PQJGy8PL+fnuKqhcnBLda/XPRIPC8VYH1hKtBzZTKHOXkPsw
ep8UQrRCqRUmhgInSO3XYSlGy8SrxKnqhjsYZWykN6SkAsjNm/+lD9IgQP3CB+NG
Mi+XvN7cNGUYuJ/1yZtyuLHn3M/HzSYGzx85FS3sYv/xS29pRQbN5U5BSjIe9jk2
R2idPhvHdwcr41LHD7JRbbC7ujFTpqibJrBiy0RMUdLupQxSvvQYFM1w993f9u1q
2xPTAGaDuhfZT3hoikGkZvs1o5ifr8ZIg+2GaFahhg0dvZBJJ/nES3XbaBkjJCSe
RTBSkI9usdeGpnvlFs+ztHcMZEhKLk1AbUs8hcm0EUfa50dI0pcN37AIbUNYKuWD
4j7UZfXRhfGulBaWX1AMmZ9ywKgYY0wvTLJyagQ2PkeR0WuCOAwKexSxYqRIrDUx
VQnehhPAgG/uKPeXMSIdH6xXFGF7o+k/qRdCAJ/NqJRthp/3GlUg5E5Yy62vjvZS
UTs943eezDVeoNZL65smT1QeV0DrSSM3LmDyulY1IM7rzCFEpdu/X8CG6UIOe5me
mGfans0K5JD+uBFNXWBPN0dvCQKIa+PdQ+pJC59vfHApyGabBme9AiriPOZJM1/i
041HJ5zIrrERk8t7mvHUVyLbYpMT4M9cCP6iYqM5BNCfrla/5fukPrL8lHYjWbnG
uB+wAYeLcAre9dyuJVJWPM1gt+IftoBGfFV0F+fdLPRUBM3KjyjA+NeVTY+H/Cvd
4amCselq2GPVYO8RKM8FTyphh82KB4b5kddOdN6WTe9+OT8HS/LKmD1CpGqJMKh3
/qWaeZfCAv1Lpzm4Iz7jpqHdkrBH/Tq2OlFpIZ3cEUHDP41mhEuNH1SPBITmjTnL
iR0kc02nrD6nVwz5+IhDM7JavGMIDvO48P78ET/AfiRmDgf8Z1QEycLFijCMv7uD
DRLi+LTbVFqjCGXCgXf5mW7ZriOfDInGIIrfvKWZuinkEKuKRxRVZWlMIMq+gIsL
uGOTj4MJx74zsqx6OLEn2GMkfYgtJ1a2Hj3xCOBWWMSymVsan7LJS17esmkAY9ZF
d+2G0vxHk1r8/ekeuWP9pew5Q7jj/meWJsaBXjugGiylv7DZV8qmX7AEkdWEGPIq
DOESUr5wl9UvYP8/sbfaFOUK3JCCFVc3Ye0I2uUIINZxW70eA32lFAgMNjVjXlWV
dfDruM2Hj/OT4hD7n/UtfMoL39TFa8TiHraU7Dfo4PgTvRIv6ZuB8YPzoGdk6f7F
0lfRJSTUu1ez/QJJ2qtaalPXYIY0NgQW/H/pCOroLeUkQJGwQPNxxh9qWvgvT0VL
QeLLdAs2latCQY3vOS3A5FI9154E1UtsOE5+T9igdZd7Jqs3GahE9w1l4yDSng7Q
rQt2aOMn4s3HcUiy+vMMPOJ517sBWlfr36bwOuUvgw4tnAHftr6yT82EK+xoO8Vv
2/alNNCLGWHbt/aCIOY4Uztzzh9w7aSu+46F7zS/DFbiDLmhKkt+Whg3W+aN2LmY
cQznlybfhtwAvLlPx04U0S1z9ApT5xT8fgKSZBf78SItxfgMiYpFeG6uGCJA4Q9g
wSye4fdcnqJsdrWe9faBPDt2EgmJMr/pqxRLg60UNOCWKzXXE3qa0SEEpJ//6LaH
vqoRULB1Mr9Vu+ZBwbwEiVqQn8F8JeJTXjXWJbolpa7nIdSx8azMJ/pOvDYCCLkG
EbUS+p4v0TmQzH8ycRm6mFBWPxqPzyX9ls9QKxm2QKHmt9tsOExD6bEyGExMb+u9
z4VqJJShmlMEtOYxXYaSFoxhQXuvfIPo7T3dIQOoqxdJ7LYI2i7wb2uYKAQoYsxm
0E4j8j31QY0gMOakpnv6zjabQwe8snFY9rd2vkL5W0CPTXH1WQmf1r9fVbWDjDS+
nUpZGfWx04aVP0ELHLIPDVUvKqsxdVUd46iAKDD2XntI3n1Mm0JiiAHxHF6pp4UG
retWW1qFj71pSoQNSaKhCgpL117j9K1pXSpS7CyYnGggRx3S35MUbtH24OENCnpb
HuaDYOn8iYtcJPgNX5UnR6ylv+dNaZd4kMddNQERU+5wY4sAwqIAqfYNO6Hiq1/y
a6qBy2TUqKLQ00gbBax8p6hnHGkP+ZJi9q+GVkhouZoEkADnTZS4qm2jN84Rwphv
NHxj7lCfnUnEKt3XA2Ld8hJUVpqwzxNrOl/ZQ1mxoNoATzh8LLGNwYztB0AOPz+X
qL6nwAwr7Y+sKyfD5bdACaSSWJcGXYMo/mmDk7ZVyHtY6oVGmIbTf7Ufs+NAx8qN
zccLW7gGCjJQgzl24i0EMYXgGz8W5Rxbzuy1mBBTaFj0g9AAIC265EQYvSuUnAEO
BSvlfkoR0dJjEIFvavKQ4ONk1wN92I9xkBviThw7/hNg1d2MeoGzwPOCGIn4l+P4
s6jC9AMyGM+9tWlU1DluY3DYgVp45/QdwBuOdGe+uQ8S/8b+lI3Gn1bdErkStvAC
on4k9D0koa6oaAav37hfpiH9HzkiaZDBNS/aF8DwvwCHsoP1yov7YjZsSD4W0OoP
jLDyvI1Uv6l//4rcCCtNjlZ9pv6hh70fO/qGJSx4miq9w5DLC3sFcuRrP62ilJ+7
VUsXMxVjnvODlC5x6QbF/kBotyKz88cAN0f6sR0aCkCFgNfo+lTHrLp+jSl7llOf
O6O0s9z4CCZmpt/QAVk/8vYyRIGojIV8qJ9biS50hrM7RmkOn8zYeUg8RWhZ9E5h
uMBb2b4L/aloTHSZf/nhSN3JOkkoqku8zxrG/y5HAcfEwVvtnxC41znwOswXpGHz
8nkie4JC5ut//Npu0Yaen50aWAAZGsr/uDL7GMgBneNGDEaLHPTUVczZv8j4FwBz
4edlrnVKYm8PpHPgxLajty2+0cPvU6h4RH5Q/LwAOxvtW9QX+BpPV9cg30n/fuFV
bRA+MOis3LrHz1posSNaxHgkEli4+CdJvS7kWhETKLl+H/VHOUI9rRydyNMKWDDQ
y4E7b1EYXae79Jm+kXcycht72walpcqXIPNWEMfiW0gMTuY716/AQlWtd10DZe0F
qLKZB4JE7YoC2Q2rPKkrSunx22kMdI4ujEx1l+TvM8WOEearr3GSEhZ7XgBp4D53
9kE2vqogmGKCk6r4meIOrUq9oa42asb1qyGLfSBMWTmo05Ji/gbY//fj4mDIbMIc
dW5Jcu4nAePvtnF+KCFVfigI7ZlTBM43iZLGc38zUWuh8BJOK1oJQH4E35YrWuyN
yOFS2Vj7HA2mSU5dZ3rR04i9DxeLDI9doztAMYFegR2iK+0f2QV4/WmMQmzTyoJF
YV/pJYBofQ8+rkmLZuoRxIcc9IyhXbJf/hpgnQAl6KF5ZlZkTDWvMP7Oo0ACedBe
l9FDBi+iKHJkNMbXK62O2FTQRBlfjDJ8SPKYgpgXp8OmYgq+w0b3+1zbuaeEaVCa
UfSYUx6FYuKNcGEuu8EPW6iujCA5n0tF+Frbl9fzqWhX3SrjRZIP/37biRptZWVt
shdlAYhIOdw1aqGIhFmSoMgAWOK7T8bK7AMqpdQoArDc+NPBfwkz39S8+dOdC8BE
NfnT+XkyMux/iGxRJPq55Y4EVcO90/mP6Qx8zh46MCVFRChI0xNtDpIkj3KBx6Q5
/k4hu9E9anwBRhPixhQCS0HLeVcxSj3HRyKD6zL9mPoYn3hi7M/rr0HRwslbbWt3
leVx83cvJycPhtomehBMpsRLrtA7HMbq+SfyAih1HRWVVjzyhCoGs6B5VrCwM6k9
b6dE0qAKtrCRzay19E6YwtDhkqB4iwuaDCVXCJrm2siWoEsZRzn43yy19Fslnxpg
lZa7f7UnJQsUwlK6/J9PoX+kwlWPnerDbCQhKNCxjepYbUyID0Zeaf0FfHio3UrB
OqUCYDkD5GU4RoQdIzQWlZ+d198ORKDVlPbLiUn7ACEr0nUBGi6PbJNQD1tpY5bJ
Xog7c/Pz/SWi9xXYVpHePL1f0Dw8VnBoPx8PfJWHs7YbPPMa3pqxMlfbNrEPhS04
n5cWsE3jb+CAjd8w3fE2fc3alrY3YWx7SsGRGhv7wfSDESsaabh/DY5chfCp8HjZ
eR+mU0xANY+O/dumudFXPLR2JZkja/VBYEKKMxg7m+RqBfA50HfalfamxvBzRDKM
6si9QiuqYPYI17H+zs7RID/Sy7mzb1TRIP2NylIPLE8vkBvpLk01D03znF2snIP2
nOlA0l4IUYZ7STMl2unBt5ZCWyWc6ykiaOqcG9RDu37tT3WANKw0/mL3p0kyo0gT
s8N3A+sXum9szucGcgetYyt4eJ4tk7wIbHK1SuO2bz4VeYM9ZoTUK9q/HfkMksEq
OzGt477yqMN3Y1ZFI5tVDFLY29SuYJ54pWnECswPisvA/F01XNEJuSar2/p+6rFq
ISnL+oOzh/UtMfQyO6db1KtZEDnKuNUL3lXR6I4a2zeiR4abvsk7tLe2QIRnFLz7
yy/7lgYhfmFt80bwUOI39vlpuYr+h5QnqAiAgC0m2PUTOFCSF4YeioMxB2szsAGw
PL0mhB+tNGiN7jd6a80iNp8dDhwEKPl3bsJYIsqcP7EUYwjfI2dZXQdZVc6kGqp7
YiisltXgfL2tDFaSHr+ZW9/l/MCzExxjYfWglhQ9sgr8IdXDJjQYhzHSBdI8kUVw
5rq3bXY7IHYP518tOzLBYsaqjgtCgR0cIcOzulR7FpAD38GGfOGw1vH5KLQSz/ms
gMkS/PEYxwfBLP9ZCq01LECQIwo+abXYpWXa1wNhl3M8PZF8+IiS026a0CPVN0Cl
C487kkk43N/S2uFnimXgNIS1o3AelklUetjnb4gbGspu3rKTRHJQ1JMB8hpkVPIL
1p8pQUNZ0/ISsNcNkWaoW6Rqy4R+ykcT/gL45Wk0YjNShB42oYe7FopKTgkKVl5y
sIG1xdFd9KG/TPE9mLYisYTzgVby8iPKFU2ig1ecsSEmzeFvUWjsiIfU8Wmw12l5
Jbrun58AEUR4Ln3HFVSK03cjOMw0y1h0ZEjnm+VFssB9P7DG88UcBZ2xpjApXAZf
7iT3hKWFNjIzZ0mfzbS6YS8cfXBJ/q/V+NRmHqCuI0JYjp10WUdd/7hacaiEBN1H
jP9VQxygcrt5SFN3Tq7YM8bFD/dq2Qi+AfJ7VsQlabp5om4sHRdRXgsFPkzubJtI
l1b/ak6TXy8yAjzaAJsJJXvst5EV3CN3d0uHr/ZsQGXWt+qPJevupvGyDOdy03Y9
jwlBHeWvocOkqzRP72VXkKZreI/cwsLNf2roVkH0zC4VTAYru6rtoLSaF40WPv6l
LSVyPOs6CtjDHbwhXSgQZZwPMxQ0OxNtJu/PSf6g4qTAeQMFGaH8AIWvXTH56RwZ
4spbaF88U6WegBOVY/wvU3lPkfJ9DhEaJfVh5yZ69QckoNfgdnS4XBbAOuNTu1VT
F9jYQxhW8O0ZCLDcGFFlUi7kYRBnMj9XIt17GZ07KOMN/HAk0oT2nvjyFiY4sKQe
fNEzsDX+5jOBK5kDgizEQjaWhtMUJfPbN6sLpfEZtjBfhSYWOEcvPF5P5T49PEF9
hC+o8iHSg/dBeH/oa8Cx5m5v9Ts5tnvStqEy4hxX8aMvcHqecObOPlG40rmhJ1Wa
RxavGiZaNwNrPPmft0GTfa1XvLftX0AZE/uktwUP/GGomaCFFMtDVYYdHf2tYmGf
HKmA7FUxvv66i01V8RRmMu2WwigXTqRTx+2TOd46qiON6vjlbkRGi9naAY6z/rGL
T2sTmznYQEzoBLoMc36dlLnEUTpBHDmJIjPUls0UKlERGUya/6Cx2XkRLDlhVwel
+UcD4yFStQJcqICRlejXe4d1bhpdndsWMJWeh9eXAId9a6IOcM26dvaajMa/Hm0+
F70n4iqse8B4/XRveVz7fTUiQX3Dwq2NX8KDg/KnZkNedjMwJzmJnIuqNMNku8YA
S7xrO768G9mZcv8iGlB4SS/iMaBNTNGhbsq9RILXHyTP4TUkvHfbvvbbtwTrOBdh
cHTgK3EmxOsvmOr0Togx2nmcYgiW+uu4ydLW3Ju/HwIjFWS7HU7P59MCYbVf5CyM
JkT+X8a7M5oP3VKIhYnI/pvY94agXRe8/WlU437pp811SjEwo+WeXeNUFUTIntRv
uV2mdi0Odk6OsqaIyyCpIRrmif5HvSJg/TCjq/ky2K5SYQAhC/Rbuw2EcwSbflFb
5u2GEQa4gKuLopJBLAqf6ElyyumGL8gx39zrOBrJvDAwqVUnEdOMEfZyVRmgSrjf
A1wMa3f4cDoQmOgVw5ylnfJeg/Uz6cHc1wX2umlNliM5MhmWN6QTvQJzzY8Xwffz
j7D2sP5wCubJFF6iKjh8lpHdbGc7YBa633YRv4NvX/6q7fwFQTU7nb83Ym4TwVXx
dFcf/Fk/VIMqaXlPX2tFuidro6vjhTK+3wUO+Hru+XwIR+DYuhjtVvfcUyqIhk4t
8uVEXFbQ79YG/KoWX0/KJlupgmXjBwzB9LeamuMsP994ejbXUatcxMV4HSMj5OKY
Vyhwa75roIsmxyqSFhhjXdNBQozxtihFzjPEA9tEVTlxFd2rUiFkzFxbZgCJU67X
CGipdHSddxCWB5CNfI9wKaMbZaloiXMWO0MCgtJYJ/OJITKIS9EinrbfAT4Mp1RY
Dyj3gTrBfc7NZU7cWtB9wDGO7Y2Mp/CStDsnQSEwZDz6z/R+SRlQ4n4Zi7vacUHH
jiZ4JhgA3jN2Rq7Qqe7Lap+04CbZqMS8ILUlaUz7iSv1teh7FNL7BHgrTh+l+uQV
n05aYFi3aWBc8N2ZRhWqhlMLAxvwkIsHus1DrzvIJ9F5R8eZjuznp17pLL/oxCCB
/2vJXtaccudcTucq1eT7MbrBh5mq/kWC4P8Rz0qyylWyoJk+I6L49elS8lXi7Z2R
0QRTIPOLyzTxYtXvOWYbT87kNYgtJqhdN42KSRjxpqa+nf5nhbqPRMdxDoF8y/NQ
MeDhyI8H7fRF1kwXu3Safq63Wkjv/sPeC5fIiq67xhu0sYrs4NpUsVBGsrWbZ445
V8gIRo4eh4TCfABL6Mj3c7chHf7XHohQIHsbs23BO/pYM2eVYPzgU73mstZrpj2W
qyzdN9VWOJR6Aumq7hg85TTGiEWk2QhhKeKGVSeoMHeJ9b0iXcKM27VYCzeolMbp
VcER3dEiFIA7Pa4/Mxg/pLbmz9Mkk3ecjt3uCY2Q7c7ltuHGIm87/xGdDl2bA/vy
Tylnd0AhZjBeOe3CfDrLqZFPp3EEO2yeliw+6O/GkrZNtdZ/MXjY1owAXgb+bAs4
1cbzHreyy+hNuPKseKff7NDyfWboIVD1pjKas4RlRYQyufep75INcXINnCPDvEdb
d2TvwMY6BSrX7AdeQ7AAixz3lAOFzxIQlFtD9J3TWkJQLSkNgDZObtpXkPBgzYcn
6ohICpaMcsd4YgqdOHr3eNylJRZcRHa6Hjsg2cFXJXVpqmyMM/MQIlR6WkRSJw0o
F5fM/kKKufc531Y1TobXoTpbWIkX/QY5TZ4igKubYHPG4ZKBbPHtYX9qDpEhku49
L+r5tF0AcVl4evyWml+PBFP5K2oTxj26x6k58+KVLcgcYQ6CtpIOSEsbcH/JnHmA
iTyVpiUPYyUnlaX+2OB9NLAV8T9frDd57WjxJzi/Z63X750icdJ/1GmyDK65+Pz0
KS1kuZ445HK9cXzp+0ouLM1/mLqsAc2AU2WnOzRz2SUtMiFsj/HJjw7plAIqbU68
jeIQeWHhP5IF8WmQDJmJXZOi9/VTKw9FtRLpW6/WXbsYZc4t9pPFDF2MC6BMogj9
59mF1Na1Nr2fYf4fKu2BN8eYrxFodo6mycPjfNyeit8njAj7Qj3fre+lGcc8IsKc
dGz0kJBmSHkrt4VYWWdDVqmlCTmRlm3vD1XJGkKNLxCEnBwQ1yffbSPN4gMZqhvN
bfoRpf2BZJnWvnLNJno8sJgwIaEBGMp6EgbVsiuqe1ucdJXid7UaAtYHOWLYr0Tc
/cohHz8YkL4oqP9Fx48zZyCN+po+XfcRzl2VDcAknKHTQOyCeFCml/1G562M1HKH
xo/oszvZ/KXtVZIK6e1eu294/kiNaK/0zSlUiyiWQjsMsDaIn8kPBZk8mKLOA/MR
tbfVya58wiq2ZFIFT4BXTbM5TMA6G/WZ8TdoISJOhTnJmdQ/4+Io3gmJMKxzaSyQ
FXFFXbH6T9X1aFD6CghRgQA19E6b7Fs2KiIVP7EgBkPB5w+GzEB+xDrQVwhgXh+N
4smyHlJSiNaZpoDaSTH9CPGYQ/L8udf/mxhfiDgTztShIxeL68qqG+vvrUpy5SIq
ZzzlrmxwTMbdZpXWNv7ryOIGzez7xz16CZNsULMQCjWCV28vQrh9QP5I+2riVEv2
gV09EFc4skY8V7gSfiToD6DbO8Lflbg6ZHk2KuevxAoLI3F2FwNxVgm8BzgTpQEO
FDl311zopq7OI9G8sr+JF8Cqyrrow4/5HvRzsGD/LT6adn0/UR5GdVaaoI1GtUlj
dmyQ4wnq4RJgYYdwytm1IclPKcqYK3fz7Ehh1TzBL18FSCU5rFojRtCivped0pfY
PIg1LKItbOXMSbhHcWrjpIRazk75WV5BnDyyA0gXOPnJCTBgDj4b1kzDq0uV4bhA
/iTOHB1X9wjgO5Icx3N42ZTxcQFdJQ06t5DCLxgG+Zvn/wTyE1QKAuqSj1bkW+zS
ixTCEBRkdm21ziSSw7h2CLkO14ep8k/DcD4u+1nYnsBtsl0qYBjLYT6A9pYiikRg
pnNSacTMmBfU5EzwiAC9iTVVaqblVwcimoFxPcN00Ve5wjO//Aa4z2NAL4dBf9Rj
5l3krSg97wbCWwjN4EMprEPyt5lDm38SWUYbLFq+2VoFi/3AnD2lOnCINbfVWYrM
v7DxYKtgYEjeyDYKWifKbht878VTijgSuGnYajLuMSqIHXURobmnGnP3UTUJcLyK
nqVMwpO1qq5XRTLs0A/3EzZv1GtEC2yNPS3xYAoHjhX5qYcfzHereVcr8/nzpYgf
BiZ9DzfVf2fgcP23Jr1+gFH421nNIvrc+iJ45bbzE3kUqCSmccL5ujutjLVbl1uk
qcFZWhBWyAlJeDwaCiH/GfvC+NMIaCcp6jMsGUNVFdygoDBvPx1SeqOG7rmxyIxL
VQJmyWZuvpmsCuemmFOYFSPorD0a4kPJEXQWb7e6hVyCeXZVrrOgzf4wRrymTj58
k+7KXcpM1ohuTIrJWiuneMV7rUFa5PRZkOhV0aNQ6cFbtEoesPGRz3YYkvngo1YO
cK2qldCU0MJvQr+Rw3i+94dvswj21+UD+a9INwjL0g2ynakYeyUunYMbs21Q2xfw
qEj8bPWwDqgTkJFh4/iwPXsipc4DTR0PyNWzMPdQp5ojSpiZ+n0k3jG0lMl+SbOj
wx8MZ6ZiDNIeq0Uf2WwYi5yvOGa/i9AEQ+sh+uo9YQLEtccy/3USlOR1haPfmy65
dk20LqqLCVV0gIZG2A4cZq1lt/kMqIs/Tv3PkN3vrOnUH1HBCWQR0EIGQNtean0c
lfqy79zgnGyo7PIU9p4nqNZ9pDVz2nnHevfgWLuf71l0r8/i5MZurLySvgT4bo6b
TUlEap4HGyl+EtD3igCRzQmmWBBf3FQ9NVrX7MUrePknkhQYgFxitHr6sRmpAQ52
jr0yedEvJCCwYkCzBKrJTwra1t3zkZA85o4VeCLkK1GqdOHcXJyjAet5rar/IEqo
uV8LwuVGJSNHqgENrDl1rOg2J7n6HyNqivNyXZrcrUpFyk92bh2t/VhOtBikrWZW
pBkBy1EgFQYAsBAVggjPBxL2vI3zCevw3lBArlDDLiPCs2TCccXMZ6Rqs6/ds3sA
lPBLEDCz3d4mX+NeYij7oqQ3zOirgenQGhsa/hbK0D1BkeTnNHRHTMEAHxXWfvtQ
mgyqylI2/G6okWWr511Gxeigv/NKBRfcKH1uTu8WjY60WPIB6pCYcLgT1rqRiMtt
qfUDNRyo1p71ks8O5A5ZfSfTglmu2P2TinscZeKE6QixTn015UxOi9NdNauGlbj6
z1Lcqwe/u99Nre7fK6LAgwQ0pALkRBFRrHPAEWzK0jhk7psy/Keq9ofNvt3ndsId
ncy59yKeEYPPtaLgAvw0Q9y4kZqzDnlQWbJeubG2kxB6/oNZwa10f0fiFZr1p6YU
Ow0hSZilMDjFs/Awuvd/rof5zTP3xpkdqUCp2wNiZloTovTEAN1EiQ8rYyWY/cgY
K7GPbxFZ0yNxiFXfMzTM1fR+XuTVhY8LSbSoYNNUUOXBtH+rvXG3LHW77R1pCvTw
z2Jqgcwqp/smQHlNibtk+dFBPbUkzgElHPm277GkGTKw+gArX3BlgwVhGJMJrgEI
sp/G5v4TOEKL9fgEMfeMdOadp4HKqrCWQo7Ed7m+ibtL9W8IyNEjN+dZrVar+Vk+
pcybTWCcBbWD2bWBHaneCc8/0AtnL9k25+SEvFUuhBDovfiwtiax2HKrSb9dOrl+
vDAMdzL5Qvc7ZKOCXKCowo5EkeIFWv56MLQkBmeI5rrYRY7B7MWNOdqwjebx346j
/FCw5z5Ij7gx7XmqEjJqI0rCQFPKgIZLHImyDKJFBTNY6kiWaSC2dJUTQ6/FXB23
tJwGPIX9JbbTrd/COUEpi1DIZw1Ov7p50tLn/uY2SeXW224Waszf8EujLDve78LT
xgZRyvCwvKXDuam3HZAOTrwuWJbE7dMEDCalEh0cIW10z7U/orKDaeQXrpNhS5Wd
tz4p6nwvEw4sU1oiEa3YzifAgTB59fW/rlrPgO3MwTjR11/at44RdaqeWa30ntBb
aEvWxwEGWhaOEBu1z9Jos81w0tHXOsRZyMubwkvy51cAz52mu4kADK+nXnwHCUq5
1X1DjUjsI3lr/17ODQi08FHSlZuNYW9cDAscreHwlgtHiegtKLiQFMfv3tyOPM4A
3k7ADSslnEj3c5RJJqVecV9oYyVQZ0zhQHm0sf3Bzr3vgMM1rwriplUMa4nb7Mve
7Su27LGvHEx5SbKlMKxGXeMODazL8bd7a7mpd7lQgFgu/NKeC+/l/Lw5ZzlFBWC4
dDccpeqvpd8smWrnsC1wgiX/6TO1OVdPxMFFxtNKRksiHHRsSY5DwxrEiDzeBObt
it/Z9ZTnKBm2Vjkxh76DztkoEjP/N+5qoWnGqnK5egO+WwsWvZQlyGvV1XnoEBaj
IMjwiTzKZHXkQYzACr6vQ7rCaIb531HoBR1XeEg9yJ1CuUvjVUayWjA7oEZddztn
x0HyzZ9JLp3LLOoC+jbKX6oB0tUkK2lsSbFVgqQIVndIoSm9Dowld+ntLQjZTtUB
bKM0P+NFpaKWRmDqjAYsDjAuMnUGRhZh3PWo7k98kXsMKNW9WKxFn7iF1rfn2Ts9
KFY7tAgCiPzzC6rDjkVLjRb/yMyuItNoMjYoRzcj9UQ0Ys0cUc7TSDlVK3uBF2YK
rIPOhoLyhpl74Qy97JNFqSNch0UD1qxcujHFLBrenbMblobH4I53eb4Wde5PUc9/
PpYTwOrbQRPQK1x6Y8AMTOvNT5xoMi8UynpahUJ+IHBf/osDkJ82OARjLqwn7Z1s
p7KCGvaHCTVS+bLKLi4pcQjeF2Obh50CgxRuRkNGjtlM5ItXLpICBLIH0SFmHUbv
QESt59y5pvVhpErPjPjtG8SkD91iQOP5l9plZFcVS931Ej4dFQ7hasToS8Mx1NgO
rvLz2LocBmey6+cgwON33HEDsHFZRmvj1O6popv9tuUh3Acca5dfF7zg52LeFV3V
oJkDpZAdG9udlXKS0YWdCDbhaZ74M1pjEZTcPaGzKixLA2V1NjqKPJDEecesKMmN
8HFN8g9OTgv+Ry2GQ2HskUqnM/j9KWYeXkf9XoXWLUXphHd3POZgqbkSpq5lKvB/
eDiy0G/ajBTqHbjpJGk82FYmHafNaKWDIv0G9jAUDJ4X+PruTjq7r25DK0gSXpuw
0XeP2oJm6DK2SFqYP7Hcv8fAW/vesI1m37TMVrUzbrWnSKkO7yD5J8tHEN0EP6W1
6GC44wQkCb65kZ7T8KK2/3j/NfaF6Z2qTrUnwce2boThXmcNvk3O6bwhgnWMukPz
e2l5KkxgEF1/OriQlAkknlDg5FxH0hU3zwh1O3pW1YicfJeHCZyervVag8hMdoDM
jdwvRRDyG5FhRjuTt5xijCmHM5h7HdibvCwsbUgMrqOWla05yFPLRVAU0tWVUhMr
kbK0qTt8mwpEmguTLN8fNyBn8Nzf4QDKUw5hhOCOdl6gKcsIyt9IF+DjmolnJleX
xVcNTogbRGebseTnSkEYVSxW4inZus2IO66UEcnuMS1DBFzx67l9pyOaoegITafr
y7FHFRS5dLjg4i7HOzEpEGpetDXfFZuReHEKWPQcyorQRCneJ0rD0brnd8HKEcCF
G/aMULiy3ld0Tath8pk8l5/uk3nq2B5QvqQVcpYDU6oz/9lFB7Tttw868CneBwtM
A6nIrtKxGmnGJdhZIH5EtptHjknVH0a8pAPLatsA+wGCxqNvDOOYRLZyFNMmZhvf
7FWC+2drmVE+pQ/JDVT5Ia5IBUdr0bmg4BofsEbf+zkJOIKnwgIiEnIrcIeQ0Ut2
d6RvvtawDy+pww/adC8FLF7DHof9G+57XJ/5gvnZVnzY9GU007PfHQaUKuOFlwly
aUAnpYhRSL/xVufozCs5u2zE0YoEr3F6ZGEq+BhJLpeJrrQd2XtqQr0LzzksbCUQ
EiL+3eaoVIshQ1CchoGUeYSB0S34XIZz7V2gm9/PV6Um29CGXbawjGGoubFGDvHF
wprtLnaHX0SC6fC7tdvaN/F/kw3JHWDMgeecTSKyXU5CddW+nFhSj7/YcRYlGElw
VnhgwLrXTBlLW3daG5i6a1WoOOeX6e1NCtI4tkkt3BXpQ8kdDy25jxQHvRNWQGTo
EaoE0gOEwhxrm8/kZ5+OIN3TzTpA9xES1D6/iZpBsoXkY4frb004jy9RAIMKG4mY
EzV2WyLpjR/iVJiHOUlPPZT/fzmyZjF3Rqx/X0MbbdieekNdVGR7e7pnPhug6jRP
DK04yb5rsnODlCxTD9XfGetaeQw9AUtt1quN/tA+B5ZoDeOH4mf7iWnYXQMeXXYd
9TUGQZ6YB65wJD7qlFsoW7+/DPUjNbqtkxnttyZU5pmiDKU69LL5jb/5hO5jtXuy
sAPgrtBgEjW62x+P/gWC29pgnfMbFDKHh3r3qw3Mz0grHAOWrg8eUVKcduxDjtnE
9MNWhXGT0XwT76B+/culARjWrkgWYdsku06+nQwBqsEeZg86iHhqmO5UeaNFyfAN
Ws6xT4IRRniwK1pvxezWVDPadU+Isrg/QA0TSpz4CmdjUY8EehSqgN+Kx3dtzLuc
mXY5EKJBSjGlg3Af44j5sRCPhYRyi/Uno6G5/BjFTo1nIWW9eRNyZ0SGjBy8TW66
LMe7pyoySc407BnRC9jjn4vW+5ZR/eLRqvHBV4QTlEjfJVAm7E4XU/0dMEl6PpsP
L9qklwCBVS88L94ctZwURdZZHTAHQYFhZm5/qmOI4eePyAKd1YU414li+ATWgVJd
4wxf3zjw8JdM1nErKbuRJ1vlgCTmGrTE3TmpgLv+/dVansqYPIqARAGaqMCf0M8F
W1CAlHT4o056irlmjDpdEr5aDADmmIP1CgOMvc3EdCZ+x/lKdA0ZBgkC9nwk8iZe
m6kXcKG4IYS4XhcEnEfjzJw97mv9cHKtAj38JvBS/lPYSljoqH8bGbIhrGIn/cIq
uKr08DL3cC/28/o0lDWNr6Yj7jdV6t3+6gFBKTKd2qfTSTrtiFJXQslplgU/0d7c
fs1zq9YxOXC69XkyA2ypOmJJavnlEMvZfANCJcWDHmWHHvrLYdmld1iX7uOCYjQe
Fxx/Wi78tBfcPXHCBPJKgIBgUELBF62TgqVSWySzdwlLGfBCxAX7mn55q3NwdFqQ
Gj2hybocwu7FtuNnZF+Ii000JczOMabkoye7cUgcYUJeNYXoaK2ev1ZONR/A9qVy
RHjAf2kUKt2uac+KBjbrRau7nvyTW4Pp3pUWriOOqfHdmB3Y7TQfEI28Gpa3I6O4
aRH5lIsLKiPuIiiEbApHbqMrk3uETm9afztBAj7z1Claf7TpM3zIzN1NPJK98dvV
GVNl/JJ2+Qs8FAHv+rBev4rMfakXG+jRGCg5ywdR5k5d6q0/OfjLPr/rMm8AF4ro
i4J2s6yP5L4wGtBwX1pqMVO6VqNgapi1gnrBWu8EsLLT6UI+oJcR6IvQfX8VDXLy
sy+GKDOAhxPhSJpMyV2npRPPWw1my/svcS1CMLcJw8DOf1rLpMRngRnqCcx8SFx5
Fa/lU2du1fD48rdcyoVG3xs1pWrg/8qtk19Wh2Xh/51VLzh0KYS/qbUwvb7whE4O
yE4qBuH7flxQFqdq5oAf6U1Q6wh3dTV8Sdj7GqWua7WyQdxB6kv58T3HrMXCAhOQ
odgvZViBkSaoxWHbhiLcrq1f4IThGVkGlGJM2M8xP13/sJTJcaTHdPjEFdRrcnbC
BsAZLs+kVgcp/JYx02FRkQ7vsnQNirb9AKN5P9jX5xZbDlp6FwDVRmOegBqkA4nV
Zfj1lkT7S61aygWUGsqoH1P5Su+OLBgbyRO4VSxjuTIol/DNvUGY7e4pLNjxxzQ1
xHPR0lF83Zh7ECfeuB9oZsrmARReblw9vkMg8pyteX9bZU1nB2OMn4VBYuhYckIB
NkhgSR4XEJLCaMdt8bbrX0ZV2lQHeFGy2BxDaGK5P33WCBzMjyDBGnJv/uJddBJU
1/vwwp2XOBjswUdEKDVyKBM1dZnpUd2Nydz+5xXS/udUi7rplPBxbi/WFnBgGlun
hdZH4bNANiGPR/WE3hb3efcIjmA2DVEcG6Lrdz1URm1HC6XaMms9Ydh4BS0eFNfX
R8PwKVXKCHeiUKRpHBjpMv0c/ZBj0uBL6D92qobdFgJeS86ShwKk41Xph5d/xz2H
075mz4zJvQGoE9upkFAwq1NkzMLxuEY2FSmCSYEgBAmV+x0SOqTsoCcMv4NL12R/
RQPDLZ4qJYpR/PbetgsY5geNzEdB5vLOjJRiYfJFBBnmjsgpaRWH3AJXD/pxWES3
UkvW0Gcqd78ycpTbT1oCuMlDuhb5HuiyhOubVCy7lnlWD+JrDwBltJQ/hWqn4mX9
RmjRSSSmRHgVrlyP8Vc9l8/nsBzNIVn2I+VXag7rorUV2i6+LFO6/EcQCFXpnWsl
fNuRtiQVGPPRMXoeKd9MpaC0tqv0Z73fnh4yr8cW2x/jian/XIoRPRJoij9OQos2
0bJmGwZgii2pSln8Scf9fzX+RZ2hmLZadEX1BMk7Kul8BQLGwhEVelTe5dhgRIP6
EgE+9L54mm6k7tYaHPrP09LbL6iXRJUEG84RUZByF48Ef5ozGv3etbVfNDtGxnQf
/P4UQSBuyh6G2GocC4JOxKd2K5iwDLq9IoxD6oWXrIF7Ca+g3dpakiy3Rv+ef+Ua
whr0WLiOXIbljK4AEuKhP/fNZUoRl9aA73gVcKIOmWOVZinCtbja8lvUHTNfGD0s
3evcZ3Awd3Qwv5HuzextJdRgv4JF6Yyxx9S2VOvilwuuXr3DgGPt6EJR+GfT+sLN
C3a77t5IFT5aH9/2ZmHOSX3IYNvvorlr2NDAnT8EatT+Z4dAMJ2mhtrp205y8Y0j
/KmVQkMt04W5hRvkAMjV1iYghSSdQILBI8b42W/wnH0YgiPTjQ/bjdiNEVr0vZVJ
qSyYJX5+58FuUwiiLuWTUi4OARDHxx4jpxbxlWrBvpP/0OzKui2AtzkhqYHYnl76
wmg25LB/oKWWZysOn5gGtq2jnuXI8cXZSlqW4+Rdi+ok2NUeBDBdbC8hopv8AAef
HRwFd8Lj9uwXIyweiqjG1L8kaFpKhZzVsd8Q/56irnhxBItwjUsBoMDGTgEIGX7d
V3iYbPdHZu2Mj0vqDeYJYxsYIhlIn4A/uMC0daCNgAQFb0fiz/PxsXMqh4zZ1lVe
jVqOYo61hjnIh3GxgyaELs2QO1df4d/d8aZaJ2Tc3cyHSPdegzxT1TCj6bExODfB
1LOdOvvOd6crGaHdEr7MTdi1FrDxY62ASO4BxWFFTgsOct624bAHk2JLXbEOa/rl
0UGVZATnSfNhCU5/FIDoaeEhMCHlCEO2O47Od85pdfyDdJymWMmYixuaCgj1kk6j
bfT6c8eaRIMQtMY+BpQ/mRnQV9XVkGDrXwLtuIf+Hq7UihQSUvt9pEdQXIT57szd
si2G4sFg9KSai1eWSUxaADLK/bxQuLv6xSj5mkZ+X+822Zlc3JZ4ksKSqDhXfUjK
CKAa8GiL1qIrXbS38lPLyTpiDjJSh7hAk1FdjBV8PxUs0eVjyRmxo7vjIZYR2lVz
mg8gL6HBr1zu77m5GFwcHFiZ3dCNL6dumFd2JnGLttkaVL+s0lGORixkxMFkYV6S
W3IHc36wvC1lHzVHz/8exSwhvDUHY49d5OZa4MyegcrBzW0S/p9g0nvV7/6afk8p
Xdig6YbPX5tEd0N89pxsrwSkYBUjB0nwUVEbWB0ZRC9RcPSVR+VY98T1QCOsLBaj
hMkehKnDTFg4+/QI6gavrkYmHUJh0rLO3EBW52lGK7e+upt5q4H259PgBXzzhzs0
HS1LSXEgdcM2lj+/Xe8gJhWYVIvck6bapjv2yE+ucZMerxtRHv4gq9rBtvALWCpn
rEbYX3ULK8Xd+ekyolArL3yOnt0sXl/Z9mYA9nuTirshlcSGpewhtPD2dVRP6G4R
c6g5PDgOdyF/1iPNaTuRy3VtCHd2sPO2yifJh+vp35wvlL/70ApGBqmPHCHHT8QD
u4lAEFfuAVeGL+lKDvkPnR6G4wbzGvHrlEqmzByMOTE7tquRtj9EJQigs+C+R67a
79oDHeek4bTEUfcLjVK/adgWX+73r2twd70nI/u4Rt50++E6bbZ4PybEEmZkUfWl
8KWQI7kcfOjQXAetpi6q8czpnP/GZUUxXsluoFbSbazPrLUqy11m4YnF+PV7az0T
MRR+g5Eqz7+blOmXyXG6yb5CCWPUOy0TKCdWsFVPHghEOYOO8kj+xgx+jyZDaC35
pOZTdbTviG8lqfZboa1Wi+CSvWNcUKaWd3rektn/1Nz/nr9Niw2G1yd9QDxiFhmz
OKQ4z6kRMfuy0g30PsDRmGQLpKyKmFiKUiO3ghEKDTDl+Wff3/uuTrUS9MOO01wJ
SmmHrlcdvFPFpRejSaW7zUHseqq+E/m95v28rE+y408f5EjMLAuITIAvchFlk8/V
MV4d1j386R4jNzBAWF9+EfvLy+X9oQfjIpDnbGUJduSLRAuZhPbM24KXz2UaHPfp
ruL6DD6ENR2cHlJuC57WJJLJeOTdkeOKS1KTsla+bQTLCuIsPtcbDM0ZcDIMRNNl
le+H0vaLx2Hbwa73O/SWtcDF1PFeSZ3QA4nJybD9hAY13B4gIhKnCTPdJMqQbewz
eriUQQZsEMJrsG4N1WhWPGbK/bkegO1EEfbq8q0/yIAkmoJWNKCyiWyItcxMi/gC
MZTyV0sgd8+T6lw5f+BcOPrownXOrGAcGa3YMa47pyGT6oU6bmAZpWIzTyDYXdoK
R4gW/1pQN4xNKbaa0xnTHlw04wgByVLNHssejONjoHaTII3NBKRKilrpUWd4AObL
4krSaNb1r2Iim/7pqaFe7sP/Wl4v9HIt1xTY/GHleMCgqnSfmQ2o/ZBNPYBT2bV6
cHtiHmGVpsXy06k0UjEONg4G1Y1SRIRjfGp3cLftQTIHZ0uK7+Ka5W2Opn1hs9Ro
oXidsJ3L95D4VynEhIR6YCpv08NdXDoAyDbLG3Jm3mhj3tuRAifejJVs2uK5DhW0
oi+YSN99GOduQ8r0WL/KBc6xEtu5cSzCcPJ88H7fIGiL765w1HAIrKx6Owgo2PrT
SExK+CARUQWDoHL8G/CLXc0d3XQPQYnCSVtnUXU21tHw4e/iM90U/HEFEH5X+0E2
biZdvWjhUWxtxC2WOulI9jxD8Z0+cn/IxcAhYhwbky204vz5ehwrTUc7LQsmGSiV
R4h7/RtYabjdxRLmSt0h/OD1obAW/EUh7s0jlMsPw5xPgJ3+w8S/EYIjmRYI1LI9
6OCrK9NMX8b/neUFmi+4kMTG3oR5hWm4oNaDnWUfJRaaaACRBR/5mfWEH6hHfvm2
O9Y1rhcGfZcKhnbBMmOisUeJSUXQRdY2x1kq91Zou9ImxtM0OFT1UWD4rluSCsQD
xIOAb2PqGB260KCzgTqu8zQJtj9Vu4PduwTcozQWOaK/qSq7PzR/tqKOTRfgqy3o
mZ9aOfHi3pQBgnR+4USU/mzYsAbD5LfaaHiHsuiDhJyOfl9gm/kfo2Ra+a29zaLf
0LagYiCfRTOMdx5CsuhuyBpqENppxZ6N2HO1J4TNdMnZ15hxQD93tJOii/DXJNjL
JrlC0BzkewUPj1lC+tBBGad8qMD/3ECBMa6FmLpktRd0U2DIoeJmE6VgwBtrY0WJ
NlRN+GygYA7V3SF1p7z3pA0HhzZf0ujSegW9dbwMn/GcN0SkqPYY1A/V2XJC3TeI
73/vRWptZ1IBWMITl1+jrzUstKSvNv0pvLyWBwP0L1ov3P1oVzpPSR4DHpX5Qs8Y
c6zp2eLFHhreOAcwDyHHNSWxY1dDGzsCN8uXv+L6LOGfCYpDuaVi7kOBS+BO7rcp
qVOEoa7biz7FYcctI+RgxLvzIrfigGfJsXm90qn741KQAyuh3lVUbTtUWSDoYm8h
JT6aBi21Mh07zaBqLJ4MQgP31qpQznBba8FaUkPb3xAitIln7BhEldpzk6x5vShT
4yNv0Ua5LXEmsvyDx1tQ1siJTCswIC5hHHb/zPky3k2YoOGOq2ViBvIMUF7LLI9R
15WvkZyygbP7ocERSTbOlQSons4JWvARQOf3eiIi+TonW4mgNfukA/i4xUXtDFqp
1WuL8JD4MImu5wp8w3d3yk8kbw9TkFIAFq7pvLr1pPmOTlQKwr1xsuUVLKP/Z3Ms
G+mn6WK8wKcKEoh5kwXZx95CPZPzdHVIIK54ny2QVGMFUAot67Dv7ZzkfTsum6yO
nKZRPr3ngCqRBmAYNZF5/NfzZLn86PGPqvWR9cx88WyTR+5et7M3SSDf+DQx0JlP
SafCMxSCv6yWz63v6lAl5vcv1kzSeOXL9fzVC3l5ZVvNuXlmKrFcqBWkd/PPS9Nw
XB7evwEkbaNaxGfH85rLT+mDmNq7CR3eIzvryC5LwaJ3phiYcTCaR9uDLlOmRnBs
f8ulZhJmWktYbv9HF6ky4FCsZ43qOvQURwHHMuv8TQh8+6Syv4mdU3ira31exO1E
L+1RGcBdJaq+bL2EsPBY6jh/lDneXYKSBvohv90xZf178FbVC9OUjo7BEAMHMVWG
DgpmbNrr9Idezltcjnd1nAzluZZiWYJ4aGZxU+Z2Cw6vUTfEgtCiyrH9Qvmg2Rbl
hQKWn6Orj4ioArLWyY3MAcbduAR4q/2XzCG/xaAHVj13ZJP9doCdM3L3KiCQjGjj
aMLYF/v0cV5cnSIN4R2CPau8osa7zq2ezbU1OVOaKfgz9HZxpTK8Kxt+bkRJ5ms9
jYTqejk/Qna1bVG0wuEHedN0e7Hqu2o002ByQ/YYOLY9Zy/q/Ht6ghvb4Yu4Tjt+
bbiMXv/F7F6mN6SM7wg5G7rw40W6w/VOQPyYOHNWGvZWNv+lIQWuXpopNdH+fTY4
fXSpu/x4xC6DPyxe6tjMGFEC+/m6M34RnVQ+vSXd3XtnBvEupJbsLlx9kS7M+j09
1O0GpUKmIQi/jSp6qLS+iPdBYgc2OeARBoZpTakXABIHx9yLVXormIMA7+aYaznt
hZdz2pyoAvOrSiTf3bDe+wm3EY2GzEPCB6RIiAZyCxyT2rmmqWapxfCLev6tPiyp
2+U3wFHl/nPkWdvXFZRU7yyca2o8HVOlB/tK2o89pg2E2jLaj4WsCZ9rNVz/c1y+
nsPfKYZoUSl1PDsnOYNFn5DR7tcW3c+x0XIKi0MH0kLs60+dBNrB4UzeQlHWDb9w
KhtT1u4jM0+79fV4Ckjst03EYcMZRYdT4ByssoBaOIxCA+b8ek47AoVHYAADfitW
TEBTiNDrZhgdgjjKl4qKVOlupHSF0S9aqx9AEkpSQZ+hMKGG2gwc/p9MAqmmOe4Q
7HYzxliILf4BQzIDukG/JVVZL5DhTYWUV2C/vAI/6tV6eShaxC/C8J6SalWH/OAa
HK6o2GFk9JBD9s/tR3sHfwr72Po+moPBYjGbIxoIKgO1Z2/L+Lr0sUinfFm50qos
FWnTCFI8cCsEqj6cvQkm+ZvA38chFGFqyFY+8vD/3Ab4YIa0FAyxbr1IoKYiHWT5
fkvPZjOHV8YJ0Luc8na62WIwU+npWo7Xbq8LO2VqNnZbGFazqhE7wrDJvkxqQb7B
9677eaenmSuZKGCqrOzzOy1lK0OP1VSSj5ywz//BIC/ZrQn1DuFoGfa4hFv1tgpk
jddb82TshhXmQ24N8nKqdaeah4ZUTK+6Wi312XcUWSTKVovcCZxqUTONHFkvrM5a
OimgncsE80u6GR+nVdAB92x0BzTGkef4b3GD0QGVy6+Csp57JeGt/V5aEEfpOipe
4YI/93v6Tmz7cIXjx3Wxyl3ra3CmQgPytzFWLUHyTmVzpbZ59uPYpcec13zLdvZW
qhIGSESfJbUTYqWX4+M1/LvtZIJ4F6QsX3d/284Mvav+lJGm992+alJ2/RJ5mB9d
c+kW7uVDcaLZeR6/sz0kUgPU5+KkGSqzb4hO2uw4tvPNzn34NVXu4w3cET+Cf7gG
rx0pRWn/3oz//Fsp0juYyC+mLPdtwwugTomSTPJ0OsLNzXo37a6eI1Biww99B6nK
t1vnaLd4epzczoUG1LAzR+lEG4/YvH7Hl3Oqc9djDMil2eP2XlFGfYLvBgMH95GA
6sSWKZVCyRh9mYhQULoIyXNEOV6OzpWh9pLDkwjw4xDt2TCy70MKdym4zFGBeiFa
EsIgH1FmWuNyk0wumxx+guU/PcqF0WTGFqGoAFiwMFngeL7awTZjWecGE844utb+
gmAlXHrGObiupJTnpX2vNonrwlqaa8P1Dp2CMF9jlRf0yeWgJ9uD9Q8JohPF8VXD
l7BuN1ktvo04xPe9TY2AsoRjRVNAgo4M1YktURlGv1rGm0fwucI046xWhI0HliCk
bXmNfdBLZK1eVFw0aeyUgTlTEt1uQZy5aRPVRuGn0P16FmwUOX+Jcl17vBxm4Wdc
6UakdlyI0ut/Pe8POIlGQFxqyKMCrud+AN4H+xM2I+KAijrh1Lmc9k03I+6z/JVi
f63B3vlwL/T8Gt2LYUyJCB4XNmYE7cP3Fsqtdr6C75fyRilNTjS28wKGmneRI0iA
7sbWzn3P0tjmxVGlQsUVzp77o9ZAXcuqd7hKvP11pqLs21xLSJC0MHxAeUKQGRe5
Wl8jEPmqSQxv2KG4RyCHz1NGvOTVVtPrHlzqQVvdXlLGtZ5yQA1M0ULeTymjDIy2
ApvVacrLZsx6aSAxRGmDcRAFjvrXOhQuqvTBR9TdiD/vLdHaAg6QNPSpkDNV5GIM
mEoZDCuMksEs/rlhJDHsBDi+k7tMkUB8A9DiX1nySDGkcASrHCoE6LQ+BPkcA35L
pJLUbNgUcenHO8fejvbW7R4xfUMtRxklWi83IYBQvD6KDvNP7jRewfnl/PqZsk9A
QdaO2If6tXH6iqIxIw8TqPkEp2HsXy0x/08rr4d5lcXHG6g3cmifyF1OxhEJj4Lv
Cdl1kVRxpgaoRK+M9DiAn5Xa5roeMn7issnxH7ZnLTBZXhqz4FAzXQNOjTxQr4PQ
C3s14XU6NNwOCdvvrGTYefr1jB47tDo7NYsaMTzyt3tXJYRNLsMbLMZDlE6qQ5Ca
2aZykhn/UmafTtDk+FTNjhemx51MgoMzp2divOy/2XSOTzrfFLFpOJNLihaIdUCL
oKhahshgT/3e9+V+cOgdL831pDgZ79EMbi+7rZr6KlYv1mPYk23mxTWVbSZlauKX
GOlHUehx6eLtQGJkvdGStlRCUNRn9Y/hiXlKtl+dsec5FHEu87Kj+3QC2H/Q6Gqj
3DyZiGNA9AqFTH0JW8leEXFlvoQ+xi+eDg6wZ3i/wJnAJO/5HvDgbkHP25HDkcS1
25bT3pnV7m5TpNY3egNS7SecS9QYkLpIY38M5xGZJoTgcRE0N2rwAH3hYbct2Hjd
tBZugQRWGX8HHnZdzZ8mJA2ugIbwfGIBigXr4VkX4ISC8TSKVvPi/oqw/tweVnmc
+Ij+6jxcAccBpS0dGAgHctiSxbfVT4kZU4yOG2+hRwId8cRAj5DXTo14UeeBMaxN
h+LX+D48OvKgHgOFaiVLLF1pLCekH6mTl8yW8dGpjjKQdJErmU4KsDOPjtS/97bo
UAwJ9jMFSG6gm+rYzCfllDHSwcPj23eRZjlBXoC1+wpUtEo0csLrq2W43kKmv5Wr
qb4OQpM/7K8XhVg9koSXEJFpnclElyp0HvDGXeH5WAoZKn+FGcVI4FzFQZ4227Bc
0GrSOgWZRwawOivY49lXD8AwmpfocE+IobXXFpjfldMK5dvp7o/QJn28xY27SdCU
9LJITddTBCfCnBakCU0T0GNfeWzaWKgWrAga4qMQRiziTbaD3dWclorRW6uCNz4M
DbHrGjcDIJYzOo4S/Al+KCDWADZ/T5UoMC51ME/t69FL9Yl0PPWY4dLFOEXoZ+1T
ZuhEZKi16flGk33bdLDe2k6oZNN7AZmS6T4ljjqL+02EJgopyxY5jp4d/llvRiRN
Zrnox6eN5JFCABiOvtaYvQZK1LG11FEatN1U5jEOBSgvKJNFI+ygUvE9Y5kD/pqa
ICQ9G9H5W/wpsnQ2u7HZQVb+Jh0/DIuApJLEs49I3oRrmi1gARbZfHbGT4euQI4m
dR2aT8XZv+ZgwBvQI+h2L8F9ER0HKnfNdB2zTw9PS41f21sQPzEyDht2q2Ri7LOm
FNsysvwwkc9jDat8kgQPwS2unSQTTiliGCODNWVhwF5gNK2iA+qRVUY8FC+jWJZt
lIL4UGZgapBPvUwf7n7NT3gF/wWDUN8OEM0Z1tn414/hmEvGlOe9vm3hNiW1j3Rg
5ELo/NeRQson59sZy9cw+HM6mWes7KfNu4glawiQya3jPseuGC1T1Gaz3yMyZX4/
JEI05CjuRc/7J7Na48jO+ZiJ/iuMfOLWsTO2H7FL077NTHrGvH2mCbjBK6ZGdLUv
HfGU5CgekNKvrn7Ac7o/QcT7kcvcMpwdPCMWqz9wu47UrpA/ytMVe9vrC4sWYsaf
RKqP8uhH6ADyIt5xfVvw4NPGffCrVYZZXIy/f6CsEXrJczQ5OZuPGJ7ONiEFJ/Xf
iIEpGSHEdEuPU6mapCukk9goKyOoFI6hZykY4RYEl2+XsOyYfWDpoB+wb6xKWSxg
9rMIjqDQzeUwDlvBh0t8jpskBcLBmOG7HMhR6HDSud8qqKpZ/dd/FyTGw9+soqAw
2gGYQUPxom52S08H0h7wzGKH+JrFIoFUQnCKBtqMU6clVebgzvfA+pdDzpFMQWXJ
hOKBhAOiH80CRxl359M6QDI3tdwa2mXD/lbZQ+oEaG5vsUrxVs/4C3I2Ov3jKtJA
Iz3rL3qebniXSG/4XOWnD1e/W/Gmmu3MJ2SLX/0RNRgnmo36mdv3i7trWCVcSujh
1LnKPnTw5Fs9cI+XTg9GQhAQA2i/6f8teHJHs/TPje1H6WZHM3WLi3R9Dvl21OVa
M7NtZGWz74/p3v+4JdczAFIDGdIx9E6R0n+6TDts1oPrOxq9w8mar04AnJANFU9/
HkzIRXo4e8CZxnooizDtA3FEJz/ZdlL0UI9ZvWAW0OPgKlmDWm8B5SQtc7ygv5Fd
0fFPhb+XaZMVgdIN+04Pd6TB0wstrvRcqZD5TojGS5ZbQydfn8lL8fZ7EarEJf4+
jebABbik3JcNbCJi5Zv1vlzSc+3X26CpuJ+X5C/cDZ/6hWrvOSy8nMDo+PlWLzog
gijt99voSGnjAr64awueWQqkiBh6DKzKx5kvsfztZuVf4ULbVOdQVfvanr+ytboX
Uxa7x786ITmvEfuvn6uOl3whbMHkTcUuGDmsUJPzEBswYezbMXITXUxghlaX9nJB
qoftrU9o89mxr3l9cZQwoffdb3O6fD8/p4HFb9SIjDOLIFsB1fIL2+VVlIcue3Sm
BFKi1oeEZutH6jOmNKGHPzR9myHdPE1A0SEuO0PHF6dzM1y4XciFdDaOEfB0UZ1C
XVmG4h6FPOuHQGbOH1DK++OD5WkluCS+5VXvSloFujG0I6b36RvVnIBfbXbEMGBE
c1nTSpeh4fPHzaT3ZkFVYvDHmLD25aoTgrk4OzBXfJJEWi/wa9miXMc5+YXi0U09
WTQ0MftwoK5WbbhT+ZHdVioSlQt51xeYxilVgAjJSaHvqOZNpAJuW85AonK35xJm
TOVPOtPlyaS3Q65L5BfSZ+gih9DzODoAEbfYgvWxLLca8l8wkgUNntG8D/QVH5c1
xkOEJNr8ZuHTKMW9F7Bt8JhGTmDwvd5O8YtNVESy3/BKwnWpdmzNN3v1pLsZm0LU
nZYIfxn9eVuVe3NOUIQXK2T1Zsjl6E8Ua872nHNAJrekiEiCkIagqeAQdg4iP3Se
tme1PtG/q3faKlr6iE+qkKQMrPUwIcKulEgn7EhmEA1g5DnB4AqarxoY3Mk9A+G6
ibgWykM2PeeXDVJjUcamVSSBl8vJywzaN3jOMvybxCe4bR93ohu7zkHyBoE7PaSv
YLLHrs5X5bq7gkWsoCXFY/lWh/+1MAZTNmFeNXvbzEqjwKGBC5UMhLGHsw96auZV
ZdvhlSwvHAWqi3E8VXcfEd24wQlwx3hkl+6SZIMY6qDeirt8dd+6PlCkq5orcpSB
kiME6NVtFv+87DjBksjvcxhywhQM2kqLxHaraT0pQvoYRfR4ukyX1flaLKFXgzFO
U/lBzyPhSYGCnsZjWKRCpXp3phSqQxuKT/3ZDG0XhqEICCOTI5TBtWRvn5kReihg
W4cvGE1oxe1QYRdd2rYChZfi17BO8zkv1gnk7bMxLtvVpiEnz/yfN2nrJRNRoxde
jGe3MpCSNQizPh+xkqTgKdKWVk6q8h2YA/9XOhhLvNFuYPNG6kMqZTlb7cISDSUs
s/KtQNv+a5h2mk4ZnNXVTLzpKr2W26V/OGzDKd/ZwbY0NgWMnYyNWbzSdf5ol583
jUJKGGkvxSw1ScWHR8O1yHSCIm24oaAisiarT7OdAfaRYISanLmGNURb4NrbTIPm
PMpD3xPn6J0armVAUOSG7CkDaIoxg0eKszdcePxDhv93JFL8ogrX6xRc5zuN47S6
68nhsyuobnFmeRdhzpvIaYXQAWnqMyKcAuyiJd1O79RulK89NmrdB7u9gd18iUuJ
EM/FxrQkE12ZyzYHWEjRv/pDb3Up02YMbW07dv0B2/z8oQE+eDWh3CgM77HfVuip
4efv4JbEhJZ9Vgthv9nGIquiWp+YsMw/jMMPQrikB2Cyah34qFBh+ylfE2qHI0xw
ipVtnOPWmDqiadXOqNx1HrS778o+pYCBrQIpZd0MmRy4Xp2uV2MWcCEUEuklSRgv
v+xfP91eivO2pA/9UmHyIQRXI+2TISvaK2WFHOG1hYub6/AfCtLsd3Tc8hHRyjgf
hR0RhAlrG5dy/UUFCeQvzjHa1yK/tjRhv36I3CSsr5ly5gA29RGKh9VGhxij31bq
C6DQBXHzjlz/XHv5QZq/hsQ4xuyBh6NORXiPhdjU2bEWyLhl9z6Y8fLixFwKIzQY
2rlnSnq2auOn74r8FvvDFmrB4439L5wvfyGAX5F2ObeP1MVy/JOzlXMuRMSMDqRp
/lOK9hrK0EzzJWqddqXK4eP02IUvQ7Y1d4pamojctYSBNGkRLeLWqZLC7DhB14my
GrcPIS7n/1rnTIXSQ79rdLaV9n3KfeNRhJfq4X6QrmReFqEMwS3jfQG5Ew1vU1ii
oREuuTIq5XqTl9IZexBqCBYivWs4B7DtILOayQZfnRB5LSxWtKJ7jg4s3Lqb5DEf
4B+/tqYDAV/YOl8Ud/Blr5l7W8M0Ydo+7n9dHuCg5jybFqB/em9Al33OxXwS2oZ8
YfKuOacrK+7JqGQDjrg6JpziQnqwkoaiDIQLDZq9poIX916LH64tgXXUM3Z3mi2g
m6sc4JEMNd5euKDl4XwLeK5ZoDVleaTF/AGJIt2IfMnkv6CrpOKehtTuKuWsOvYy
gPKawBqglcn+sdU2fJQLKo34CN1Q5h8o8RLsA+jQLa06/OOHJP6L5bWks1TGWHuL
pXb5h/aeOZlgq6MQfH6LnbP9PyrzO2VxdsKRZh9EDfldim85umw90bEPlvaXDOV2
rGeoOioGrHjI3OpkVL2b/qErKa69pGMsZYxqYt6yGRKBORZAYdFIF8lH6olxygSk
U843anwUTXQXvrdHsXN8quCG4BrwW8yQHMBxkElejvgyrb0/cmUp2y51ToyA3KMZ
a2eXbSurVcfprmWypPijAjXvm9jhEoLNsgUUnCHoxMczRl/MS8CxLxGKb4e0Y77k
i9TgL1vCNg06Vc2cBTNcd5UBJIRKogr1PwjLMd3IOWIx/WPUiYGRhVhnixgBFgIm
fZkjQeEIKPjFk77mZT5liVxoTWzVeVGQs1qJJoz2FJbQac1pY6rWQFR0SC7N5eCp
CrUhBHviVWSMPH+Mk2hB4bt6EBKbup4vXpeAs8z93EO2VREmzHlmZhf2RpPdadtc
27SafcYmez6tqdChVSxWsoLy1biEmJdLEZ+K2CUjR6qEk6z0cZ6Pe5p5WZiUAbGu
qs+hJ0UnNDuA8F8KlEEThSWipwi6xYw32RpdfYhMQeSMdgfoEjo5CQWlPEjZ6jdb
wxsrJtE99KdSxiseFOeGOA99dWG74vfVCdu1pbyxWoDCkyfV7y1PuDjwuPNLBVP6
ozcxoeAUWJfCLbppyzSX+1U19VvtMglClYbYMhrB8fPWTZaNENd7w5964tTqmzv4
n2EtrxDAKh0VYVdrkeBMsinkcaV1iRwwF4UKbVc8bAWITND2mK5qqpAyRHZj1gED
TTHDMWkE9jpl7VukbZziV+mk8D9WHGYjXZvpgaHTlI5NxHG4YQY7k2btlBSCzer+
ubAgvFmfhG7UTbYXsR1+uFphXsvLnIEcUlRg1miAtolsxQxPfem9SM5++UV6r6yP
4+REg4C54ZH6yHPPRfYlziBa82831S4oonLzVUitp6qvYQXjf4VFwExDETjmkZc2
AyFzvB/7+PscF0uPgIG310+Nfp33qzhp3jsziQj7enqdx1UEV51hR86xsbZUhgrB
U1Q9oioXIFENX1uMdbWZVGsz3qcxneIaTnh0zCA7sEP7DSKHh7aZ8pj3znlVcwwK
Ja7szNhl6t04b4N4szv5/dAhtuQHrYSs1YDPzuBCd0AeXrvdezlIhTC0HmIgAobk
QjHifUk/vbvRttLpxWXx6IozqZRxtuBH9NIW/z6c0TJg0xtKuSAQGJIqDzuIL++0
KERmblHcapxIZD0lTAkHTus8qnhSh3Z0Jfh0axIYgaM91ousXYCIURgAs2QeK9Sm
VN5caZfTQk4RdET9RnH3GRg9ogTypmviASId51CZ6hOmSBXFJHN/CZ1f3imvtYL2
zKbrrm2EffDgeJtDTv4GgyXm7mg50Jht16lFMjDwnNHacEiT2JZ8BxLpemBisQEu
AJDrYDaQh25egAv9Ij12luxrXMHSnuHOI985MhGFFuBVW/Gs72ChzVHG5l2TJ3lY
jMWhxnFyehvlWIkavl4GJmWw9xnYfgBHxpXdxsU6zxd0NW6p0R3cmTcH/4g370aD
WyQO0HhCQ2rkBx7/aM9Ydlq6gysEU2ZcCCzON60RH2VUO4epqcAc9jQYuDIZilZ6
zXpZ7wjSwZjGdTFfgenVx96gk03NxzbC254ONXsCrnhsK/72BQj7wIOL8R3R7QnZ
JbnqZLFtWmR04tGeqLNrRxP6Q1k01cXjsHLU7SSZT8/XD1yoogh6xb1zItUDxchk
z3MFN/yaPfPFwVMIc7CKmuH3k03ZLDgmeqyj8XhsK/PNi4jH+sKOqFdSaTjEll5M
IMr2YKxqqMP30qJ32PdGMK/14AHg4mzvJ6Cao/JynJeaL8XKSR4aIT/S+Zzja4ka
reD8GDmbeGTn3K117GWPNc3I6s5Hfs5JH+VoxOpRgZnVtF32fMu4s18uKUb81pnn
X6Pt3a6AJofTeIdwbJqD3DpbcHm1khSOkFolxugCyak9/bpYCb5DxTeokjhVM6zO
JIDDs5xdNjVgigrOlwyx1pQwuMk7ZFJp77DCloE/0Upzsbm3vbmGZZWwxhpnUZnZ
m8ErOPGvkjAoGaIIJYvoB+y90GYUswU10LoRgNSceNPIdYNNevb1dOf4TEvlkPbi
hcawDajBF7Tk6VUAUwftKnokF8ZamBdjrIL9XccAV8DvbIIRjrJpt5MRsvnXCZfh
GqkWh22QNKFdjF5qjE4DCz2vXWqGRg3CnSip5PF3TFgUmuZAIBdtMb4N8fqYg5fN
KMUOgYl60K1VUAoGfjclvHYHx1xhsgH/kvm/2zT3lfry2mDfSEBFm9HO+MQnU9b0
bvJze0zmbBnSavvjppVtCQoPkIDXyXqCRsfv3r4S+nIXz2wctLeeVvdDUPLziG+l
BYNFlxliT14v3Hub9SQwlIvvsow19V1wNJREOGnriRq5m14i4Cjol1zoMnVrKYbD
7wUuFG+3CvTOkmwTD3iTZq959PQlN9FUxT3TE0J8YyUsb6qudEIIJ2sTMCg2n9J+
o6/6mx5mJvQtvrZGLA5SzK8rIGffFFB8PnjhXODLLx5VkJTvKPqwTSALsqu+gkLp
s+1geUzhBSulp5ikjEk6xPPi4VT143E67XVBI5VPdnfcoYR0hf4uS2t9vyk6Xnqp
CnZtYuwU4zyEaTcHdNdvtsXHZUCVOH3Y3DruohEaJc/uEM7ycrHjskwniMp/jPng
qKEQx873/LLOqt1QCOH7o8roUn+1o5uIq/lTk0OF8yqyA+1WgCpXxhLtFF9d1+1K
TReC8b/iAjlpEPeOoE4Aq03kQ/DxI+KsW5V6rctBnKJ7x5ttsHFNsmPpqZlQTOE7
C+F+IF9MBlISJR39S9dwnxRCg/1moaYkO+iLCtEerI+lxMsCGb+NiIYUJJT0/aYI
fodva1sL3htZJciOhd4+pPx5IyIJG5pM2IcymEhz9ORQMQiudhI2CmiXHE0Q4nqT
6CfBZ3erbb8LorL9FycI8Bjggt1U64/LjIWuWPN8fRT0QqFa5p6gO36+1wcx62jf
C5G9ZIkWuql6EdFl+jeiM0zcmRaPuVYL+1kVrWNaaQ4AstMH5m+jmkcUIGOwdewl
8vDnQ1Df2nXAcLAl2Ao1Xmk7f7Ys4+A4d649SPdzUavxC6TfnEorvq8vH/LN1ejf
34HYl43zjSR9gYIIBdBUhys6SPa6bn8fKFgrEf7VhXKt73s5E/0+FnQjfE6k40Z8
1Y33IjYOwPWkmTbWsFbRI+eydP4yc1mLZlbXjSr2k8cyzvsM1XdKa/ndXsvsqRTX
w+BpffqzFu1oBX/PxmWnAivYeR4+A4c0XCsZE89TS7fWEJgYB4cz0rC7Qc8uuq12
Fl1VATwsB0PZTVqQHIszU8gkc8CB9ITGEqMiE6McEQndELBgT/dgMBgEs2WmHkZw
Enwzl4miv59cOwUmQL4VkS4vS4PrLGDeTQJ+xcrAh3nhPJ1zEEVEBIr1oXoFwBLW
rgfSpiWS613wZVzyTmNr59KETf1DF0wZeta/sZHf5fjmmhOOg3/s9nPjgWZpGucw
h+nQvqQeWW01xHPBMz3kox6Mfd9H+jqC+5c4lcK4KPdo+00N60128rrFT7ys+puj
9/mMHdax5b4Mv3bdN1hy9hc+ruJB5JzrChHx/HLSY5q71m/2lKiq1ltHil0llVne
IOj/pyLDtf0WteU86y58KaROZP/ewlh/cRM7Hsk9cO+1fuaTDCrm9Vd2w7oEmCLl
8t34V8r9BdntU62qthY6QZj8w/HDE10wJusVnE13Ni7By8FUWb2xn1NNA2ZT0y2E
cEZECUO53ntzIArLJ7Bvm6dWW0Pkb3mbDvOTeKs1gQ1NKR1xkRMQ47a4BMD6U6jx
aJyzBUaDg3HnCfoP/dStqyaPeWXqRbCJZ0vJpKoId4YRJ4GBWBzR/S7H2oK+TRfo
NHvZoZTbKkp0Q6JEKGEmD8RrPNnUlgM+vXnRei1smlQKEt+roJDI4sMCkAt/hFeZ
Oc04DZJNcUdE/Oc93Jryt5yEDEA97kJMB8OAAyhC2qujhFGUThWYQ2ZvTJfgtzqm
QfIU+QCxgOSdy0eY+kH/JrnHX4AAcczrr2dWnLX/UBYd/Jbqtynq6MZ61w/xXgW6
C1rGlzHN+OSpmdC7k36vnr5jBOnKGIJB5G4femD6cqpltCZau/4EgKZwsIeYU/Kl
N3yL7D12WbH3QvST9Y2MjaPZDnybRdIYbJmwcqzip9H3AR934Qy8uuRJ5UNWLw30
X9cSj8Zat0r911s/v8aT120W3ptXvVcRA1h0LA5gggtSeEAro5OKdiReyz/KcxdT
nDKQLlV9nwg3Rw+s4FwS/pG/3Uxy5rU4eBFoQLYs28rRfWOlzYreqpteMtwcHUiq
ZInCWC/Wh36P1Zipv/rMA3ufgMtJtB5vLF80yNQE6jhnAaWZxzx8+J8v6YCrFIIu
zHWn5LW8Y533WAR/73sjAQznaQnNr+FD1pXplbv+UZPtFUna6EoVlsS9IDssknLz
e1Ef54s/YzzsGnn9S0pp3XHQcm7VQhNCdn8otMjE8/ODiq3Orsm2iDimi3giOAjD
yoctbO+HV5BqcO2yGfwNiu7NZKJieTVW5zNibt0upfZu50wfkK85g/xsMWhlqks5
s/eTc9tOVzJ+7qhrj/xW8JaUB0iF7HeElA5H8ncl6623khrYke1LkqpJavdRhCvp
E1Rz4dOf6TOIUUSiUURd3LmS3lhAX/v5MCYV9L1pnZPNSOTObGFy8YyMMBO8m/Hy
nUlsniaByu5w3lU8QWK8PufTAVnjjPpoYnnc9wROc+0jNBjBMwI28XAVeOwbqiy1
H3uRsUR7KmaeEUhLO7f94AgRhxPx4CK3TqLmlkN55NjeXJuWWW5iBhRje8vve1iI
fWnp18MhuTDjqxJp16FtZNu0NXw9hkAGMOmAyfUDl+gnIEdSPjaCJgrifnNg3ifh
QnqaqGVyBiorvUft3gYpn10Vl9M07Dd/Lu7CU2ZF8Mrkzd8/hPIG/rYSxflApUlb
wAdXLEU4S5IhfZPuS6SJAtj7oUeSRwG1DG9ZsGRth37f5q+SgqgXOFlPfmGdU/M+
glm2lJyIQpW9+749G7QeE5Sa7RY7FXqg5ji8ZTC5yP1i3/soKbUt1tWUYGQGxNqC
l9S19p7orfKKJzywbtS2NF6WONdJWY0XHsP3CeA/v/IggjA0iNBy5QsZ+FzQJRD4
DQAtWi+juPesIOYLdUUV3GVxj6NzWcO7sIxOXD5dvy/zShdU4Czvdq6Bp2xIdyfy
V8eVwl0la+F13tLlVJOE+Us84UUrPkic3FukktAoaAVJ+jfbcKqDXwcInC6zUeW9
oveIpbh7kE8W6piPe98tqgNgsSleYwi9HtfhmAlRbeFby9tSyCODMOlMF2lYP0Jm
gYSgBq2+F8mvfYVEmxnl7UDD+ObzARKvlbe8ykPKTUN5tC57ibUbU7SHwNq/ljzm
JASKyVKKiNlFj+MpMqrbwIDWPO3+WSnvzdeLDmHNVxEV457nvlDWu0IKVM7VKXQo
RevXM8XuoAD6sTAAINjTAXDb6Afxjz+pu5RjOlK/bCj3UwBvFDeQa3v17hA0bzc6
fUwMqh/Xc9w4yw41O4tLwlb2A8CIBFlOj1TOj7WJDn3QkYayMqcA6UXR5PiozdaT
i1Vhj3XUPobfJPH57cOU+4/cjFoSey7SCL0yTstFYXbaWKeauIMcCjU1sQ7g3LpC
gwpDePb4IG5QihAnmWCI9HGJCvzBQbKv4jhqrG5KoMqp36UMoXe/Yu6CYTFVxG80
bmU9uLzRoEz77NxbrT4kYNzEiCcuuP4rEwPckvqe+CJZL8uY9h/6Uv2TYtrETujZ
8LE5c6nxFivQx1dueAK1/D4PLB6b91KUPyYTZBi/XTBcmqDJqfhl5k1SLAxXmTz7
weKySTgmDlcRxapXZTD56+HubPmk+B5Ak7CbhujkN3luRpEc8P4/M2lgzOq9uISH
H1/1oMNMJ0p88ALo90aMq4m4DncGyWZOIq5K7WmMG22rXyIHiUmWljZoWUwpC8cj
o2705zTAfV/D2fZ7scTqsrh2njp9zfaYAFb5bf4SNPTr8RFP38Oj07JqaWe0iepa
Z+2bmjEqC/jZ7Ap1i5qQKI/B7Xo0Of5t6jTOYb0P2GyOA2nb8SyYmQVwfjUlJ7dF
TpeiZSkEKdxPIemVwsR4PCLp4Fk4HVm5w4HrAev4uR5O2gztW16TM6TeYH5invbR
YYl4LWrG5264gKBJBQ3TWkGzyDIOpDd82GmLnmy/UlvffHvTYb27uu3gvuI21xS7
Koic5cbWo3SH64y0P2lj+2FdPTM/ES63UqyF0wJJyvFXJJOXdJAQ/jIW+Eu6njku
OGwijLmv8ufAwjYtxYtlpcXzEk2h0LH/g8eU9sI6Ph+vcF7GufCZSuMV43nGUYJS
03DPL+A2mPZFbivAhkEyn/xYr/4F7VOmeUQgCO8Eb+btICK8nYJcWJHnk5WEQc4Q
BejaCWU8GttiXeHzMtl0OyWwte/8Xoe8J+VqD5iNHQK/TtBlMk/R6XveL3Lht/89
q+Cq/r8JJ2UU6LK5ntilbskgXX7UknUE0Vid09XaePpQ4hYBHqaKHaua5Uq5CSix
1ikJycRHnNPSYDMJWBOhkuMdWqj21872ANQS9zmY4QIQfNqTdL7st23yUfmOwKgb
Ah8nc8b57xc9lRQZIpn7sfaWiQsI8VMb6CBk6I40Ygpot9DLXNChRPpFuBf2zcfJ
CJFqpP0VVYFoAXcvcmyMv0WyK8xPaMr6g53SxuHGaTA7OalzgdAV+yYUsLqxxcRu
Cu+jruSst0AicnQ7IKHLDAPU5txb3SobHzqPLqLfiJZjtUM+B3dUn/7ihpra+CWf
zD2qjS9JjnBLzAEMp8/kqDwEF6CFGBkmlpj8mOcUzj/E+591DTtzJ+rx4PvN/P3a
7U8Q63+JcZtwDp0VRfJ9wqgjlepRU1se6fw7p02v5YPDcvSJRCrxM8hah/M9tLus
vcuNzpcumJtbXdo+8w+at4ZsCCrIw/57tdIo6L6c0flvHyTaUdJRpfAiXRusCss9
9G77RPmfJvYHD6aJRFeXoD2sV8UpPvxcxQHabKynxl7OTYQx9Xx4+eT5xwNJRGRd
m1scge//acUrI/8QED73llPPxmYkaP8kwYxsjGRsNJqsqDD5ll66H7Fjgm4orTt8
NuriUugyujYoS+z9z7+LfiNiX40UtzKKKZVbea7q8fTqzN/KPCV/FrlRNx2ZVPHu
8XC15TlBgVT2iIgmV06eVDEDR5BF7smERq/iWmeiRd5qywdRjCO3F8aeHRnuwzPh
UQvtLku9wPmuiE9yEBNqXVIa91WNdx3SvoJb0k0a6cQ+CH39LpjhvmcZ4hsLxDIy
rPmx9r8ma+fivwagztAUaIp8W3ee8pUo6iRPCUlvDMMlJNtorfxE7EVHYFPdHmWu
WzsVJp9GR/YlJx/A8Gn1oxKGJUvvP2cFc1qE2eRIA9nL9XkWtoyPYDblrGsAGBxI
6KQAtjy5oPUmYG1ccPHN+YocCPhMXJ0YiPeVrNNf98rLpDOCW5qZljPY9k62eyTv
PLEqC71vN3Iy1S1bEr2xvgb57MmN1ZpFwbjXE2IVtrzUu9j8zzgwNY1wugumM+/f
jt1JbtBDQykyf3uh5Q+Ms6EpvocH5opmgEp5u9PlxwG0Gcc0S8Zcb0DFXXBXoNnn
mC62dIn4di6l/olLCinPGWxK+9W53OzYT4H/xuOrJ9ZqcbCqsAx385xfj3mp2KqT
0kvi+j8U2h5kcWnbZkCcNoGpY9GCkfvxrLToxFuU9TLLsdvUF7xs+ewiXfEKhBM1
PPrIz/WbB/BIV3RqghBfzxui73s+msaXfHM2kZI+KeTwULYf3WYb/oOW7rymeMoM
PXK737bXbuAtW+L3omzZQ2KseY8EGFILMB5tVnfXhtPlHGMO61KEF4vI56oF1wc1
qNL3CKPkUElSi6T76yJzqKZ4tP8E2Lym0p0rjYThYb6iW/00UxCtz3ykx3h2hUbq
ql87QIUfiCQUxbtseGIHEjY+Lye8nhSdsedkMVPVEy8OWtcsWiB9YizQgk3zc+9l
Td19lTQQ6minfPJJ6M9PsNkGcFJsUKp9dz9A3x4F3+Jor95c0xs0occkKaUcDmc5
gxGY3rLXsr1jT7t90RhYZ6zvL0+FP9z7nGhTTl9VdRQa8AxmHfyh2q3tXwRNEaMs
brQcBG3yeO9ih5j5p+JaJBi63IdyiL+6hdQGC4dOkmUr8OMBnvlnSGxuqIdj/Tnh
UQ7LvU26FyWJJXSSC2q0/Bs9f3Z2DyaM7BgRM+jQpvTHNXWcUgA47NVpnyFeeggQ
fs7xSJy0b/p3n2KRwp4nGekcrx9j5Hk/fv7khTI1a07MjOP40l2XV/b+robwDg/v
eahZ7C+O6Yp3XIEUoFv4Uqaa57oCo8K52hJCirIUgLA4H/4cRGe6oohZbnK9hyyU
B8kPHo+6xwz4nLxFJ4nI5ivMEvTxJm8YgcQ0M0o+g1Mv1atAibpS/kBXAdifzfYX
HgKQOk/XT2NNA3yhD4Fyim/ZLX+t1/U4jbR0A30q+lfvU/gujIIh3yVDfCvG5+v7
UTq9hzFUEPiw0xLtXH8jpz9DNCk1pvKKcMRNTXPOYJZRYkNgkVbpigmdP0JWuqKv
FUzlP/wYTJdlSCaIsFEig1NTdxTxFAUIW37lbxx+BVWTwOaExKks+bWgELTGy20s
L+qHDS355AM50rU5XHPkl96eT9YQfekzBCpfzrPG454HhYtFVkXYiSK8eNCz1pEK
Sw/RGkbLmqqSIQ8s6b+AfcWSvbzMoAoHC0mzWeWGp2oSHEzIB2W01v+vxQWjP44X
lDJwdXtlmy3TIVLLrjj5x+FjEBWY6EVyodcCOQIpPc8nZ4mBIaKR+jH/GXcQFuJ9
KyE9SRnE+O9DYEl/TuH02pAMvygglxvbbGiXlidh5sc1WyFc5ADEq7yud4DSi/yF
Jldb+HwrxIBV52h2EuYvH4U10yYeBL/75bD0JOG6ez7qQ3IvxrP+h6j8iKs3bkC0
rS+xZ99M32MJ+1aR+De+7+oa4DxcMzD7oVN1mMubDI5L67VEj1CPnAXpZ8BDSu5h
cKnEZ7p5t09f2kQj8t7st+YsCOORXcPotOGFtHRYdxu/E3j59gElE5FFSkwx5Wgr
SW34HCDBKACC4yeLSSG+PC/8/G2UXJqffH5ciaYLhRu50zDIjBcJbtFLM59sB1lA
/1DbPuPzClQlKahpfoGHiQ0CGaFkX9h+xoWjjoyKeIuBXUU0C/Mx06Ba1rxbFXPI
VmFwSjf0/G96SKlkDGl5MmrhDLK9neJZCqGOrLWyFtpjkxkeZdUc6PaKYW3ELUbE
07Uuw5ehLMpVX/ZxFAuSHYldTdWtKa8umxQTG59P0ZX1M7nNdX1X4kXn0qhLPsLd
EvkpbbxHamvp1++qR3VEK5bpXl8CG88sbNWIl38hHu/jlLw3KPEkn1U0GJL7uOFL
Y1I6sa2hweLhjJ85SAsD9V3g2EQfKpFYMYdWfkNsc6cPzTyQgCnZJ47N+XIjaEFD
hWEQSegl4/R7qE+oLIg4JX5pXTns+M8x2el3F6j2gd3BgyK7eWbP334iXAMeeHxQ
gSxgCwCxXXs7ZBsSDaZ6zDalkOUWpPx4RAAi2BwnkGjQM22Fg9R2mWVyCvI9tR10
5CYm8cQDjl11y70frqCFJ/BOqv6RSimooq4U/NEXjIIf8Onor77D+HSQIV/J1aLy
i6wsyewe+R+ldcJ9eEcnsieJyyckqfYPM2emydRxmQBuMH7KHzvpQee61aWtSKBJ
aapUKjUp+zjIbPU9L2VgF6pmlAYXoxE0ABbKoUS9XLmO0YFq3MoXT3IOAcocOyJa
zvFlJYRR8NaPi9NLZdfKFxErh5mGGU438va8qcYfx1criNGVPVodPLBycv00+8vM
b5IiiIOazUKzqJiLmvOHAdSKxKrIVIYvQO/z3zbnd3rYzjDqcDmseNRhvxHopCyp
tM+5/L2ZUD2/E9csJg1NCrTrZ9sRTRbTqWvpM4ARsvfEQ3g/FDmse+LyNNW/NOrY
j8NDqEQAJ5AhB83oCL9XdskQdKMcVnoQluL6xtrXO9+TlzFtDUTKNP0+XkGzdqg4
bNA31+nNvwzHx3MnsTzVay5rezxeCBl4zi0f0B5t+V47G/3W8Vt+6ZbHQUU8IDkC
/p7FWx1QNxvU5qu6ceAnNiRRk2y/o1RCqkncoLjuSURZfQCqsxjk5WvxQ3vrHmsW
Oq3ZZSRa+f+UYS2omiTkRDt/uo8IoPPZjRPFxKhl9EgbsZUEa+i2nzvSw3XrchaM
LJEIjUEzFheLdIWdUsjHGGvJQuF0j1LekndzBJc8Nx0VlEG69NU6PLxDtnpptMD/
q5o989RdiWXZtsZka/vG2KZjxAS/9uMub6RYzs6pDrCLwe6QcUIk3RHCX2ZcBLVS
yMFNK40I/AaqQ6FkPnel5VqF4g8xNHdU7Q1KVMsvovU+dCGo618IxJa85uzlgY6D
2EoxaAId0dpgbjl5OoPh3Ww9Y4jpHvDeKqCUmW6N0tlNM37DGRt/7BqBlvXkH/lB
ZTPc9yPFHS57UdXSlBztcZt+0o4RY8bzW6BoZjxuFA+GVFDoMc+d0cmZMMMH++C8
MIWIWGnfjZF6plLg2dJtWK5asML0Del6K8NGh562bZto20dYn8Lohvt/IhFvtL3I
TxzHIXiOF//wcHeN/rR0xJ7btetDLEulGdH5GS2XmDhf0i7Oi26iKSxwudhMIZjb
tgb20de5TBJGI0h7VhrUFAiBNUldhsD0XPOdcp4XaBMov65hebrKhAfK2n4awewr
l0Rt408Rw6avQsdhqm96TJ9QMOIOLkxF5GYKuIe0KKyP/ZDWJKLuBCnAl+paCjbs
bAXPimJVBJxHE1g5/PZCIp7YGcn/gAZNfRg0p5ld4jGXFZqt3IbEoueq2iLrYpOZ
/NIRirQdk8lpwICIufBoIioyz4BfXgadXYFalSW6VsoOmxiz0/DE9GB0TnsnoGM+
6XeYYGFXysTCP/f6guqzM/lSaN/e7nr8e6RxwPSO+11P3Stxk+whfqkfFjBYb1P7
AkKjT930VyjJKd1w0GaOt3JAJqKXye6Htc926hFphrdf20umenHtpuIxGGRJcu/n
UvLCLpHnv8dbQ3C0eszr2wVK96YJAAedHfF3XxU3WrfPJBpXpGDTONxBPVsAwQyT
X6r9fflFl6nyQEwmw3ogXjpI6D8Y3Ipei7AWtP69MyDx+EVpNhOmdNRg4sEoqn88
v7sJWBJOjO/CQxUtte5kotLOp84GK4YP3g36m6wCFmC8HpTdG++g4T4HeoonqTYN
TAwrHlBt8T1xyQt7CKamxbMlewj+rlFlSpkX8DlNa2ZA73M9I1BJqPrPR8WvBTe+
4erY0TN5nD5hBkj6+ZYGUzk/gOV/2AWo/fhgIyAEthSky22Y0JrrDCXRLYCx93OF
f/3RD/Bpak+NfIpqDrnxbzx65su5JRmt9as7xg0fWz+G8UPo2/CldnTsdeMRa9/a
VXGdLl1mDrAsNLfcijrgi8fNr0tJsF8OIomqAHqR6eZsOgFT3JFMLiwwMRwH0QN8
5eV3zyZ54/dfKKINy4Uk34nhsIVk73bfNEsZ5NAbAkw8e7pfojBlPcw5PtayJHhk
rCBOIP8k56SmPsjpClXZoMVpcP7CS8g2eXp6RC5tgromyHcTXyI/2vbt73gCu9fE
PfYOyMyt1D9ETx8hOzmcaJfbFWn3LhgkAxGwEVMKXgZ1h7/bHB6TalssVwkdPujw
j2LKA95EUVuQEImEzP0/XahKXUwNOu/gFcSDaRwsDWoO99zZQwbzcnXoa36OqhKk
S3JiyUrsCX1Gy/8vqrNLqUeDOXxu8vzwdv9mhGs4kqg9FCIM4iCT7kD+2w5Gs/Sq
pTG7p8AqlkR4g2hlo0Pv1bfbpNjxDcq+LrTiOUkFPh+IQp2K1suzmL2rP5M2St5G
d5S6hG5uA8NEXfmJA4qItk2hWpsS5A/fxTIUB7llGhXFVmYRsLJQxQLiXt5KdZDi
igZkWH46YbO8FUF0HOfDgzVxtC7a5E7Wn0toT0toiyGvvkfARk444pX6z+YgUj+f
pnp6RoxnKfNxj81fsPz999H0NVGPfvSYSa4uUR3V1/kCghpmJzb+DBymEX1yE71g
PPsdHxXYwKthWgTFgtLAv+1W/NuveGWIJnpk83LX9uOMuGwTCVlliDDupbs7OdKA
Nuu+ko5d3xB2DfEBczshbUf1JFsWmtDB0fE0tdZlgHWPWaw8SNJj2+qpu1AtlLOK
M5Nve5PPd2IDH2SDI51N3/P9pdKdF/zugHovNLBD3IXYF9HZnQLZsdpdbj1LYDyL
c3WzOqxhw8xY3ZANpsVnOmTBofo24itUJogNE/45qLdtK4sog02Qbh/8fGSThFOQ
j6AyDFcfKdHcza7zd0eQRVLyY6sLEzUQDvlZvHjnIC+BtCuD+1vrr79B9LwmoET1
few8rqGzx+Ym9y7NbvYhEvCd3UgUlbEaGOfoBaDg7GAaYNri0IuCeUpaV2agKcfH
RdwZ7evaCXaji5JGXJK43/Kjf+AXdIFA+TvIMTiWpC4GlMl++xMdsMJARpMeFVlF
Mfk0TNYiKCDAYqvsUTjKJnmOT9Rm6brVUI/0/jQZ2DBMyIrdoN54Rf+UCPgN5GWh
OeAc5IjjdGoMVw9P7JyuswbdeG5UwFRU2WLFV1dhFIsaw/w+x/SB8U2/UCAh0s/C
ALlIE80IxpmcIlFkrM3Lp/S6n1Ffbt/IPp/CnKbKKSzMs+ioewDBAZFWunyMS1O4
4rOGj9nAdPNuQbVLe9wbfog35KhDXmhTXAWF0BxR2OIFW0FIlIdtuZEDhl+fVqed
Q9SJXrCp7mx7gBWqKqtwJ/Ny+LKWPjm2jS+FV+5PmQStfV6schlHgtrz/T8RsG9V
xstzmRExNal3QMVr9B2hYUuepXIeHK9NA/BvC591PmmcKe4Fwi8UN6lpJnr3Vuz5
im5M7AqdNZzwt8xCv/KvntzWRvxogRntGAqhBDFXiTIyNNG09pXrbk/pHDt0IIdc
mKXLJ7j3NXEK9bu+8YjUdaGVTCXhAmgaotNI9kMKXV/AMWXkqIG0ELMmblBBpbu1
7bKimMYi9IR0c5VgXVa6jX5eOvAW82mQ/h7foffHUfm6IvRulG4OkNXxaRF8f2F6
vTqcDdbWsv4uW4tfMJaFnG/Sn9ENbsAf+z3Nrj7u/dWDyWUoanhPRQWslmzX6Xk9
bcKQOcM/7JFq1cga0DUsBR8kBHzsKZwETCeYnndUUrQ+yIwgbIaydHX2KMPOIxcR
2zJboY2kWhQyDm9e9l4v2Vg3rzo93c+LdNsy5FTXb4uUYIAvXto1DjeDQj7vXWZe
3rID9IIlkW8X+1q8Xn1cHx9DTgSl2SnphSE+nYxkGM9FeyMwbJATcICXbMu1l1Pu
x4CAawnth3+zkVNsBOK+lwYFWrm6ZwDWEyZSpbjoH07mhFRet4/sA9DCNHc3UvzM
0NnjuqroREGKrpzJKClxcN+dNbgXUHDmcRB3pGhVJZ6gvN37fUj4vkdqn7kNTvKX
wnJbfm5K+CoeciXF/mRFdcdmI8AlLCVKD4aHsTtdKhx56ulGFgxvgh10vo0TcLsW
iW4S48eBVuNbNM2zWlK1LSApP4C1EQNfmV9oEk8RmvWdNfEC2dKlZYjVuXemcEZZ
79q3tAxqk3rU7akKuUmPFFJ6x9cQQ8FgVSxseQ3fY86sKG3kWfFfXSkOM5QjlP8q
7mx94x61MYWvZG2ZM2qtxdiMqlVQ0dUQz47urshoyFJwMeSRc1cT28gXgINvl0ql
Jccy7uepWJUkh56arc53ScIHJ5eemkuE2A2uNl58bIS3roypAATHwGeVaGv+X7VT
+cabCB9mO5O3Y3SRX0WkiHbQlqishM1l6Zgs47jASkSpZdvrkjhIif+C6G5huC9t
RmQgPbaL/9g5CZs4OuZtGnIFuZEV0sRc9MVh/5GTyX9oiMW13DJCeRfPljCO4BsS
X8kCklGyOQp7+XB+ZraC89K1I4oQcqUw7FiTeNGqKbhcTO/GCJ0GIUDTvrfMiv2r
PCCNsMD1gn5gqC6HVlWvDu/EQ5spAtvlNX/9o1YiPEbBuya2ZKVDcYgX+KeLP8Ah
o3sz37ySorJU1rKHYfSGItuwUMUK/ZqoQASisBOvxyehzA8OeDf0FayXTog+CXhP
dqWZlPItbj7u1oRI2UYbmJ5S1d4dahZ81mYbNwHnQNOrIg9QSvuXDlOK6G6k4dby
PZ7dSZILy+HPBZWLn+IbE8RloVmhrrfXkBXrx8YC0hJbDvMYiJpxi0yIafUuFxww
t7FH/BfGZOWTitevgcVTOjRKfxBm0ZqzNvtMtHfueXdrQtFfxG6qByyXOLTlVRvh
EfTlMtdGrgmu3ve47HNrZOoMzPHHqrJOuQ3TR+905HZcfvhmbGTJD53LIUUzv3bA
/oLL/bi1Ou6oQ8+YajI6WqTWVIVzTO/v0ygsd/plCDHzk7NwCU041/oQ3tuGb9Ab
CLSJRIOmBvdabntkm7LGqj/fN/rF8aDiaKT+rIzszD+f7PesnuuHRoC2yj1zDdGt
cvEiwp4MHM+bDlDQzKsB8nkhQdZzLM91AJDcYBPREf0ex2/fdP6G9h2stKOuc4tK
HFx6vn0IKvOKBc3pz+ZaA7nDD/wGa/y4Z4cLIt06pa/7AHjOR+CjPqxJlCy+BA6h
NwcYCiM6z9Xej/Am9Qv1dx5LgMZrS21cspbOfNAbbaz/kzgBfM5Eoc/WMdWi3ftW
ZVugACmDNDhQOPjH1JJZOn/9WeYbU0ReLqIpSOT8uhjgzqDepwI1AeBat/rLgW/g
J7YueKxREOKHCspHcuulJrDvCAPc6BwVQWTKjtjjkrPtJ+azfmkQ7XWcC/JIX8Dh
SQPwpp342+XAGdHP4sAyBANgnfGEhhz0R8VYXluO4XjjY+zLt6JrdNtrhHzdHn1N
gOZdEdFFBJnbqy6DAuZTfGGTaEXSGaQ1h4xF5NGxpgwze+SYUEaYg9yfV7NuG3v1
gy9j5Bzj0f5voJ1RnNLHLmGrFhgJJ4p5IznmnZ2OwRt1tjv6yTD/Im5e3nKvAgEf
W0UN5BQb0UsNOp6wmhs0ufgCFs42rN38RoIrTD1MlZT9tcQa+SnQ5vBXUBwuZbW6
N8BVkaijlr7XyPRmG3aASckmNZ4wMabFTvW900Kxkm2lQlzLc52VnfSy5lkcNjrZ
qwQGssA5e7yAQEesILBGC41FC5gQutqDfWgZmTgAfL82tcTsPmaEkkiMo/nG5dFD
vm1dOCB4voeiFlR6CJBOEnhl5JB6/CXGRv9Bh07Mi5B7UCQIjpipgGM6JLYmVfg/
1URAM3YU9bKlXCaS7gzl4PDa6rxl9LsFJmp66sPzvRC6tvrrWTHfXH2OyKohy1cP
U/RXhqymacfVDD9uyd/IwEYkV9jw3Ik5SJZLJiovdxDDAdqgaWih4Z640Ldnx725
VAS7PP6ARLH/Sjd2ZUAIg6j4QwG+JAG79Pua7opn4fzojEbEJpfKJ7PsRfC8RHB8
1QJuK6d8lWLC8OjJyCgjf8o2X2HS9vZ8M7LxgEii5Lj4oIvJjkSWiBu/CbN1xe8A
ctIiqHU1kVQTszsDcxa9m5rCef5rIvVYi/cTDlKuDE1ahL6BBCW+L7xl/nBilf8o
W9EQqsrbyjYy6A9+1HWRAikx7+7aoF1gIgrMxoMAOE0CIwj0Jebt+ftzIXBF0I4z
aI4J0Cp/3eWg8ZwotIx96+6dvgqSkmaT4NtktefVb1ym8L3X7nhRl81TEZrSOBNt
geQEUBh6u+dsKVhjlfEmQjYA+vPGyrBrAkuDk8m3XeqcCcHhxHCluG6jnBpi+rkT
WSvZ6gJ3FRH6MytlSIEqNKk4ftLbbe69BrO6xukV1Np3TOKGHdmKG+vv/nbeRiJs
M2+ivmMDgaldMlM7JvCQ9BQARclCC9R3OK5winghOGFgU5L8yeHWg0RtZhCf+6dT
0go5Zt1pichedaesnEiZlGoLpEsuY5CUrIBLth/N6HygX+clneucDRyKhd7h+vG0
TVqjL15v9Thcz5/J+hSBWPthmF9PgxHTBAoB/+5pryF+Z8b3KWRZU60IqKeEYJJv
v+VsabLbotZBSk2GHHjkarkFK8oWEbixfENy8M2i6cUCLD3uizN/ysBLzn5KTEPj
OYqzP5TL2YNwTWM4s6sZVRK7piQ3K1KNy/FiCxhXxuKKy/ZEgKIk/4WxOvMBXhA4
KQYsJp0/El8hdOYe5PLIb90hfV1+q0nJv7cAYfCHWQR/j+8oCdNFMrUOwR+G3pyD
ooFOe8s+sroES4uqfNqLDgE3yBbH2Fkc5sy7kBjze2f/10sChRRF9d/VMPjIUx0F
C6oJ/+iyrgHubu4clYs3NgAW7m45ZZWvsy9Ww9k6xDH9Sd8N3WwaOyhM8mMUwFwn
nmPzFRcAxA3YJi59NBJ5vH8zCoJBt982VnWUEdUQqcx5LWwsXMwjX1Cw94VkZSqz
Emy8f6AGvH5oJb5uA0DQJpRghF+PUsUC6LfjUcC+YFdPv0y9BXWRLJhu3uDs8vsn
4yvd+vsOARjJ55AbQtNSx/leO9UOtJ8iuJduINCy+2tjQT+YnmaNwpwX9u/QQjdq
kP5sONElYv6ALVZx56XtZCF90cbRmeGJnuy3vgwzJ3dP1mrqPRbyphbpdQ1giDpt
bw2fI2gdTLc8ED/6ufaq4aJeKjO47wT0ui1HjwNHqHG7YbvFFhv+xEpjtMW2GTed
VGCmMKmNTUmaCPvcjSKeQTcfZjS+mk8aU9f0A8X/N2ZgvHjMc7XYRh0LZomu0oCK
6/30ViUpC3veAcUMDuEw5cx861giEhqD18HLkVOwr79D6LLZXeqzcJnBIXSqwd/e
D+O6SSvv3jyJGMIP2FYP+7PWMTtbnQhymxWCNPU9umZ3fywQrgr+jKGdRkemNB8f
CMvGZ3O1FSWHluFyrKWod9u5+Yy2n8Y0D7LgcnYhIkUz68nZztpTJn0BnLiSA5gM
jMLrwi99QF8pxtvOuGDh3WkITD+eqtUgugRWiojK8V4HsvPl0j61JvZApw03ZpoR
qu+LznIan+2J6sq/xmzbt0KjWVQScoDBEDF3VjOUk8vdB9JdtnayqujzRn1PzFqC
Wv/2gMCoZViUxid+sxyyxThj5HNEiIpOWooRzu49IQp4nmGbbvIFRdd7t80NHb0V
umA2WMMYaKXht1H5T7zREVQedUiFkTZ7hvKq4Jio4BXUJNm2cWHU/grMnzqHq1rl
3VjV+8ZfMKVCUJuEmjUDthfnxwt40GDbZtYBdZzh85jqzNDnxQSU81UsSUKFcebT
6sBfHVFyHgebNhFgGYIzObQb04vGu8RyaWcjo6DJVmLBplG/FHCboXVc262vyOri
6K/2+SlPHfm6agZ0JayUe84diFBHiTbC2HSS6Nl9mtdH4WvFGO0+3meuqA63ConC
i8lJ9JbZ8m4n0BQ4iL/DLNecG3Y5vS3TTDCd68mBMV1Ui/u5LMIdaOZxNun1QGrf
45nvwtaTvuANqq5LCSMfOnnX3Z6H7LH9Hkrz65pHeJ8HKCIVupJ6Wdj3DFIy5ixb
szvBQRXbzNkNW6dK775emOQmhq+dONoNzQBGJw5ILf500MZK8/QwnKC5+953txuv
/KIDZZYRfS4Bx6uTC/nWYyjOY6zBoSb7VX+5ieeexyMDcBLowx85C3gE7wB131s9
T3LEz29K4pOx0vdakzwHThqdAkBmQzCUqOrOyqU8FD5xRRbx/H8nMRYHpgZkEBhe
AVFGxoBV6TkLoqYLsLhejZWREIXDEGUIu84oq0CNuuEY95PYh5DrFlFHVaumK6mo
ACnSdKxnN+4UofcEII2P8lSJYd3wceDhXv5PDMVRhMZn95813KF5E6urrwK2DOdr
VeElC6WnMfyQFN5zXK9dy3LP7r64/bvSRmfvkgTCsv43dOcwm//QuFU/9YXYJgGF
427t/vmOFW3hD7oQuTgtWaMNanN00HgTTlkuFbzbcsEdNANm3X0j8OVFt9pZeDbu
etnDhB0reHBvz2RQoxl5hZlTNoQBzeOdX2wbdSLpKjx2/vMOSEmC4J+8NfL1BOdb
+5MACqR7LRKuF2rn89Fk2bN6efTgUudDtjWp1LtKK++gAfD8/Sxs/BkyH6q1cXPb
EOxWLO7K1KHC4PKY6r2oRAEGq5bhkMfIchctjz6iQbdlZgh0a8u+h82Qfd7/NM31
9jZfId64Cy7gtD2tZMJEWi/N0JV+bGLjzfYA49DITelzvO8mMX1Vh8qtIWUiGb4i
Og8os2u9/xdjrAklR0JzAbGWqqmS7kZxv/QzI0w52HoS6AY8FIoVJNAn6aBT7DNV
bRniz56sufjS8nH8Lei0Ure+wAlJ1Te3FRubUjBd8chCGn2kMQgE/pzQZheTB4xZ
jQmsWxzUfH+TkjHGTTFj5xioBGeYW0qgWCfKqwBH5inUHYY+DjXt86xWcgvWWys7
RZpQp8A1VVEsHSClFH9QDkW1ftU8qJLhZRJPKf2B1BwJRYGgsoNhjg3YO4X1Icrp
q63Z/lRgCW7+fmAza9xRFzT1/rHIurWfEe5JVx4PE+r1vhxiX/hNYArp+VQ+7Ptn
6PgSBGg6rQ+1dpWYFpa9AwHXa9USkk+8ZHugCGX6K9dhZ5SWSKWVBqIhtxpxeTxW
R2N9Qkw1XHix+DPfIjmrZbQBY/veoLaVeTB6a53Gp0YHaf0ZpizIiazvfkc14jHO
InlBNiNVr3S9ZbKOsl7NObNo9r7VExo0xgUXEFclzBaS+bymPPkDhAVg8nFhBANp
DT68HN2mClmOq9zd5PGIFDJGuXrBFeVPQdKLZ3XJAzrH30JmdAbxV0hYar6i7O+I
X9kaoS3+yknR4DIebUVpfOa79VLGOlbSGaG1q7j25sAqXKio4YQTYgyStda7wvuP
ujkj0DRdQMmg7/4jiJZrC6x1L39s4KsxlKEU33nKgsCOcj/ft8m9H16SBH7YYlTv
1iYHF8RwjkKr867IAYGIMmYOlcgkmhCNC8Y6KKC/g42aSNe701TGyOfB6O6+j38X
4aLgZ326B+DJRrgWb2931lLcawLUkU4miDY3uYzUJmE8Fz5Gu4Zu+BXH2ycK3KXG
MRSWvL0rfRBo5nt59Y+vcoA5Bt44b4EIBO9yyg1vEYwPIjlDLGAyF8Q77dEYC6Lo
vZ3C2qI6T0daWa+q+rRQGkumsmNBnKHQhRwyy/n7Zjz/uGJy5KAfn8hMngVgrtaJ
QELuMjRa95bw/zTZDpqsy3TTQiSVTYM5bXhqlfnXwwFla9bnyWTntKPWmEEObB5H
3ZymLQ8OhKcw9jJ5xqHkLJPZr36SAF42WPaCtAY2IQZEu+SchHMStc+aVTxQRy2y
iDyZSA5t5z0BTcz9l8FwJAHCPlVG+JcDavTjbEDR/IYWLHnWvHVhwLCrcf9hgFvf
l/oC50PiXZTh1Lc9/etg8KN9kSckIjB+bSChzTWDQyb5qytGjZ9jizrRNWap1POl
w2gW00zYMMeBtSh8t5QWWds2owgmEZnfDKhx7f9hzd4D83VDxUW/oVy4N0e2G59N
u4C0bCnFa2d5sil6kLTTz5BQkJhjxTmRrkYtFElqkpqxbq/pWWX7hyS5dejTET0V
7426+PFJXUiKVvWbUAbv5dAB29uupJuQr3ez2Et5eQ0HRvsnwAwltBU3JvaHiV3P
i5v3tpHlLRXclkHQu3CU4m16YFp3frbKNcH9Qaz62dqWYgskPjOb9E/b1rcqDJPl
wTeOnTnZRmL735ToOPJcRkq18ppDZ1UZenm4C1QegLHuu06Rjwl20lf4PYcWITB+
xCiB3S5gjHVKjF00GnFh+OjOEOjOfe9kIZIPZ7sHh5uhu2KCgkNmkw0L8Ut2xNb/
v22GLW1hx9e96O0OrgmmK+ivM7s3hj2aOwtC3URgcYKnM3Ytw9Iak1bmKXO9xqSP
X59iZbKoL1fgQW7FMp0+0H2r852fBNh2v8NfIZ8zvQDrOmlXUIwhIRXIVFeuqwS/
BFZ0+tUlEdfntuTcru8zrnGy6c9N7Om0erqjb4az8PdAT4hRJ77wFOf5PA3A3tkI
+VylgzyQmLZhzb/Q23fffO0+puqcMVKT0f/6s1SsOmbAcNSvpXc0RXNKLWokbLqF
UD75vCT/0PpIJQuysH7BjeBLHZHVLSPfTmEOm6lJp+nCZjkAqgwX8X3GcGlaPjRZ
Dr3UEUW8RU+sKaXsBkLa7UfYqny8o2zMaf5zA7lpin10idZeREbW9uwFCOC6mu4h
VUWA0A+6vS9GO2vVtjRWTGfey2F0GuQ4EiYbrx8+Iv/jCbO+ZJT2rNeTacYhsz5w
LqtS9pTA5LO1d3OhGRyyM74QWgS3May6K1/Z8a5OkxNlwCZbGaH4auDAGduwOrlr
vv8wuQHix1SMo3RXKPK7R7rvjaafUejAz0aQ/FDhI+CbXP7VUSNn8j+gojZ/BVwT
C8Q1rg1JFiwhFoSdQmk4xfjRXLn6szAoa6fxcNwy8xrI4PYlLmOnp/+h9NsPyyXc
WYQbdRZtQM1XEONrTT77qizXNU6c4nBzuytf0VUBE/K4B3IFxiqTwd+KlT6I9H7y
QuDw5P69nZVqpjFhMt2ZNOXmOVwMftv53I5vp8rYCT9RO2zV7+g3NQFMJZjYFdeo
2r8qAkd+ZpoHWU64FCQ+bY/m9sURKdx3hCwQL+6DJgIewLvXUjui9iEltP0A1j7d
5UvdX51ntdywZqJZ5YV1bm39ufOLjMt1Jz12PGZQfe5GBmESZilH5Oy7YcoGfnHO
GdlkJYRFr88HmybgPjGATL7c+J8GWGwlivfYRVEDgf4QgK95Za33Awqn2TwiVtp9
gkFq5gUE46DeRdsQ9vOutew8dou3Gt9GUmAfvESJxn2//+Sn/HIwM92HcuwblgrZ
p6uiVCWWMxS4rGeCrku+XfOJ2FpXKrf3LwU6qJPpX/BAe7SdhT9SbXgItEExmIe1
wjjDiilwXyjVPk/TN9zMsgn1irNQjnwxa4wfToGg5wTKrrcUOaDjXBmP5Zyyo8ba
qfo+o3whQdJH8xvAYpI5b0riCaMKI0MD4R8y6huWOE/9a00V/W6IEWoQskiao7uD
wr9o2RGlEyW5bgjSzHxD7XivGvoVR2QWxcNVxNjRCgqujE+uU6qFOdNyeCzztw1Q
E/W2Ha0kGfD3EMEhXduBudzXqf0LX7tMcJ/CcgdOH8y81Kud3OQXIf92bjut2fOT
mq1RtvQ+Ar2rzVGIuRnj9kb6YJu2x8RA+vICAnm24vOxri5kwm8zvYskOig8PS+2
HRGpdQi1ofLe5vmir6w1XOGs7O2/puQzMf4Cgm6gwBatZwQY5aDyXCIhVnDFL6ab
r7aw6JcT1yhcMcZY5Grb//+mJe49/Eh6j6vMUH0DxavJAuClBFqROe3Sg7UimjwU
qFBP4aZ6OcakI74l0hAQ2Zjxa1mEy9/z4XD3VJeAfN953kbO+FI3gXmgO2s/czC7
wWbYJ+srauFxYMejHthAHNKo/17qg58rqNGEtcWtesdBtc6QnR4qEm1uCzEmAR9j
BVrZKFemzYD2NEjjrSFZIs3q4qVNxToOYAk1vC5t+z0znoGh3KLqPfOweyAb76+b
Ihclzyq5ZlZNBBpJTB/uYAOPBzFNmLt9Sd+DChhLbGDpWW5phAgUHXvCtmAq9Tu6
/dq198Vfr1b4WJd4K0WoOQYYLLQj4r2wutL0Ts08aVV1ZAVNBxYV5vEbu7OdKKZH
R4KdsRi14i3ylOQUm2Lywm18jOBR1q/gPf2WAdPEdlCRox0E6cB2DI2ahVBE29KD
TrRxACCBQgmooZdniDJHr4Im0IaOP/u3XDCBiHwksPMDeu981xT/ZBp/55if3cb7
Q0MQPFnDR9WvBO6Vg/FcczEShlAsF+T+HdkOl/AkZKYsro+sm0SkV8z0WhhFaJ1O
pHay4qNqwF6CfNRSR4nMvhwW/e/KIvq2JzFOrGm9c6itz3mUjUZfTJ+aCItlf8Us
Kn8FReibjxd8AGRE246gWI79cnNrnhKXaw87Iwi1Xv0f9t76cBRBPxBF7EckNTTc
HLL/vR8iV/TNBrjSVrR2Hl7BhJDBT32dH8NTck6qOG82y0dnvisjKAyxyY3u61lR
39HbeaASu7J3n+DAHHvEiWStwlwuD19Kr/h/7Vi64cE4bnWKHJW2fX3y0/rbd9v/
6E1f4Z2/3h+hcuHQzhq2ekhdBCDdfabm7vtHAhqkkzmAHrTFHZcUMMY9f79lnORz
l4nVxs4Q5pPRyJlXnXshvkD8lbEpZjJrntcc4gb1YDR1jQaKNhZOTJjKNqUGyiF1
hbQYgD1VjtOSazPjCmOr0d0kJyMBSxSfOpQwMAbyWhR/WOigea0wqB8nkcLIzLMU
mipt52MtfJ6nedpO2eUxXEqrybmKvTUAGMuljibknY054QJCEMNmnLzX71s1tL5q
KTrKGckBXU+CTjaQGyzK2FJf7PE7ETxz9uZryvS9BlIrmazAmp05y9fgjx9OnFSt
cA56RA8ocfMpmWaBkTKAjlaJNQfbNIhK7+4abPYdt3TdEIloYTVYahqmLaY59ozQ
TPzbt46PLtBlS5+Njl/eKAO0Gn8tor/Zn/BBY2ZZh7hMFdaCKSjgMkg/tID/15Dv
ZatQJnpVvwKx1NNcnkmo9W559E9sS6hSKAPugSoZi4KzNcT3LW9MKC2kNJR9uESB
7u6amtD+0zw+9gInYo4XOYBT8TeHLOnucboC6BrVn1YWeEV0z7gYOErh8AupVVrE
/XV91q0XwDYLAzTYZua+4PU2/UuOwyWkCCX1TJFtElk9ysFCv3u7tD2Ctk9xR+oY
KGsAk3DePeqw7Q0Jq0Kdv+5GNP9T2EMHhxBUzOtwv6zWJ4nu9YfuAfxWs+kDwqgV
ZBP3b4PGurleWIKht5N1ivAWccdyWGoC2DUZsTv4hzM2aPy/C+TXQwYg4ch3Ju9y
y2tZiBEldrBuzZBf5pY9KJ+QQ31gtkhNJohS+L/CbNHg+Rf7suDhHuDqrGc82VmZ
Gj58Wpz+gFd6ypz+j7eXQdyhRIwumUrZSR3ATX2Pmqj9uU0n+KRz7/hqd0SHgrFk
atjThUbBq2ZziXMPRbLBeGPod1DeeC/A4wbHPLHXGcH2GOsO2MRKyCiHs7Z/4dbF
jze1+J5xzs9AR1QM94JE717tWxBoWcDescryk7nOpUKRyxnxkkmQzJ0SpZxG3440
0K+8+AGs3g3Dj1ZxzSIaVBjOlLD1JaiYKgFe4VbZe1hYRgm42lhTtRJMlRSI8QJZ
5FkXcuQvE0H4veJ7k0jJXIl3kYqqB4RbNKhiMqVWnGk/k4SKr9FyOFTmloABDktT
7Tvb2HuuLzR0XsREdhyfrDAtTuc7Ox5hX7mJsMEySxFAYU7/03S3DhnFRGpshz7L
yjCwv969HynN9XnWzk5U5b+iP4fCOyrMNbh6cm2u3af6EP3OKxcLtcGo/egoRxbA
YzshXqXuewKpZxoXtLGu8wVrHe4UaTo3Ge1MRJH0yKCX8TbgZBeze+gcpVNhCxel
wEu8F4U0rFKYbsrpLEMcKcxA6AnnwUuWiZsleEoApoquskw5EZuOnhBUES1ddvoq
6NVSH0B3ZRdEktXNS8VUDSMCnVN0j6Ml/oZpEW7xLTT2yqIlaXC79PT3eaDIO9Wi
Wsm63WuA/LJfbH1gAiLnS822TG/cq61votwlKgEkVXcGJUhJdJ1rWObq6FiMk2iZ
E1R6IggV4WBrhQ/GJz+xsk27xg6mNYRl1vwMOkoVxdVOk7cC4vJrKbAMMyYtiwrs
13Tt7DaK1c8vLdZLrru6Sc4AwCgW+PLE+9D7WVlHBOaaRCrsREUsUOQ4PlvLnGmd
nD4Xwg6nvbKGqhIuuxIRUSg5v1VsAFGDSLVZ6BEVtKM6mWUSoV1UFsF8j2oF7HXK
nwsQhEml+j1IulMsMso8Rm6aF1a5ySbM/4vI+JPlbcgL3aejrpoufE4pMFObySBO
U2CGB1Dm5QRkXNwQKkTO3qZDDyAtmpmX4/nTyTKXy42478VgpEFAK3EqosOSu6LW
ewxGBrUwxF0Qhc5DHyh16N0EhIHY87jujsYuWqdwOBp2+Xqm/9x/ua6hFgEXsoQ6
TVPRYbhl5ZPuSUVMahWCduw+TvvKaTMz75DYLCbFh3uX04pWfAZBfoh8PmjOSiEb
941pJ236W3IxABZxu5gA79yNDrPv6G3C5H2q8rIbaOBQbEz9hPSjwPpSCTLVzqeL
9vqzveOCiJdcroH2GYxhOAUcUCTp02czcvaFvyc/c0D0CnK09W2YxD5tjDBXz0kQ
xUk4Y8QYLhuQwwK9vuHWsgKqg9Blr+PSIoV/gWiSlszfCL/sUBLpAjk9vDPU1r0f
eqshHBpfzVeVDlFRd5QyflrMWfDEauEAJTxRMyMSKtMGinm3xz4TIx6w2S6amyv1
pSqQpgD2RPVYoo4VLYarKzM7ug9KGjzwJ1VhSt6IVWRNuEwABuMP9oG9ImECRzTQ
Y4okm+XUDPz1VWPdEBmPU9nJaOl22SnQaXAFl50+o+paKsoc6P6HLztp20Tfrtp9
FMlwnfUOZCxS7ZfKPsOAQYCfnoCrID/OT0onEuGrnE/lGjmnRUK4T/DNjYyhTSKl
PaZ0ojpG/H12///09bYxO7Lo9E+C+PnM524K0vUR9IAhDA9UZCP5IE0FG8AQyW3J
AtplHMseXxMVTQV2m5RSl+NF3gSClMPvYu+EYWU5ufb0H0h0inN4GeZ7HuIxJneO
2aq9cb7uTjw0oktBh2rAixR0Mdrk4oj0cZicS0ofln4P34mk/OrPjQC+al4K6BiQ
lOO8xzSAC+3xsabMgfn7JPQI0AGEgAI7opoIregIDVInupk1nsGpbmjQ3eFeKaGx
z2ghpks/8dj09jWqxLMyYKA6vis5jtUfj8uva0d7pzaRHyA9fXDOeXZ66fd0MHF+
+U5pPgQz6Qn4hTRZylNSfdUm9xseN1Q+lgds9k6PMT9qtXbLFI4fmI/JwFnN58Qt
Q8cHepPrN/cPyBW2SZBQJl3aPP5E8arrOXCmIY0XS9/MlX/R3Nl43aezrhbrPVMy
Zz/Ro4oXHnGYldRj7pWchK1NxOS0nOMIDw0ECe2mk8CO/vNf5J7urnIOngYPC1Q9
10FSxZtop+OiO2xwJ4/NA+oIFA2s+kgx7HVgbbqRgVyE1I823I7HDr3h88o2Pnyj
kxNrqudiHyUwSyOuysqgTyK2CnoopVW7ZylFPSC7/UzcBLe9nfGOizin8JrvPN1J
tvbMVL3rhouS1vwA1h/xHzRY79UcRVWrCpB1AxsYAAAL/AOAOolmVrm7iZZuW5cv
CR9FszTZTcFYpy360lXb0NOVieBhn3DKWQyC4RVNa+weyXS78HkP+9phD6pfYFTH
V0ESCETFwSbDCKtR49j+OyjLzEvu7YW6MHxqo8L2R6rEJuzogWcGesU4tlN/pAAn
9E0rtebNeh/rE0yJ7DAjdUEsUmINKfcuNDurSXYzarixn1twYrgxjr1zoRKtMal8
eRXZrdoXz9U9F/1yczottguQlRBKGIZPxqKUmhWRMFJvnXY5RqDPUhIcHlt1C6OI
W37YBuD9G0mBgZ/6ySU4uvnXPzSqDWBdIyPvLetXcJIvtTwiagEGY1zBZH/XU1V7
H/V7w9TVY+Gu3yLVZUpgPz9+liyiDrZBfgg1cGS9MC+FFRg0Pb8v7+QYHbnCR7dr
QWWr0LMMyYAIdWOAmPf6Q7g8jaxupEqR2kE8PqghUQesNY5yuI5ejMhRjs/0xNdM
r7KPTRlEa4WpNBycnF4cW/j83vLRcDYPE1dnU+opI9FNZRmiLw2pHfRiewPKxZ/v
vQWluOdnOUB7kRXrwY6kq6P1T3FXY2XUJUkGIwH42niRxvmf4C++wWkWThbN2Y9s
yZbd9NOO5FfPmTTNEr43b0LDBt9r2h4rKkhAZxx/QrL26hDX7Xv+onRtWWolyzj8
0jA1vx2WOV+lRREnr5J3HMXmS47/6wZFQbaWfn7ZXIsuR2pObyAYRUfNwHQM+YhI
JFsL9W3oyEZUPIDFuJu+JN/NKq1laDT/kiKpJmEUyUBuvsSQQlUx3G69LxOqlmUN
xvYChCOvFm+U3KUWeNoKcm0ZW28CUoo7V6Xs16i/JDr/KcW18U9QLTqz/zu5de4P
sZxZ5BHOD2IEI1ksdVd/KTybTD8xN1FHLlhbsE1oY+xeli1VCRxIt5c3aGvQID4Q
t3SPeKh8oIxK58iXTucG1W1mCQTx6HXfbrVNL4H/qVmJ+I2D/nnsf7oadlbR0iYa
S4eXIMsW/Jyhzu8j8U3aHKD0j5MJ7Ho2ApV2MHL8F3mHB3bxiNcp5LwG9NM/a3UX
W7C8ryq1CCaYiHw81B3WbYun5/a1pRCB0jNN8N9vbCRH5TACtlQf6amtUe0pzRQE
fw6hNCSBZeJaJmtSCDC9PX6KllRBv0SFyM/PMqzCk7FJY3yF2SPPSFSLHRqat2n9
QlCBPAUfot6itIKLEFyptU3gBPapVg3mnAd7GQtz2mVdRSWGIwiqf0ufROtml51X
zGsgV0zenTyP4aWDfF/j0bDwXw7j2P7Rek/uvQJc3dMoL89zQ0YItI2TbER104ka
3FhmaGovtN4eh9Ilozmpniv0pOq1P0olD6hDtQFs25m7ZbwoE6Z7I1gfsxH9H8uY
N8/hVphsdzj/r4j8LGvDNwQjwKET8l4kHNRLxsfQc2eDVM+45m8iCM0jreARiprz
kKKRxz/CCBIMUCnwospfAVQS3v3YnFFai+5k4WM1Hvab6gs91K4/gWiAN4tnHVVY
fpI70RIuwWFQcxxbD5rIq/3+9B4BiAYt+oNVYwcwFYAXXxBqlZZWrS/k3MxhVLDR
qY16AAEqA3a3Kwvb2yFx4/Wyam4Luj4zQIYp7MP0x51r0Po+GLv6dirq7C8/bwhS
1C3cjO9wxGLv0nCO93yXnpeV3cFEJbZPfUvtCF3HkzRmaYpU5hif9jeQS98FGiqw
Vc/fuClYt+9sbn+lmAuKp/V5gtBx82R4wHFWA/34KJGQTiPbg11Sk/jDFnbCjQTj
g7ozW+CuyG1QT5DEhUnPsowtXnf/foqD/QOw2uBt20CrOpWDh4hxwgkKw3kOsU/C
Ph92vgejTysMAF4HF6RTeVdCG+9qKap7mgCrcFcitkAVitO1O+XnG5nno3MypiYq
X9U+JvXOObDxgZBU1c99uWdJMvXqZqDP2QRp+ZpYqIj3C4whEdNoNw9L+llQk8Ce
ELL7qcaiaawV7plb2tteyJL11mrj/ScIfp/CRfb+YvSYJaxuJgI4HGRK45Ijt6vg
YIsHsQCZvIEdU0BtXPfEba+rysVClDTUHG+h+a+TLEBR2csiU9hfCQzDQy5cF5ZC
ZGbZur0BTQ89FaJt45rhr/FYAUOwDQAUczOvQsASSNiEXO8cJo34UH5r7ZRPOcWU
BucXN/r95vvW7TT/S4DIB/ZbuDf1igFBUERf6mDwUKiYFcH94h23FMT2u6H26E1/
N2SijRNTt9BLFu3wjxqyIVlVjsa1Z9P4hA9lICOSWGsAvjGRSDvZcafqyXd2dd8k
kCpCwgmrbLGUniZVC/HoU4VVt9JG3LnOn38pslhGTNas1rjYJec6xowXK5yCTTXq
E/jm+nQfySmcPobVAHKv40Xz1cEvtR0Bcow9WG3Y6I4wQ3oOP9umEeegvOwSg42f
DJFGTuMnNqD3aX/9xOeLUaS43MMR8o/O/2dx8VBuxSPfZBcf4oetaIijrWIYM1Ea
X/Ph6v9pLVzT6nkPHKFXdEYqup3tCC4gt98fmJf9Hk/OGJ0QL2405OiyI9g1eC3G
E5PCvU6rBL0g6LMATMh+k57oxM1wBU0fL0XSRRzx52/I/VryuFKRpD7sO9c67i38
T6/MBMwKiGkTkIetw1t1QYuHe1AkqQehx8MmOz5ytT4bp1hh/D3pnYfanWTDFQar
ViSMVlDsDfI+r+CcfrtJPCeZY8dA2iGgmQ2s0RNdoP8XwsNBwr6bhSO2vJUUkNsd
CEGyFNclW9OYLD/X9cKUmdjXiLFVB7C1zmp9iDRqf8xVMXwLiRL74S+FgQt7gawk
gDRSaw/QuV5R+0rvURxsayGj714UsK/E61hYigaQ8wjba5bBG2RJMOOedGmb4lcO
tlnnnq4rZYVl2yFBByCZDTecbC+7U5m+gVaHy+OGHpE0oeYlH+L4HfUEGrRKjiRi
p6yyi0luzSumVFd0+Wb+m2BZkAnPkrzZ+pNdpd8A3RDTa1TVF+eCtgcdVYLLa2SV
1UdBnUCsZlOsfa2Tm0CKyDcyhmnQJ8kbS/Dr7JMkfaGf2vfhr1/6YZcrbEfvsCsk
6CEmEjJh30QTS5NQljTZgQNepcQ6GjhfZhhBZVzKwLgz8THn2LsB79Q6kRBigXP3
efr6HcJFcwO3WaTN94gqZpMc6hxDuArhUUWSK1+Nz2/96IVGB2iKAbYM5ytMkoyL
ebfdFcUS+WISxttmY4LRz8qq4hqrPafLM7elpyD75x3ZbeP/M+12rZGhQBsQ97zZ
aHxHFCmBxqT2ed2kJJpszx3II8xRChnfoNlVmFGVlchT7MInnbXQ9Kck16L/xVHd
6EDMXCJZCLV9ICMtVgWcFI8rDaBnHMrZFL68hpMSH1E2b9TvLHIfKE7nlpm/ocmi
CpclOocxUJ+13/iqNSpH4pz6og7lvCA3sWf2j4vs3m3I6wZ0c9WScx19NI0PtdrH
1lY+w0B8lMhGwYgnVO+Uu9UZ0OxWTAeHvsiW/8XZJo9hlA0ofMDFa0WILzroDBI9
t//453ai8Xe9N54Ht7yML7QvH+hcpJoucckJZBAx5D/kUVcCryemZN6y+sWxHvVh
1jSH32GmgLVgl7nIPHqfY917x8Fcj7zniRKBcBLzhQkppd3zfacAlweApZb1+COF
sjJiWRo0iw+Frhp/PdofVplm7uSmEdT3OHHhgHzTuA4UUa3kVgKO2p7XDwiRAl24
ujjyLKJJLHom/3J6XCHI4D4dWEra6LA5Qw3C66rqvlLiC1UkqUfSbh4JLKEcPWzd
BUmmOOrYLWwqNrt3kTP6bVN6sJfI8MRwMAYw6mB+rZhWWr5PW/HqMFMi5gRjacbm
6h1R0YnMSoGxHbTInVkSGtXJNxVezj/HtkKvOyKIMPrJT7fmTQGFMtUc3cJ0Fngh
34jyQUy3MZfZ23uwe7+zlBUqZ6WbvcY7215khoU/yRg8qg/dvs5zMYW8QHCIP6zu
8+N/9qAQU/6zBo+mqiBRSCnknLDObhQRD5chi6MNylY7Yj/PJyAG4sP6LCkLg7vu
nViZoK7rxoVwM0bqdcZOGEcrR0TD1MpTyjujOtBIKUoTTeXqL7dFF+NOod0e9VcA
FMmRmIQFLQEAm8iHIOpaKV9ZVw0NrZ4vY47jH7sDTfj0ym4wM3q3UX9gCiYvQLkh
Rd5dmv53tJaB3+kZTb4KvqSOfzyEBQtvpbqk1/lGVXaOfmMJ+dLO0LRDKuYt+EnJ
SI4QFkXKdOPR0aMA872R/vFTCe/mRKtl73KBxZMC+AfJY6ReNQXXZ2O3x3LrEFdF
X4zoPfQJQOe9RmZfn1PorziRrmznCXY1FLckKred/Qj9aw4Y/9Ce2wic/x142yJi
C1a3XrvEcz9YCptjkZD0MVz1fgKWTQHUJPzlLg2zLhQK9SwH5O+WERXQRsnA4qi4
i2U3NIrCsfOkptM8AH3wOGmsKsZzkpGf+6ecSN9qOFh58p71ZhPpJUgOmQqrKmzw
jtt0ztISuT69cINZ1A09iv/xuYaroY3k29Y6LFDFSBkssxy9fsrW7GQ+VWAIpUw3
wCqmNU+Vk8K54YUbGatlQZQGn3O5zdovZIWTZoK5PJPOvxgZxUXKVhf9CBpGKEok
qxd6tsEn6FRHV4Ug599u6iwLtzVmdXmBBi6zR7+lgUOrgbsKI3Rs2egwpeRqCNbN
L/MHB5gs/y1G3K5YDjGrPCJDakWIX4IuXAl33nM6/q6Wq8bByW913xqyI/nCGzJn
q6YU9/QkwXAbkzeKlbeLZbQ5/d1n/EzjtdMvgJpVAOO3tRnW2Ckr/5C0K4Nyb71g
UmpeH7Xc2L7/ASh7ZaFD4CxIXcn3RCS8gNKxK5a+/0ZUGc5QOIOxm/+38bt6L5N8
IW1o+ezz9hFq611awvBqdkYF5H/93X3YwAGQY6FmH7uGjo8ih6jTenjvooYt0fJ8
bsngB4siHaWd0FZduiTRBBGleUG1w0m4caOtffNWIKV1bsTHH59tdqUmqTBPXWwE
iJyOfWkkjdR85T5A2IcWVADwJEPSqQa+eD56lisV9OJhipyf7eKVqXNQR+y+YMY+
Qf4HIDcqPE+LvaeKFbf6/V0cMtAX1gAmGi45RvaY1UYdsgBO+j62zhYWb/7KuvoJ
1NjsjNhe+4pVyEVm1q/WzNhJTflm/SOrqLsMJ02swapfieMc/SNeSEYX8AeCngb3
dHhSHvqtu5utHlVlpdHuQzTCOu80Fcn0ssqtlBL18pUlc1DjloCX8K2nyHA6EFWB
ZCqZaV2/ux1dLdcHzijJEOpCwbPOIx/7+n/M95VEV9AJXVNHRkQl120TK8OZHREk
HKWftrQkfq3C3avvz7lbCc7KBubfBFAjptfYU1K7flvzpYmcEXJfjaJeP37zBHBn
ZZqR5HHOsJI2V/Dp43plEAN+XhXqYpznPpDE3fW9zCQs528HPzHw7/TzFRVVlWhN
YXtsYnxJayp/yRTQlzafwwic0rXu5rVTFidkzPRE3bh4O1n3i2I9jS3vXZCXT3z+
Q7+OkoDqsm8lY/TfFqxJFzmqse7umeAOh5wrIQAbVOgaVeg8jTWZWEO3wgp6yUgH
DLbtqXWq4hIiOHLVcQ/rG7aW0N7Yn+zic/uewbPQTZwK3gOR7gTrTN4bxK2YTvxB
OsXS1CmmzN+pdnRckmDGpozcaXeWHSvnkHNAGKEpW5JOTLyqZMtDT4HhFE9VbE1I
YjqLkMu6LlLD7ga80ZkHNArA0NHWNu9nvxO3ZGgU4hAUMYbx6e7YTRfB24vXk7NW
P1DQ7KOf98JwTBiuY/GSCF6gvYETUaBjW8rgCdbzumc6OimrJn/gTYS7eNeK6640
h/9i1XB/hd0ur7+3ucqV9gtvuVG3f/01dTc9h4ZYPJJ0zFM69TYen2uLYpN8jGe8
R3bw97WMGrDZqn8pfbsHqAbFmEuo6zJtMTRJvEa6rf53sUIdsQNo1/cEQMjcBDf5
u3y4lLoWrA3IfQ1yx7Tsiq8JAiwvY1xBoo6vmW6N1yk76Shg9ot37TnScuYoQzzK
zeMovqi8mk4T5CgapFGdjJMeOsu+kVEW1qPMgwXgffC7wA4P9lKAWzmJghsjDTAB
y+zMFCdfU4+Z4+9oIquxo6k45HNq8V3NbXu/MF9ifETntPAhpC6wKHoUvXB22JKe
LhBxqUN1wl5eVow1kXax4NsjuOARS3Fo1oNckiIaiWs958GZPvkZtuLmJDfNb4zY
LfjyQ4upvx8dugBN1FdEnVaBtLhO2H021KFWZEFSzceLZ3Fed2go/ACJa0FyRTZ3
k53qSs2fLAR2jqepBNzGrH+ZZMCFVhoh2wE1jWjvvfJSprlwPzWsT9sLptsuRoSU
nYUpqvycfxsk1iHlW1f7J9oykJv1KZ+s6740iUu1JCg+PVlVImM6j9MlsaSJ1CP2
wF054Nxslf+YgAXEAL/dkDsPBLOWYZ4cgKdpJg9Em0d/srCN0CP1UVO0R1LNIx/Q
c+cYtDyAGqL9ylNY1oqMjhV97XHItJNB1TXZM4MDAA2vFoUnsCQRIZ8VE03UXpFO
Q5J1Lf9Q4FKK3KXaoawXDkBjYim9zUKOIEiIiQIXF8fFD+qzJmdGQwiD8BMhaWQe
6inmX9ZgpH/vKttPvJ56/IouUCIM9iAYegqO7tuacKWAnNKA4po+mE4t4kAvTvIb
4h9k/ju1C39h/A7MeUS6efVVH/nkKbuKcNRYZNj/ACNAGBHK13c792acSJgRSlTP
uab7Ng8S++ssfb7ovi97F4ZiHXG1s1xqHAbMlIlZJ0IuODpcCpBKKmyltxYGYFB5
8cCBeX1zlE7guMZHKcbF02fZXYdRc77t3u1ld5WIUdk94aBhrxLm5QagKfhWrgNs
bAOexPTHTHmuFIBMJEfPKcR5dqmW7UodKBHxvSi1L92uS7ltn8oXGfc3C0YQk0ps
p7m3u7MmSH9TH1qWCSpUf7laGUTMLqbkSMMwjyAV2KARseum7Ig5L/UJhd/wM8Vc
v9NUPMZ2jlN3wppQoypwVn/UbhJu4f/55V5zU8EgZ/2Cwo/wCRjdq203yU7jG4Oi
sbtbHFRcdpZwdMNI75QFivUIrpKHFRthmC1h1zpORLHRhQHPzCeU44Clhsp5+Inc
tfllSkx9SB8s2BSv8SOx+PTbxUudJkyFx0C4I+G7GAqwvv4uUOYlDGAJRsnzoNZl
dTT45cMo51J+4Knoq5ilRmfXS/ojFLJpPURM6jViSw4vMJ6GZDnUFcS+vB1aKJs/
mFjinfNBQPJmA8NBjt+GMkeeZlRCi/GHdhAPUVJV5PW8/htMUA36WdbUvVM9u72J
+gOZBaBtyCasqU/73AHdyFMASEvsJS3ohkiXuAlIXAb9UwbpZ/NiIny1cjKHdZc2
Qlcuk29KaGQHXVaewda+PllPkzyLiBMDIrUY0GaRZJJ9U163T92VOo4Qyrbqy5HA
8CqtslXzok9PEEUdQ5aXGjub+u9e0Bt2KJlk0jxqVlSWTWQArWMGgTxcitPEOQ5L
QLqOTBeWs0oOH+/Vah3jX+2FRvdhonB5g59NUsqu0jGMjjV9OqYVhFFo5Q+5MAqL
73sYYKNdDOzLWetG/l4wZAFbOr1pWgyId7Vngn6Y8v6et2qJavtMuvRWyBMTsnYr
TDBfswD6hXfkrS365VlCN27CkazwFR7NML4YKhf5tmmU3/NQ1E823CUesYkR5QCa
yGSA2NxWPhDwQpfVqrmOms/Nr/r+HWNsRAwhXIJQ5cDk97VU+g3e5HTZAXgnUN+T
Rky3CYQ2e12yuXoHYbEH8f9VWS7BKAPuVWsj763ZHDzn3rE9fdFGc9ux/aIBJnSv
dbpEgnwmR6Xg0j6LLcaDAO/vCBjbbFwPl/1yBulKuZr/zFrSNLEygCQ8Rr0oSjXy
9cyCBFRJ0huESoth/kW6NzDowI8SSB5iZkGoYovn5u3apnVdFvbitBUIUR4eFxUQ
tX4M65Axz2gRXRApXhdIUPQobCM92vRiuJX3/88X59dAi/j8OjsW3ib4nw1/eARY
V8MUfVSUXuAo5882UKevgyPskwsFew+xs5PVb8UsWfplv84+sW2uS5WAyCpfhIrI
Bp9EFXRChc9bC7S2aiJyLUyGmlGb+9qcy6G/eSCyD96zVzK2nyuGE4Z3tUuBkBhx
49tvOdfTrWXi8PKfj8awyYpPjS9LfJm4mdSLoMx+fHdIeZfKd+eri2IF0KPJjz/i
z/uvowlCME+8S8uYojxp4BjNngULFIWVbiY1cP9Vl4fA+ZXmeSIPnDNlB5HZYZLK
kNl7dFf4EcW47MxXRMoQHEK0WaI8P0poAfAFxKIptVFpE01fqkcSHJS0OvgXBc6l
/SY41G4asrhOJP8joc81xGur3rvmzhEQQMkDTysvfcGZ0jNlDC+V9lpYvL0C6dfN
MXDDRfV58+kyqCD7oEJGgHWBkcJ8YUeDdNhmwCjbz0sCTIyXrClQytQ/3TXKsB/1
XCggIl3iUwbtzZR3noGXvq+HqbCAVkmi0TwhlWwwBlPTIJYHlxV6565O77pi6DPb
xRihe75fQo1NyUEbvioGpGRK2Vl5jSu1QfOEA7UguJ9K9+iymmnRDxLQqhRC/5FY
p9ngkK4KltYkIamanl/Kw7WwNaEmkkHkgZlSLkR51TNyklb8mxMCyRXy1TOvSHun
inYxMDzFm4PP3bgF9wAIWy5gAkKgpzV7hlueX94gLb6UCfo7ac0nP7uHNZRiBHN8
UqOAFm2AcdazKYYxJH/JXbEt4usaP9tjln3tTMWg3H4XMhgqevc7KUK6WV82+/2p
AK5OjkG5waTwueIbfZzOvhKazz9aJZXDuMZyGtll74H/WqSC7OnpP995y8QA8oST
98sqJWclRzMhC6uTVZlKBy1HtyNia3RGSqS04ZHEdjZhGmSAMdQKy44BVxKHc2wv
T2mvAPjs1RyD2UiJCoODTI1W91+MgW9G98kq8K4wVSymSqfYfYJZwW+RJHz9MmGu
76KAxQ9Y8p0YLKKegIA8Un/oyUN2RRekqLwLjILDVM9eeHiBP6lmtFD75WgSxUr+
gsKZTt78aH9YivJ+oqWivhVd1j6x+2+nF8Vt/e36jXtE2Uq47ID0nxNThPosWwVv
gVR7TvCiw8mYEjWTxhaqjXv3T1+9WIrhN03QK9xSrFL0nHd6Pnr0ftq4zAG3h3fW
QGSH02tf/+TGpjC/ytDZE7RlVmN33LJgjFrNEk0L6h5MG6L9s67KmSEqKRCJomdA
D04Askm6Gw98HN8QtzQNPzm67JAd343UUgI5dxs7fhPG6UsQzfCwhrry0iLOyRHu
M2L1cwfTlIJPifwO1XWl+29Ub/ReEVnRDjOvkpuaa46L8OhDl/gnFiUTmSsyv5uE
wOmiEQeh957T7N0IcIK6ZTRovjudnN4ScVeYIlesFu1+uw4pN9nN8KParKU2Irli
43GUxCfKhQnTjGU44xHWlssOb9xGRNz+QTfjYj5P70LhuZZSsBxvqQIwt9uOXDCe
mMP3VzAws5v9WFIaOGfuRI/6I7/FU0QH3sOyUM1a0Lip3XJi8KhY4175/CfT4FTF
cq7DiN3v/bTkujs1aH8lfkouYQ3rxW4V1xhYbjlokhHlgrsSEXGLKaA7YhkcnHPn
AjVKyW5VVNASZia5gVrxzvLY6YVatvtkzbZSfzD+7C3rCKTpJaq7aHWoCPlmpdsc
tAyiwQ+G5QBncJgahSzlM/Xd96kurd/rtu80lDYSm0jAqdmB4//B7w74rOSEAQT9
sfjHci97DoBSuttY58e4J3iIx+1U8FpKiwU3T9ZD6uPv/HxoamMAf/w8610FSYpi
4RHAw8Fuqqazp2AZUDF0iQalP5Zxxf/dsBrOTH3S85c64KKemcSlDoeNM2QsO6GW
uMYmt+//twbh2vdemBWdTS/BPaF6Ia60RNalVv57tQKfnIQT8SI+UIeOc6DFVVis
iKqG4uW9E6GTV2lBcKYeP7qCI51Qa7ZpGkjBUBbuascgHBcfic2nMdwgQNW8qnS+
q/f57QzMDQqVs+QRuMHxw8E3dLA67s6EWrCM8DJZdgeDgRAbhUnfXQ12FShVsfYD
+xsiXZK6u6DIbiOuky8i8TNYQueglSjvVfa/GzmyMrcae1dv5MpGgx0ycxl/aOQO
pueVQ4Yc0ZnE2Fohaae8r3gAColfdBUeABIRW9oSiHSQbVj6e6PLShD0ZJq1FJkN
Bef+QkaTdzQ1yPxfeGm3yziCk3E+w3cYvdQr3nOUEl0uakrKtJlxmGWgi8PZq+cD
2unCRgJAVkpSItEs9eKHL1jUkdhrCGUHBZmNFR9MzqptHTYxoNPtHNfLo9IHscls
9Tl9EufZxjf8rP6IFQREbCJrL31A11203a4fLdbUaWEh/e3dQ9CmC1DqwlrIVrjJ
Eq5omeZamH5iHr7er1zabOW24RqLVpyzc8WygBDZwOIUt9ZoJJL+pOnpI3lOsDri
OQ11eCOjMpiseb2hnOZePn2IJi5w+r0L2dMbs7FEG9XyoaCp2NjYb+7Pzdbptf4k
CZ9CLnGI5BYcRifN62KR+iWzz9PGnbGvZQjek7CfgDF4lhZLFAClhTdJeWspNEuY
Yr0uCgEBZH3QNqptlyEX/5XV7famHdCegZb8lnW1vQTSEyRaZRWOt1ZfeP7wYFXT
nvn+lN17fF2ETX0yjWjbQbjp05IB5RWZdag+ZODlklHAecb13EDx0dq1vszZZcOg
cM//0AJunXFEFTwT9Ahn/g13JTMZH70UOvZhMyfTch5ihZdYnq5K2fh14wfA0XPn
d3hw+mLdQkZ7BusN/R+ODwc11t2maYWoILWtUWWQ0+5nWFuGNLgaEw8NMIa1iByk
9IegoXULl1vVgybakEUEixTioI+QGnyENnhjJ5Q1dUd1nmzIBXCImmYEwQarWV5f
DOGr1psV02wF/BfBAN6w40yuAwQK4wfwMUk211qmLq55hx/6+vkHSPiO1ENVdRfm
GVhC2wIG5+p2CvBPpy1SxpY+UGgu2tsDfhvYESuoNM4ghaXumDYKYSZku7WTul7x
ZkDvY9Pbu6dJj57sn7i0XMCgnMpVgq+GiN/kH6iTCEDwU9S9tb3/tsdeBLGJ6P+T
HxeRc7vWVA1Ghj1T815acG82YZBPbyIUfk5XI/qrBpuAfrxHR2DwivZm5+bYYiah
Jc/biWY98s1rew72Ac29QSEZqA2s6OlxZ1V2Qpci8ioAxQ0MnRTHL29Kzki0EMwv
0TD8Pd4Xt/8UIHdYd5oivelATGEUcnok8q1Iktu78i/K9fPdPbFmrLTT9lIrWQUy
39E3WW2azU4yH009gOIKX+oZ5rIF7R7Y9O5Q8NbbLiGuCQW+LqvTaF7fFq4ceN5s
PpWQNUTEl0PEX/DKnapqQenJ+MxHsE247vVs5rfOpla5ZOprBcLK/a3drUgRWxky
GYBbZS+UZxg2o/v7Llx333Y2lmZfp7GOvkY7TpmOKH//Gst/zPf7xEO5EB9FKa3L
XH8ZhbtIvA/HTx3PWqX/5Tax1yCWOizMhNF/3a6UQwG0GNIl3bD6sqBhQTu+hqaH
zPIGyx7EPQLvTLtrClABzo4vFDajqFq/rbdJvy8+A5Wm7XTltlQOxPix8CmMFCzW
v/b6frZFtxeqqf45RwuAgDDb9egxt0NOwKM03bepY7appUiOOm0B56ZSs6MdsHLn
mymSIcqn3nzGK90S+5Nfif7GITCMEvqUbGmv00717Iki2MoSApd4tE3CYcufNPyP
hDT1J0NhpYg9QbdOOgHb/IuEl/fo2DPx25IP3DvJ8JZ5PMfK3+1diUQzHpp820SK
37U9H6LjzGT9lZTmf3ypcUGKzz2gTlllu6mM4IbHO40REKPkajmg0LPXrsC+WWKq
SvEQL1hScjloqsQsyXOksiX9tm1ETDZSFkv22IVKcplNrdUYgDQaF3qTP8BcEBO8
lGVkN0AdOLtJJaN9L2EGL9pRWg7viLvh1YtFljXhgOkZN2hxNCkHPJ5qdkl08gxI
v0kbvMs9FkNg9v89x6sTolPeH+lDos3NT4cRe1mvFwu6KSXb5rhLZfn3vQxfjbzY
Slcvk6myWnhHTcTMYe1qxEwqgUueg9dZIFKGPN03nYuvWM5fAHagt+bM17IilgB1
rHC2xk+FZyz3MyP+jvkqvUJ8P68zTDofL9q1uEdP+StRJPV8v50tBdJKSHOu8Mtx
Qd80EJw5N3tHVwk1eLj8yknufYSZ4U0Z2z1OTXIJSo5PbFRvfZq+Yn3rpfrBF1Sp
TEFRL9vWJttIRgwC3YrZTYiUllF5e3o3dYuXy80Dqhc7KebT1NNRIivMARfCCIpL
RgNwGHfOzE6ZDp42q9FHIyxB9e84W8+JHxwjsAW0D8i8gULhcOHvTwm38bL5CDHz
MIbcPoORZgINh07kppv7WB5cDsW+8JMCbkho3LLpodXu9tTgBz//9nqQHafc2UUo
vJA599O58/ZubDe6/Yoqf/jQcs+Odnpc9dlIKPz6riWMTU06StPp4w0/sXcJ/ctl
dfeoC22YDqPzlRqAmYEvLUuaIptPvjdHbV/+6VjvNDr19dNf+l9k/RqWgUS91nM/
VFZGNSRBSEXQmWJ48qOnKfHlQB3SOrFMJI0PWWl1Iyw6eJ7FCnojILGfcLoA8WLO
Lqtxb4+JumtibrxvIuNwUzK1W7HyBzCVRD0tg4U9HX+Um894zkV2sm7eJ8uGBRKF
JMKuNbpx+zG0ySpKrdP/+r1HmEEdLR3HS6Z1wdn67tIEOGRZP3GX6BFB6ASe19yr
tVXwClr4p9EbvdNqleczOz6Ix4FzCalMYHgamiDvd4XecyD+BPafVw3Ir6RSxp6j
biBTniO/BeCXTJOjJ6oxNLl/YhBjY2OzfVipO1huYTk9/Jzbjfz++NkaaRqYIb8t
5oJZOwQ0cS9zRQcHJIqodV27Jgq5yNfCtISKFASkw1AWQ4UR1C4XXx7WEz2iHvOe
Jjl5DnnfStCN3pGrkWtPYgowSpLUCj7GWMKExGMpuK2EIWnHIokApWJD3XyYBfob
bPBKky7XGiJlsj2PrXnergL+x6e26AyYDShXBkAnOlX5SrfqIaZwGb0SNEs4+eWR
9EMZyHyszTk4xAaPKzhUBJowxp/7NKdIRAIEtSCbBd40DPDxab/vZnS1pUASJ1BA
DnnC8B/Aqhi4UrEAtPE318ZpME01hij++7QhfE85979nnMPW50lmM+b77mDCEEb2
3bKpJV0N4S1EM++b+Z5dQmHjOhFz59L+xuS1zCa8OuYOyI5/mQpTklMlKti/4mKu
he0TsDmgmgCsqCVJCqw10YJjFJ+1uB0AA1+D3hemRqdO5S7VH0drO4zW1e78mFJR
En8Gl1L8VdzGceSxhJChzdxHmkd8ToAb1DFERChZNL1i/PanyMYMI00KX2j+/Ral
NpTwUd8BP+LEvWisOpDjKfh07PURQwMT1fslW2iSSqsEO2fU7VczYEn8xZONJ2B6
zqCykWpIxv8CskbVqeKvCfG8K6fl9Nl4clnxiihzBTb6FCpCtc9F060S9jNXAoOP
7tf2XiD6FxzS5qbbpLMsK0GSTvlHijfWLUeS/zRsWzp+3P1rnggzaACmu3hnR/VU
YBT/Jl8wXSlWLZf/mcirZOe4ouQde2qZCx0Oa+BVzQ9vhdRQyJx0Wtgfn7hU8B8z
8GY4v/AJQLAmNaRkXn5PMOqkxBEDG2kaJJg2PH9TA+xmLqBbmUEXgthZi3FBoKPv
/hhNS1eZyObSGxqy7Gw5hrwMYq+sZR4+yk3a19OL4uiaGQPM5LURej6ZSwfstcQ+
fGlsnNBTIc9Nzcwo6eyqGhPDmcwMFMd3QVVPg/Zl9clu0U7Jd0cXyi5klOvXJGQJ
ShKZSc1jhLdc4uwugJVxZoOB8oHUt6TGHJSkaJ604mZ/zTf6CWCuaO7ww3bR/JYh
25KV7Lz6Rh49fUfEBUqaqXS5NJRwSki98he+hEoDkpCT45nKSjfOMR4XsqfqkAaA
6yNJwZMCUz/KFfaXAtAmYjVB+oomFv0OYySSTJG6RTNpWl36Cv80bSPNkuRnc4G1
i67YukKc77WK5QHNXYFBV9Se9mR7SRL55UZbH7wRraSva4wRTQxlS5DifkVqDo1g
TKAgB7X8Y1TFJ1PWwhTgfSQvvZlkVSqAiI6imo9S38dUB29OkYU+GcYzO1GP90F8
KP6nVL7PUVFWi6UiuVsbN4TyJO6AJdF6j/aAH9mxk1g3DHVzvFooOMdGiFwHk10E
TqtAKcnLovwKhVZG7PgdK8Kw0vmS7o79Isc9CIryM4AxP4XdG8kHWbg9qwl2hdJ5
L+4pFwolVT7DOdzPTOHBOPCeMHXxdL4hDq0j6rLJr9CwzUyCz6Sxq7o+On6u3q9Y
359kXIpxnnROkzgAXj781kalAFjH4SkDAQ2G4mNRTD9jHRBIXThrNfC10nCeLKTw
PWanb3X7rOqejFV+wN7Dtd7X/b39XXnFsELT6itUGGcSAPHuGGfd+VFtnWdgxzLy
qGky8rpVF8a4mv6DRjFDynztTxlRmRYStRZpMtuv9mz3J/1e8XaejEJPVs8OPxqe
+UUZvZVCgpcsHgBu9bcIwifbCK+ZhTAGCLLBtKJdmdAf8LT6KeyL0/9vb9ITcLah
OquLDjsO/tJ517cA8U7AEftsFPDd9Kq3N2U8lcb7b+fiHRdPlfnTaouCaPGHGgZ2
gPxzO9vp6mMYeiCOYzXsfqTpf/U52oTqOpAaZq+lsnUV1G5ew1epG229y/tj7nQf
YQQlE0efFGeNujgJJBuGyqPMh722DEQwGD8MT6lD5gfJ5da0XYVDZGF0whVfx67x
5TfNsSWqDUzvMGPiStMNow2ga06PGE6eO8whRtydRxUTn/ooslywEWpwzEHphce/
DvmObg0L6MdHyE/Vj4dSO4bf9oQo+MlZ8jUCoXWt1LddIeS8OzLn6SYrZAc1e17H
gBi1bqNjKKXqbCYr+wUqeg/ezllWBvFryINrm0HTPQ8CsumKrwAFtQLHvyeVC/l+
lXS8k7MX6uRg9sCxPk+MJ7LMjLBQDIoTyHR1SZggUbs0DbC+hbMkQGbgur0rXJCl
BTOFT37xw6eqHzfWZjOh0Oy3qg/sdRwkRZOkjg1IIXqfhoP6TJ6MFt1ladIK0Srp
VUCsM2nGxOOTYFQT6PUqz87VL6NBTtlHofR5/MwiXoijK0N9N1evWObGsCs1mhWt
/eTtgtIpr9jA+CZBJMfvdjXYWwt2K6I1lJLmQAYxp7srifr1KdiIODpC6D8UprBP
Mjy6R2IRplSzUyDeo8uV+s2qddGlhRBGAsEs/ltk846zn6+0jlicqEvKWhqRx4nn
Dkkrt6KbL/6QiO3GrdX9qqN33i60NkKXgRx4YxhFwdw8kesnDB6lPM7qEV7QHLIn
+6CoaetbvaDA07n4/UrDV+bfw0a3lEL2BkIK0tTLB23y+z3fWcrFcvi8RHi+tZ6I
Pb/6cGb8PmkfMxQ189tfdIsmemkfktxQKB1lAW2gngda2P532LyShKEfC8NZmxQT
Vtqx83OzubyJddzytMAaru7GNfV5SBl4HxAufyTzcMdGdIvcfu78mCSiFxAT0BKL
7DfYHOrN7hI3W3BjE79bT0NAplj0yIB1TZaQ3e12JN0yg+JXxdbreuAJBzXieUFo
QRrj6lGxywaCA4Qj+JizbYTvkpElS6mywAyn6tbNf8TJWKO7kR6XSg1vyrSG6Oqo
/RhxEqd0SUm3pqlcmyzfModBDZ3keoiVrU/EXP8frCZKP7AgXL1+B1VB/Nq1t15w
/xiQJK9nTgbIwkkjvZzqgd1xkvqu14qGMLEYsCBI2IYycHUzeuDfZYnD+RIg+/RV
6XVo8jskiPWpykq4JKbhBRByTF5zZq8yDtJ5Re5StXdZVUWhOJT9y9JjH8X6AooV
YH4eAOGUyAxwsAq6GGgJ9ups5XCJw2losymQKiQspYftPirCXvJwRrmNu4mtNlK5
pG+q9PTb6SKGzDy59jVBZUuQ8xHB8q3SaZVSdhx0Uym1t5VNP/0rCGz47cpX47py
vQaMgrKirrvHFXIMQzFONB9ljfy8IvsWWe3taTZfM3Tvp2YkOONBN275u/UfqRJo
xq3LRiiFuPFqYApp0FOiUE0iacSpu4LiWArZcUYv4/rM5ZywYgZ25AN6bDaFMQ1o
apTX7LL8szlzenlQY7sqUDUbGn2+RHsXr1nQniJOgfKlMzA81hcV8FLwvnzw54ie
w2xM3a38F5lisi+3OYlwSzXNvRkyhNwYr3gwiAEeYEcfrsOBh7/oad+0FBj65u7O
HdY73bCndFSQQUnkg8jLdOgsGQbTTCSzKE19HnYdQVNf0ziXvDnMRIetLJuSvhTj
jaw9YH3h1nNhpw+fn9e2a64zu1FPD6heUwURnJAp92Brn+ECFKSo6D7IRrxn+T0Q
VBeBnHEUApCmhqG5oeA+lPCcWghQEEw/ZfWXcmC5uAb3H1Enz+4I2Jsx9xa68kDg
nqRG21xMJRwnNpLuiLJf1wt6NyNaE2FPRLz9/cEvweSDTwqMMBdpLEIKBQQxKMEn
+IFtH9lrLhTE+/fnR5kJchr6HMRlmVUMyfB2P2wZpW0rx6L7563GsKkMi1/5nUUy
6yU3OAXlQ7mguRkml9RU/hwt/VidTOFoSD51NdXWYn0+sdZNhHHtsEN72GEYc9yc
q0HF1i1aWN/33bef1C5D55TOgOo6N6fGyMrA/u0m9KiGkFgcng7l7+dD1CmL9TQJ
E0NTcY2urEiVdbaTiDfMG1XJQDSnRHDTvCL1gRh29Es/OKPRVUenvnYCY4jyLzpk
Kt3IjWKwrDGrK3BbszrqPvDLCAG+N50gnvxYQaJepHo+WEoTVtNQgPA7dxoEw+gx
uTa6pGGNcWeqtD31SyGf3ZiV7tN1+ZKR4AYi0okWZ7HPCBMukhEupkXD9MS/99vj
RR6iUV3tZptfs/HICjWPNDbEAl4y3N2bo+L4Z5p+ze2L1BBjZQj/H3IabgcuxA5B
kBa/tmMgZrjwSrfsHakrnnPsdsdDXfjviPup5oVUiUFdbRWSzZIpjR4aS2lzzUtH
gJyo1EuWjwvLPtf+RX7Xczke661qpf8bLvBz7XixlLCO9aEjqJFL3+pvg2mB2BE4
mvAO2Eoa1qVMfaaNeGmN4cc1lD015FwU4af6SFQdMlAwQOgVsevtxmxRSO7MY+wj
HVsGg+ZrlKjCXSd8vE/ydfc9ZqANwzn+BeZvtVOBMXeLkuHG+djuI22IplO0SJlm
4G/IrZo+hQ2o6XvWuij8UJAebvJAkkHp8K2oaygyPvqwHZMs1A613pr5YGOXHJdq
p4CaoESpj5TS7+L/Q7Q4Z1cTQ5hKobSau+vr0EASRHlJc3XgzYjnENDZwbljgRG8
bf51ZrS4RLsERnG9F96/aa+wr+O7asiJJAhO+H39uoRsDJqVE7fvUe3OXIuDDfU9
WZTZBxAXMJyPJQbVF/VTek7Nw3eo58eRCiR8tdGZLrE20SiQMZyNkHt4rgfLUSHV
JYPAaFj1izIlJasmUa0IjPvPxztHtTjJa1P7Iu0oH8Nagr+2zD4wOzhVHk75JVB7
YHX0EO6TZYBWUobK4+RDfTgdOtTRF/cKfuibFhkIJr19U1DXvWW+PlEx4fv6n0wW
hpoBOuXo1Q1lHQyLTFN8rh9xVRcs6lLsCYXdFWFPyugKB2CT1Cdp4y3G2qWTyRzf
FeL2LOKvTMcnSxZl0m8Z1Drghal5mvdr5kXfUdWKE5mOSj3aPqlofPWc0zqf1se+
iubbn5nGUJNp1PBdJb72IEfeB4OO92AfIszBGKKBO+xZLYdyvQuRJo9IuTvSryv5
p0jI4klcvzc2oAKc+woRVvO923D2yfe8VFjP0p+vli3xpyKGiP1qDC6/C3G52ybz
s6H0eeSmLpaDFaDKB21y4DWn6sdEcsJY+z2/oEsvhLDor18O94ZWEJ/6AG+l/oG1
ZyTOArR8Sfle0eYhmALUYc1N05grDMjD6QMSmS7xnqZdg07yb7PiFQMI/8C11ozR
7V55zbMZfVb/2SoW4EZ27gAQe9LPVZu/cavM5qXYz2mBOaCmF1SPRS5uXg3BImmb
Glg2g2Zt3hiQ3x+CunJGtuAPIQveyiFJPg49geERzw551HR0QSr09tQA+oSdCI4E
sv9Aiky+Z2i0fNKKAD46Z3W72f0F9Qd08a4P5r/z7HGg/dEWwVibG0k0sRu7o8sg
JQrNeXaqV2MyCCFPPBSP1XyucZdkfgc8Sc6UDzymDe3+e9g53or47TJ4wF9uiUhy
vC0LOazTZAbV77ltS50cdkPnxUrZoWc08KvnvKlEX3BYfEbMf6Qp1U2I56T/yGMz
GTROeklpu58O/Gb4B1fPgRRJZffM/WI6EA/5x7OflL6wOms/i2c6xI6D5uL+upr8
ZeEtN7osdIufWvt3vIgxJuQPlFeOepYCgGowRKCh8zLhnzp5IBSiNxhPi/k2jDze
oBim8lWlVh1oufQ/83monHxB627f1ouFyUHH9lDZi7crM6g0rFZKux1+/aDgBUos
gl4wsaeTm3Pa75VI3x4L1+Q48DWq1VIh3D22k8+yDhpSd9QfNFzw6bL6WIvKFq7m
AGY+z56ViUh4sYQMC2v6vUEudMLsNXVhvK2eayhK+M6KLTPBvpspMSgVeLNFhoet
L4GJlL2IIrqokFXpjjdGzFO1DWKxKQD83RWf+vrnGL1xbIH/pGwKx8o00Yeswlr4
8KrREAvIE4TeZnKseuQvwYvJZr2sctpOOc7kscJuxQEYIUubTbj/n6iD2xlhsqin
6m+QrfbMwkB8GvpfpZBQ6tDAeAnx7kObkZ1BcBWoYqjEoALPlwJcOANhNeyJAdz5
YLjoz8nW8WlfW2Ki9kRyuci8oW4m5zOdAZ/gcZF3pNgnw23LabdHb+NgK2GagkhW
nB5neH5pogcZZyP6lCHNaMl5vKPX0EClEHUet182E/T4QifZQCaIAryCCJNcA/7x
34VXlsvXc1I5kT7q26GW5GGPlt0YUH+nZKPNFaXtdtf+41n7/VONFMBMn1MGumBz
NOaB4ktHMZUboBo/1vfM5AcVIYDM0vcK1YFGXA0QKeLUJ5dyqwZ6d7QY2RZAWeaf
bnj3ud2Se1aXBVRqQfryFAb4IYjLxBUJVQai8YuZ7ry9yLd5ZFhaTCkQLJLyg6Qw
/Rc298PeNwbmM92PdqCp8WswM9AU0NNvD/BQ5TcA36m2aUUwh2ILY+/18S+9/2n1
AwntSiO9SEOBkyMdQoGpZkhyjmBi1upeW60Wp7knhHHaHHmqcdUilBgiDY+LQ/Oc
u6/8kuVCQLTPbY5sHrCCXudtP+iH0UEPGvf0XdYNt9DPALn5WceIYkofkuKNm5pK
7A8GL9GKNE6JQWSVWNEGCHloYV8lQ/Aa7Sq2CNZIpheOJqHHcjeukraAwKGcgvQk
xI9FRphm5NEP/uLBrkCzaNY7gPu/nSnHE1DkSGDiST23nXwYpbJMzbES+FPeTjM2
MxE4C/s3xdpUQQxwQ6Mv/IFYdfANvtCW/C7QVBWB8C32vPlCf9cZOuV03WltOFpm
giHYiFM4AmnrrHUOKVfO5jKeburNFggHxQieTy4HPmx4cF8ts2iFXQZDVv4FLyNd
whzFuZS9Br6xyai6mboHk/M5AFvUCYcAEkxmH8T8G56fXExnImFaUHWv6KNQ8ial
9bK7oLxZx41jfGOlhwNEwFoJ/XgX+Ml+1dW4r4hxCG8fBjEvzS3CGiQHokFQpl29
Wdc/I2t15yUyNISeFaIMqzG55KSANQuWK2Fr+7SSfA5Js77zkSOlArosO9aFCQeo
ZSu35WUkdUa9rnhCOILA3Q/WXYMgKSd8AeecVt7GZImsfCicplLcL/syyLT8Z0h5
RklurWts7zUAU459ryHraH/gqSvknLGzY2P6yRM+BUkD7hnn9i68owMf4BS1LzR+
MNTt5iwD/rzYZ4q/pV44WERbvkc8hebLjsG5T8+FCCPLQUWrTPjC7qiZOLgbFR36
ME/mcl30+ulOSdtz5g4FP8HRXCUUO07oBlCEeW5pVGzwHJUpiFnEVEfXwhNOaD1c
58ABfEhIdBOVUNkaitbXVCK7++ZiqSd4DT8wUlPtVq2E+w9t6239ZiDfOPiUnhGN
AjfNJsdhuRTxwTGKr2hEaGS73jzSxdKpmxf5M5k43uUtqDKqOBV2MfdginKP1UMg
gZHa9N5wDfosHRKXWvZr1n/xWW+aNzAiFWenzqfqJ/XJ9DlrtinJBSE6a8cFjZl8
kTXRlRMa21QTYs3hHUBj/f5hSUp1oW8UJfFuBvTu0c1ZabDXJQGVdGXS1SzK6m1l
o1UiQmbNREo64T7jocGAQrofJl/L3RrEGgnjNg4emq6BdkkAKPW4J/+ARHph64pM
hFxf5WXLgPWp69F40b15Ljx+TVuPIfiVxyzvyDU+XFO6dUZd/v8Kmo6cDxZQOY3E
HbSd8nfXNNkzH3qNVkdwJtKKx1HpkpzMKDnAV088930/R8anA4OwF5YWfJGpxG1s
0rmaMRIXuSGT/oieBi9PZ0hvEeCbrulV1wKBmL5kiq/lhswXe8JFzE0XYow76CN5
crZY/0cB1+7MZllgNqKTt5n0WUqE2l4rdbnLGiX0r2iiPI8AkgMWGf0cfLOpIFtD
1sjkvH9xaZc3k/h8Ew7Rh2VVoxFl+l2KDTPTKFKNIltKJmgsJzj1uSbf7T1Lt5dQ
tTEy5W4W41wC7ebk6dCxB0SVMu5elG5idODXUIc5TzUKAngIFKzfZ0XIjUCPjVZ/
rwKZ73ok1zYIL9nCYs119Sx0iIDLnCjlSA2m+dN1ME6tUSmYI1Lf6EzXJPdYX66X
G/zPQqrgKQoICysPIyeJDdkIn7lUNWtva2gvJE2PEdwVbAlR1QzwZJ3boIgQwKQS
N01mdrdQczfyvkQY98GDwnbKKIM3/64d7QA13Lkl0ho/9JOo7NUeCk6K+i6HFcln
Ixei2LggYHVbd3JFBT1n4RS5wQIMuhYgCd/oRTXA6dkObVaGuLZN0uXWhzfm59Q1
SKxr+sB6mY8vL4jWJPUCwniqpfWeLKpZXEYkvyaU9Ov5ZzQwB6Iw68tJELqH+jxI
LL02Uu6nhYEqftpXYzFJx7lmPsLBsiu2sc2c+20uoBLTNVjGfn4GNmKJxgCXvew6
WiOeU0pkSWapzGYrC/kXHBbuNTFfbEjSwW53qQkFWICbVUrX+ZWzGv02WnEiaOZY
8cwLWrezv9r23/iMWEBx3eMW4PDrK+JP5YyEhjiBu5YqAF3rKpFVTdlgusFRboOV
V5jAXoItOvncBKpMviTaAEZDGN8Gl5ODFK81/cBjfpgjVxc52igxq9mowzjGewzT
O5dh6k/1T2Ti6esNcBldkL85xreK3C9fOkjhTaEKE0uMHE8QaKctUSOblNJUJ69g
c2TdA5NLHxGWd8w6czEXop162Nmbyn8GzthzWVedJi0FsPsANoIq4tU1J36HBWLK
HO3+mB3JVayGWinQWkX3hcFEHTjB7oFOHEilPwXz7HS4Fut4KOWVUzdQXfYj0bA0
7NZn4tXDq2UJt/pJTZWv9+A4eqQpd/XBKoU5eu9CW567gt6iWQqVygWyu1JxWAXH
+alddsewQ6aTnBgv2VRtaLn3sSPq5aPpmdQkMcZUdzSc03sXG4FGZkT6ddjZtYYy
dQCRKUdKsS87z6Tudur+g2saK1j0iYLK6PMrvIlrKmaVvcNh3zvoVjvKvv0Q9a71
RdNAHbgwsP8+HBassTl/BvW+lDKMv6V5ujNUKiJNsfszv6cBicOHFB9c1Hpqhfe3
KxAwGvf8BIF+Lz1n9LfcgwNnZK5yEpPjH0licwcpMW85KtcySw0wf65EiBvk1mwi
0PPM8gBlQKMWJ9+SIaLoCdzm1bPgLXqyJhXQm5INlgc7fqi+K57bF8buSTH0bbzE
zkJ9vS+n3Qbgz9Hfr9HdwReH5lXFxgI8l2gDMKdHMi8tbnCZpJBadmZds6mOshwO
u229L207ENHNulX5oKwH5x+2QTmPPVMWGhIflAongkEgMLVGwfBUSyTGIoAaLaV6
MgFDGjWdPUHAcUS+YFXBHFGtRYV/S0SL/lt3p2xPeHQZ2Mme9NVhMpCO8kH9K1ci
yEDmkuRJh5FBDoFbMUQh9nhEjQyEHd8F1ILTliogmYP3iXRvwY0p6xTdeQHgipSj
yPuckIE62Isq52d5KL3mefR6TQU26taayRCDGrQXkavmcERKj5YL7TS2DIv41VEI
8ZXdaPV/zPdGTxjzLqlatYVXTbpwWqmucPxuuwPxxyuHy0avv17sECxEYy1zr2xN
mUZBXGvY2JOWWMldo6OiqT8w3MdfoCmczTrxwbn/8gDqFUfEhJmckN7g2JEct2jS
tp9Cgit62FsrhB1lM4X653x7fCWaMk32bPskQkhUUkTPFGCIr52ApOczytdUm5Lb
PhTIzKdNJvvIz5aZ++Uopb3HI8qFIfxlehPdySHOmbmR9HImYlZ4PcTf6XkOKJv3
8lMtCJwLd7MMAXks9qEMfxGfsAPUAzPgPUurUzVZdHNDuKBHkCp7qxYr7ZFBi66v
MQwUG30EbYJXgzt7voSwyOADwIR/lLHBdGHf7Yaqk+sASVoeIe8YRcEXzyFMcdkt
TLzTcrmaYu5W+idcqC/S67Jv2s+8FfgIs3qr0OjIfONkMfKG0PrdWQMLyHU7OJL+
hAXA0DWOAW2ZKw8s3ua+vB21NJ3CbmwRgZ2krR/NSUyZiDNHXeW10lFxnW8vZ6i0
q9aMJv4lx5I+DNCfmxTIQSauePYEm0sIef7atq/zBgH8j15HJ3dBh6HUiZxGkh+6
XHVqrItiwyNgWyHl9v7Lgn771VSEF+CHmsiaS3Cnav2XvstYsDPdcYx3SbiCJDxB
gRnL6VJgAq/t30CrDHFFvXScq9uXmNHxxkccpMm9yxHSZHtcHt5pw1jxplAWBD81
HbLcpcPBMsa9WBbI3EN2RIOr0DNnXBO/jjI40h078NySknoqk64nblypjeu28Ble
Yj+kfkfanmsjvLiKAxXdZ0LvuTswHDZSFm8KX1BwvLJgrHV6s8VB7J0QLIkpQqyb
4wHkVe+zVDbDj45vKF5/nykDoQXHD/jtmUDWdW1Cfi6U5swwmusbp8udTaO+DVzP
AwW/iKpF9EanfC50Y38/HjLjJddWmAgKzZFGxjVNd4rr0cNuf1qqPg3IVHLgtT2I
mqfRC4fRFztgJXj7KYbCL9GDYU9stJ+XbJw5hcP7jbdT2kzrZmr//UVGA1fOf8Ua
dftBXSgNRI5IbZmRB+TNb4fzqXRbKtGG1NIKr/ZYjkbpem2VLhThsWKXbk/2V/Pv
lJ2XMcHRzUTf8+/ZI3ppmFmFdgRniPixZvJmOEk9fGSLH8otSmht3DRE1U6hUMbB
wr0ckklXDc7s4iQFyQ14tIpW92jzpfvYBEd2rMNhp6ekYt3zsYSTaFyEZ0u59cM/
WNIVJWNEg7Dvy4KKYFm+Ya3lLuXRE4B8mAMx8D3I1P+NFo0b4dBGbAswPgQE3kyZ
BPGA7KBNvntTXjyBzpfSjuuy9PMtRgzTxm9n8Sr4f6FKe8Iij/P6htKH3wIS504g
p3lIol0HQFEzUtZ4ov56vDTF2yZC3eH2ZASWyuYtUy03OyuPb/HAQmuMhVnXXTZx
GCOoEfjxLxwQHX1wKCL1mG0egaIs+nv/oSSH/4Q7gdBC4f6h+lCbdn+PS+0FGfM5
bw72L7F0vdGKQAF9dBphuHnOIQ5aQF086O3o0hrZ8yJ9A8anNPS+p/PYv7cO2W5z
0dquhSBcF+eHjDBLvpKu7br+eECCeYklkLaf/2gQO26G43Vfzjqd1VNUXBkM+R7E
Q0EFPueeXhUqUdzbCv0xLlTmb4BUwUJiF5fQqNlJ7YSdlwkoPbxQxV4S5GkWLtwk
nB8WuYM91tfcNZkRC+F4QTeNJ5P/1t5GegN6rRlDKeADFVayLCx1qokaHvg+eXa6
dfmu1w2EDj3KcgpO0N0Ry9+yVtLVxzKwv647mX4ItkYsIwmQS+dyJYz1lMQOhhRY
2pnDznK9f8mciC8ElVRmZuZsmtNRx4v595ZU9VZLKliDuIPcAT1apadYGpDTX0pC
E/KM0E6+8EFY7819cumuUVeoOv+GID07lYpJkM7BK54Wkwbh5mHrFfrA5jZsxKBY
xFGebFAqqVfijQvS8K67bC++XZfgm8FPiq28JF16SdjZzA10Bbvx4+Tw1zOyyR+3
Zq2FjaZOrlMlZfdomPWomIwu9Lhm8o3z2b2wdWGmOXJX7ZgvWRvhHkXDQPUk29/3
CQ7vgSsiS2bX50UHBdbu3dD6373f2XefIj6NvgNKCT1/r5s/1ylkMWts0KPyhM72
DykDPtvlRVfnUzxpZkQhWu6nr2GCm2CbjWwiVdVtu7FyNY+2rFY9jz9IHB4NasC6
MqsjT9dBA4kllBpJ0F5A87TQ8r4YiWw51vhR3Z5IB1xwLwxr/a04NNFHQxtFDjSx
HNgCVfkwnR85ABKycNvMiskT4ULIHtgUT2flaEkOImhzWI9IFhHtsLxYMA4yOjVg
mg1/hHJh0CFjcrGhLfwdMtTRfRGBwvDlxEZ8saswx1xfPMzQiZSCVOJpyNQzx6o1
kQn4dwUZWD4kbSCIKIoZGHauINAmr1pRqIIAyeLUPH5AXNx4kFyn7MXUi37ZRDdl
OQJ6mWCmYXT6JQtzoqi+74XEcw+9L50icwIGUJCIj9ecsx/U1a1Tskf7gYe7Z7AR
hKbJKq9GXiZ5fqaMMLGnJkjnhGi/PRHqNDfx7/YcwAhyNPckL/LGlWOFqRON11WM
0XNFwb31lCo1df2Ww5dohIUHE7xjbSRf1agnaBw8qs8/RrbZWkmUjxk4JuLKJtL/
/4FI/AHwZ/50EockAc+6sT5fAdg6Nvc53BP1VWXmxVojLqk+PGPsjfaDFxkXeRHS
LJt/TfWB69s890HWbqJ+NCs+M6B2KcWAlLrYRh4kAhtP1rbhEy72JdQpax/AgrDt
ym2pNzxkuM+9PZdqOA13vGlkhHEJ7NxqszaOrGlMTisxAwI5HE5ZFkpoO9s9tAzp
sPL92WjsIa+2vb5QhRuRdtPKrmlNE9Bd6UscfF3Fq1g6knUKZPt6yeDaEvDVGaTH
aPcVAlOrm75qWePSymT+fzbGjGpCjgOoyCt7H9p8zQe9x7J528K6tf6aW3RS3EJI
vw1ED7r9YS7nsvNq9Qy3UGSfRUjCEwzthu/N9kyWFuzS4w4GmFxul7ZHueNZS/8T
PL8NhpxiVfKs0uResy3alAuxwV89AIDUvEpWHwXg7XGQl3rwDJjvW98qpkN7aPlB
OHdctGw7vGNkEiFFPVsMQxKe8eIoEnbYma9pqQ0YTC7QCQJjcDzQMCDSi0ySJEso
MPwKC+rtioDZ7240qT5o9StbFHb9In3p8PfMToquL7naoCRGG3AeWrke0ePIMPuG
LE+qcBoccSZy5tfPmf1h5SBCbELWCgz+gMld2mX5A0SLSbNp1BFzMrR3jVhvWkkR
Hehhyl2Qj1PbAGraBs228dTbVuJfWHkx3/N6LqHNCi4eEB6/F1NDy1gjYdjizBHj
YFRde17z8l9z8cles/uN+D7f1pIt1gBTizMaHIxQPGKxWtGzPkymjVA7v2SV4FCu
kA6chAAWDIO7GvFgWYGNhy8dP44fobbSX1tMlzZknq3Wq9k4VRWFVRtgLp3wPyiC
7r5W6KqDMb+2GlRSg19k1fIH13n4HLNB/hVKDHotR0Gk7O0Nz4J2Ae1U9hvTDN/Y
Gfmkavb3jsD/o/zwPm20bLIs0CBdziOG6aZzGlrRFySdF5kUA87F0b1ZH8qZv5YT
mKrVGPvFevUe2ADi39PN7Bgkj34KC5gTaSGeLQ7+XUI22yEI5NxSxNGYHFyr4+NY
K798uK6J2oAErH0eP+oMMsp2j76oGTNkDxa82nx8myz/evNk7MBFxhs2T6mijXWO
/PJNUXg+8DrFTH5jIfK30JiycJchmNocwPCq4ZcP/0VlgkTjAX1FJrt1kJ2KbZmb
v+oK5Ab/aw0O2ohd9fD3AeNdE4pTKrwG6VHf/szmpqs0zJj+5EC/QYofjrlYAfFu
8e0hryDuYSVRo7+Kvga07VTRvFT3r7rJUyd9HNcM99B/8O6GWarwllIf33qD0blP
t+OudGCwUItNaLCR6Z+LMQS4hMxSH7o+gTKMPsQap0U4jeDG3FBoJLf2k/OKYnZY
QhSW+i/j8PGh7Yz9ng7S5OAXnFKCvMfB5WVz478aNq3i3Ozr+ruk+KeBPzM4aVgB
cTyABgRTO3NcDCSLu/33AvkydwxhrvM5LNKBr8o6Z+Zm2r+N4gudiyJck8ucZN1b
M8xNO59AquWXXz6OWWww+toTIyrWvLN7DP200XK5MYilAEJYnPusGJYoFQHD5Ow1
tLUJYREjF2EP126npxDZxkTtLVYUxFvAxvxLqnuvuBOSmuIj+/KWYLozKqxj0Um9
t0mplUzHTonf09c+X2Z29b4A6UxQA2Cuh+vXlDxcXNx0mI3LlKbcxkLI6Fs15xvJ
wSFfMo6z67HroDpSoiGKdXImxrRLfbVLNstfa3PSpJjxivNULyqgUaK89/6EeySo
HYP6tMaedaQIn5RW2tD0LZPVY9uPahdFcnvRCxjTkZpdiLPfVHxWiq8tvblwjXj9
ID2blhBrxE6eX19qsAaA/DZoYfhUbZp7JMrDRsy01iH9GAoMctAmWjjP2IcxSk4P
18GchpayEkVOqMCqCBZZwNmqxspvfI6YkZ+E46v3E1LB8K4Mp2YbevPYpIN3oeWD
7SquRgTNCvuVLCdtuqCA69ChB8A4+dX4PTcMxNRRXg465IXhh2Iqq3bptkKZ03aB
RgPFW2yoDRcIh3JzOPyWV9sZwIsB/glSzRKFmXdQt64kslZAaa+0P0F2+cqaHTIH
b7jppMYT2/abI1HkaSdjvQG3/ABL18vXyWrpK6qjMHcSSSlRiAGKIZmMAgxL7cPg
KYYOJFaAPr12vc+2CWokD2IsWoSysPhVWIwsjNM+H4f14oL2nvaNG5JALh2Wmc2d
iMxECJd/tEosCV5uBc3ThWfQVtah5z91U8H60gaQh2XmxVl4bnHCoJT2the59JaP
jXAVRxoAp88+ozzNEfkHFjDkihsLXt63NwMON0/YkD2HTCdKOBVlQ6eugQ8oC59w
YQi0/2lXYRENYv8a+a+vyuRJpUFDvVSg2DVv40xcrkBRI6Lh6usImuL0UYfcvDMJ
HH2msrNmhHoqVlUgwx0oQYZsh8jesPKV6taYMBLO4uFCMCGTHv6rlcmnqZzf5L3d
cSd5FZ5GAtIWmWwGQfnv0o+m2q8KYNUk+3IEQsRL5hadYBAJJacLZH8kNfyDfZMv
qyWmPd8MMPQt1ePQfCi37ceHs7qm3P4sfj7+X3rg78RZaiJF/LxljrH6wT1Z6pYh
jOjeu9qTBCbRYqIr6jwU4KK36fab1F5p87VFhFhk77MEBQQiliduLWP0IiULgZ15
v74Tt/qEZLH9YgqUxF4RtZeQNZWATyGLi84T+hAUlvLSVAA0wW3TtVlpVN4VyBq6
eUThTAyMG6RgloaLI2JxLnN7PtF9J3WAgAKJ53WQjuMEPwsYjJIoUi+Q+AJJu7sj
tXM0yqNSCJWgS+/7tQLW8kU5txnabXT8kOBXfMhqz/j+EBk/79kT6EJXGFErcVFs
iA5yJ53wAi9rnMMzWSuqfIHl0tQ2hGDkz9xD9wMwlqslybIkiVcNNojS5NkYd+Tq
50tjiOV3hYERUwk/nymnJoDKGQ05DAy5H7Aq7cVn2ww8s5Plg565xgn/v1FWXJ/+
tSxp4UsS+bjS1VYm3e/Y/3nIzrQM3ot6AI5zzcapXDpcP+PUCQ0DLpWrlWcXdyQE
xUVwXahTrFDb2Pk/HmqeR16Z2xP2l0Vx/wzcG7dhtVyLoXUNOMX12O2v4O1Fxwo6
gEs5AGdg/jcbPM+RxW2mX8P1c5nDJD4notCtTiT5Jpq/YkOl4s41kOM9mAqM0r1v
f/qGobgip2C1tBMl/gakkAVLgL92IM3h8UkloT+GbWsSij6S/XZCrOlmeEzFG72f
KLmRiFM0P/SsWnKeex+D6naJ051RSsW6S5qkUqLqoOYuCfnaYp/qY6fuervAEh7t
tfWRSuQbjOaVbgourb2K36L4MpGzRbHANP1WaZ0ByPPiAvVHVwCEZwwcuEP6QXKf
SvYIoNMBqyTyHB5bamWySL2e845CoIRElF3JvAKSyK/smYXTo06jL/piV0VPcOh+
dxR/y6hYTNOhWxAoMN+Wn/nbqcD1UCagOrC9AYmEG6RHMaQn3GTJuFb2LwVBCezJ
j+naqIbSEBgMXS/jvFUhVaQ+7jKwy4CcoaVggIcW2yvlgCpyGrWywWKbCihGwQ3O
7kEh4ytdMVHqiIuDn3xwD6RUHwfS61xzLqofckUMKDmX0HaM36hYyds3E33tg+Vv
GaTkGj7gMTH6w8pCf5WXOhZrXJRvlU5qd+xpu61Fc671cZ4JeO+Tx3HkJ57MnP+G
kAUyxJioiwOQOOIaUnEuW1nDi2CEkGtHVJAJdXqZekhhLSO4V6NqMAwZP2XhywW9
1MezugC9mMUotTQfM+39GKEtbxbcDoyITGO9azwwNTYtdLGTZ6UV9djqa006NOVt
NG4df7oElD15XTIjrsx0+T6UcPpJWzS0VxDZyo+4NPGJW5Ve8kbmq90ghSDCNQ7G
y4DMvHhE8TZopD5/Nr1l9ret4lJ1Y/jbdIidSLHnoQkfIy+DRdCm5bBRtk6E/W/0
y7yQ2utY46KIToubKIMkUz2ph0UD1C9/txf5EyBcd7xO4/VkuJszm8n+fBTwOpOm
nbDS0HXk5JQ2kv7iIv7tNMBmTox4fVMg3g6UnrKFmzRKO8bsYQxLQ9uHj5gdNM3F
KuMcNnAJPVUt2jB6p8YNslBZnUpyZ9VxMsSgEuhGYKy9TwbllhvMOaQ6hNGjWiLl
jF+gx7oRehASYrLaYHJxPLvitt1X+/NXWUGXe9PaPR1Mk42XSKNd/qWvEL74Nbd3
nJlKMpUGQydSjcZVnCStULVoD5qAaim5fn4Ng14rVW4oZnqMovx5q3OKpX/7EqJu
ZiMFHi8mfCoeUMaderBDRZbUGDMi57mdYen7chbuAWr5YW1+qoATJauOcfE07P6b
CdxXMnm+RRpuKoE57ZqymtH/QZXjpLJvPSyTKQywa34ImkgS58zoU92m0ABDVl41
1oDv468jG0XyrWkeyELWt1uyT+7qhbrjjV7n05lye1L2rJV6/u+T9pCKMtjeTL5X
poGAKY4IOPtLNXuwA00QpGAFiPxkwZX2UK4XHPhHHCoZWoVJI8PJ8h9uZg+OEpCt
cv22j4w8iVZlDuHIvaU/93/TlT+Q4/0R3pv3mw/PM12wQ4H2UX1QVeHyacCINdbd
mEVUYU4Lx3m5IeSPM8D3iAfXMrLAAGP/a3T6ArLAV94S7O6RnHRZXKz7jfxdOXHY
BGOmsnD9WqqPW49utDzAEe/Cf/pwhNCj+tJnqFOpOEdMtATqIkocH4QZReFfnRG9
gGENze9a/MSdPfnQ3UIJladE1OfgZ9zRIJBOtfelZTdP3LjkUmsqP/446McdHaRF
q7ZWIbBHQMuP8kUV/Q7JAwM6HJP0OYHX+ynhsnx/ZWgXZrXAx6w681PBJYtkDfFL
s2vjy6oQV2z+eb5drYNT2kQAB05qHe6jOnGYQPSMierPlUSY9bICE/ngZRUvsRGh
hTpuXo2OBDX+X7OR+DTqlWNgNv9XPC5zL0ItrbVla5NssbOJIlXoZXSILjLYn/qh
Ar4Da8n3j+ykp2D+ncGKX2D76tIaiJAP2w6O6Bh7s8C2tjyKsAsjNUH8XqizYpc4
Tc5JwQEfxxh9GFA0DqjdvRxWE2HClpMaFmO4eOwM3hhor53SeLuNssPaPqB1VX8W
/uk3thk7jNRUQLKZmdXJXQxdhzpTzA4sbgFwGW4bDbkYzvoSHw4YPJM94jcuhK/h
OIsDLGtx64T4wfchACTRE8IGtokTG0hQ1DoqsyFh1Q/Dn9+Ng45Eq3Z+ZR99Ygyw
5fCDvfhp5H2Z6x3rNxe/FT5/k7UhCYTcolfyax6BFMak4eKnqFtf1JhSQH/buWOr
tzGse+cNGLybbwvkye4btKsZDoVTMZRl6lcsFe5k86DeN92NBcJvMMfNtbk4e2cJ
b5YBsywApl9IU9ubCs5XWux9ZpV/n3GWhwfeaykdpVk6Nu68zluGHnbHbHG6kfwW
85i1LYs1JxOM7mv1AMIC13nQ1C7my4ycDiFHe2EVGIc/NZZhhtuoMXSBVyVljaa4
nZZFlGMALd/R/R2qaA1P7+5uEPKc2QyXHJn+OCob+ye/e5E5sVSHb9mhOthn27KX
EYJi8SCZp+u/KB9EAcUfZ5jXvLYS+Xgzi9x4fX7SaUvbbsGA1qgVd9b+AuNYlABy
I8OUI02JMBdmwT4yIHZuoejzSjlcKyj8/zGs1iU8sAbJWusw751AmTnbcxC9AhsI
h37hHs3Rrqel6ihG8RDHP6SufmtGQ+9TgCun3RLwc6ZThWl9g9OoKJeZxImNfRXR
XaxcV4232X5KykbSsCi8T1JgiiQbDfl3e0q/3Xomi6zJK14xTDdyPESgoHHCDBPS
mnSDGbSKXR0so3WRxKF/ZHoUa7mw728mc+RWZsO53btGNo8SPkt6FFW+avLSgHa4
+ybCz+Kn5JpttPbew0iPEiuyMmjaeuvhaF/VDk8zCE5N1g2xg+YY5tXMC18Vgta/
ytrVl9/5AtElZHAhOSXMyuMpxkuMZLFrxcDoSmFlhQanppViSQQ/GVmIcZmOb3VL
mu2dNDBieL2npxPToPqXtKUqfJiYOYn+xS+rvQCSFVNQvtvV4k46FYalUnys38/c
gWc5BO8lNXHyy7zHfy/2Qto48/zxq6AIBcbDe/U2t1Z5bCgbw4B8FxXMc5hq9r0N
0rqzo8s7g1OoAAP2VNh7JQP5NC0j4TmnZMzHFGdGvdzC9PFTqQAg0jNbHo2YGN1t
r6smgOPwPCiO+9zk9QB2udnJqO4HpPS/iJrJIQBEN/JuLcIjsNFquM9WaWmm/WPy
4Z/27WZ27S6U4H8qxbXF7b8ZxJDzyNmpWW21h0YrbOHqVpsyGh7x235tZD2bNN8M
pPfy8VS/ESxidqzl3xcv1Jk9QIb7fvfMzhx7mWgA+XWxy5qH0/sc/kWIcova7eLn
YHza7/88wKW3kOkp2fsqW0cMLPGILvdsI5obCk+3omREtWeFt53o+NXG1B825kY2
GwgVKSFfbXC2lmPPi7paqjEAUfyjFqS7ySBEKCm/1E4c5rMxK/nhh3pr+UOY6PUf
rrRTllAOM/IYUNN89dIGXaAmrcBcBK42oA9hn1kP/DsHMgjg6zSSRFX7+YeR3pCw
uzB/z3Mc18NTlWeRNXdjGeRievei3Mqfgq2OckD09xbguvY5Fl84PvBp2zi3gsQp
RDAp6C5IQfcga2UduMKINpm7e9DNIR+DoVUxVY4Ll5RZxkVwWhbcqf5DLssdrJIP
r5yZAtwoBwmGaj0cSWqlYkDXZkTAzfcDbBuQ0vCco/WaKkI9GamI1NYUM1PAni46
uw9bRwUBAOhpuYcoVOSxWPYo8zFtGltjf9WQuIZzO0eOgPQcd8e5AAK2P/7RD15I
TgufkFDWDmHsIf+HUwfIF7jEXFhA32NqztnM2vM4Tsmt7cyRR2uV4VrHIZ65oBAz
nzBXgpp8do+xStw7PMG8si+jEKd/JhAFd82Ac6FEchIj71pBnqWQTTXJ6ILzqaak
M25Bho97Lhiq/rcJQnpy1DhQEyrbujl47NsVn1y2MBnAqpRfwXu+hVBstIm/zLTZ
k14OshdYSZW71bmMiyz8GLkGX7Hc2T6rBKARhBwy0bhrtr2pz+yPPfkk5Jlekao5
JW/H+lKs7sj8bduP7ovx45CjO4qhyZnloDXtTND+TUXmA74zTWQnhp2GpGWcOhap
5pGIDsRzmUlsuVdWblM7GKooJJ2dU+jUtpwqP/zcMA+jOjr7xowxwIcGnjsp8wr4
zs64f9akk+Ovq11Al4SsEPpWtaqnW8U42qA2EfmZy7ATXgZ6Kw3Yfx2i1XpQ/L7s
/FO2Ejvk6kTUrhqqB4oVfCc+RkBF47gi6yHdq0DiVXGeAO7xvmMjzeaSYQh4HRhq
cQcVmFcIXBctF1aPwLwHw+3Rs7OVVVwqOZYtG73DwwzuC269E7i1U5t6I01mWMU8
ViAmWcF6x2+JsR5OcQP+WCCrmQR71AIS27RT7M4Bfpw31mGwPLBQnCnXL5QwR/pW
3Wg0wmgTzJSAQAgyutZykRaAReUs/qt/0mXmLEYLEJeQEe6kqA+iMFMkV5lhX07p
7xs31npp9diAOuo7T7DdS6K7NKfo2pBRS+xyFI0FENPL4xXYNEijLtjr9Coj1LF0
H+Sc8a+3qIW0e4kqfXkrby7VJi1wgd0557CoVtmxJdz9aXab9h1oxhGqs7/8H5Xx
XaIDQyZcV3PmF6WYvFSL8yN/9Yt5U72o7rgF3hfEV0DZXQdWX8N8LfB9WUaQfHN/
wUalU/EG0SisjnEI9C+mpZO3Vvm3jSuw8mHleeb6oVSZS2PIe3w8Qb8LvW1GAsKu
sLytPzE5APt5KHVmPlyv35WV0qEG/RbMscwPTqRCDmU5uiQA+NKXLw5/ZkIDolrw
kj9NwTV2rjrlXgc5eyp2hy9JEoCG0aU1nrLw3mSXy/2Diud09iroESAzKgSSfnBA
13DNFp8lp6R92jToLbqNUhTslpshoHg+Y352z/ESuSO8GH6fT39+WLp7th8m7MDs
sD6TnPVHmu7nnpGM9miJ6TvQ5hMLBDqcAGOY9DFep2s+Ci7EUDG1n+0Sd4+v7SxW
Yw7UHXlkteQO3xOiAlyePeyl8CnNfDthXrs7wxoJNLPM+S5J2ka/nEYelQ2mN7Lc
lVnXrHSOaKhe14r6gQx807QbrjWoc4ktv6AjWfigJR2D1y3l6LFUw6wwRzqYNzQ0
gQbbN7D514aUnSAwm+HhKbekMOrxOKwAC3UyNEZim3awlzCOH06eOtpUjs5UT3ft
FxKPMuu9PWDChSw+6guOIdOs4gKodBtcEIdUbxPV+vaNHYDfPb3QQOJG5ygFU8fT
GjmPPqTOY6Xmnmt1+Qa6A5dpD81nXxWd0Gg8s2W+wJ8PY1ACI+PHTfkgIqwbywLN
T/vQx86h3zB/8kcFqhkXYIg1vpiwi7GSSOKMtmC0eMdBtAN990CJrdmQxr5uxDER
lukmlMMjSWJUYylmShHoTMeF3SoIvY5XHtLsC3EJ3sUs0Y3DcLMYMqxX8mPxu6af
deEO9YrfDeAoROLu/z+yLVGOUn7LWSshaRWV/KQOp8ys0NoldPzzhFOWOZAapPft
P2CRtHC5OOfpdO6h+ZTnSoqgEhrHjpa/XUsJPpAG3bvAqmx/wA5B0M1QtkGLJFFh
yHvBv/LQIfnhbCN5ecrtkYwr2dnvA0dDQ1FnUJS6qdIY3+OyWeiM7LV1zddPgBcY
XpYSNPZ4FB39Et0zhEWc5VjD6LZc8vnLNJo/l6IviJqVUF85+w33Ug+UDPmLA8Hf
QNOOEXHX4in2Hq2uwPjVGF0iImzhTIyy1OMj3+/2A4MO3Eq1o9l2y/nONs51iRqI
GKt611KoUMp2i52elqxUq1FAmoiCvcvDuRifUfeRkNXPAig1iMQTVyIAN94eC9eR
wIYxX0GgEHLfWyKHQK+QDKV7BQwWv7aPpDahLX0n6Z8vVNnUdlH0ikB6ALPVitWJ
7v5LEr9pwP404utWtrTBEeWRdJpAsRAl6qe52z+l6ArzUqAWt7rjFDaF96f1Sr5e
s1KXR1q8Xq8LV+YAlDFcp3YxqHYG/gsiDGZs5ED0MmdUtyQqz5JSRDJekSyZSLmW
z6lbhIypub70Hgi+Qr/cuQC1pMIt6sB1QhhnPbOe5NvTuvy3vArrwoN1HRlc9fNd
+pnFYk13TDy/I3Rr+BtU2tR83078uwMOawk+Fas88jKBTWFdxyq4JtlaMZIaPZ2H
z+Ie6GrrBZGHlu+KwzBEfkzZKcef6QydBjWKI46eNTXUlxT8/tseOqaxOOQSceXS
T0Re4HGBCe9nhcLnWySl5ILGyik6Vc5nleLeaT0Re8hMWQDRUu1AXRDBCtMSKDOH
umfoisAKzAEZOKQ4kxkWV1XQec8+M+gX5L2zioc8G0Z6eiclm4BOku6a3yPZD3hL
CEACkIAicZjgFHxEW59YjkHY6zFHWXxMYc5znCeqp9knHU94lXDrrKMk4PTK2Ynm
B5r8rgslQiy1isdJzG6soz8k8tqoCl75rgYw2t5EwWpG0R/IPUKQ6TOkXKguh1rl
u8XikUGxpe8Kntmu859DyBysrSaX7IPdW36zcWyJjSwM+C8Yy/4Xsq65VwIVxFo+
x8iMnj3tj7gTAAG+56p/pSvOtA8TEKsCxv1gsBVTGPTQC+u5k03R1NxfUaWg7xC8
KoZiqO22bOKWk0s7Ghc9AwGFAfHAR9dTaB/xaft2v2HBBL/wY0oxFfZ2FtQmZaPC
IdssriOiO6eeqjSnfTFL0/3Nz8NQ5AuYO8yhib5CAROkr0m86uM/fN45yjqfsMN+
xJAN7ZqPvO/SUH9sZTu4Cwy9PgfRSKiJ938Qh0m5fcXdoK8Ib1nGe1JEiJirqmwX
GVavCtxyr0gMsruYtNTLpm6tX7MydaJR/YDZo8gF4THC0ZenVyjygLqJx2mZzNzj
i1ZuE2cMXaAmmqD/iLNZ1xyBppc5wOi+YhQeB+pbx6vretn1ezB6kUmvNPsNIa+s
yzmQfH+eO4bmPtnOQ34hrwBirrsOstOu/vk1RVVxw21KHVoNWGKfDalY6B+HgUdY
WY7GaRfb9WUu1JTYOtk6qfXZO9QbU/fmFHcZWi9wvuCngMspDwM7HSuNZ59XDw25
qnnbLfMLbULrBtBAwCB84Yn2vIVAcm3xy7p4d4dk6Gzz6I7YPymCLkmcxSFbl3hf
DNWOw/8PL98xtpbAL/PFX4gjc1k5j5V1Yu4MfZ1f24XTxUOqTCR6Sb/nu56LEeea
dOaPHdACsEgmnqBfbq517Op+2855obqRh3SNpIHERrrOTZzex3U0m+LRaHNrfYOl
ErKQQmJ/0mXawKYAUtHn7DKmYTdxorm3DixHTbmwqS850VV3yuPjTzFYplyCwSXy
bZryTgUckBr7hNhX77i6uaPYVpf3r5TpgSZOfn6AKzl3oqELD5l+I7QOhvaWTjLC
QEK6TneD9W0sf0DGljEaSTE52+0/USZHsfIGtbScm4aF1SCIpCS0EOIGk8YLfNFp
kysoZtKJLJCORsPoMgJrmnNkEOoy535+DK46Eq9qatSJ0brjpAHbzWZN681glk+Z
Jc8v2Tz/X0OwAl0bBayRpkZZ3ZwnVnYLLdEj//XzK9cA4f2zaWI92KVY9eZbQteh
HxutZLMVDOPTidiKsLqQuVLebA6l6aep0uRrQKpd83IPYlwr/OSrwgLIC5fDDaFy
HowpT4Zv+6X5sTpcLX32v71EzkdZ5Q81G/lEp6yStcvseTQa9KVuQdm+WAJAPi9E
iXALlgqHxno+1FRst7bJUXl6GEMWxu3ZivdACJt8Y2NBuCYL+xU/ta8MGpQoe9QX
1zDtypLDkWmLnXtMqHqwD3Gi9JDvT7crXPg5jKGKQhx3xFVHlCBDPWJiL9lEITaV
QUH+GuFbvYVHWtEs6Nfdtfjfocsm4GHp2A7Eb4ByVhQ9z9nZDpNoR2uCqLagL0As
p3oK+bO7c6mTxfYJkiwMTbwUD8qDX2AjArPyOQy/xnZG7itNk8Rl8FAp0SFDG4Yr
PqlYOIu8RrlDpK46pn/10F/kZS1AeA+FkQVZ3wwj+pYe/CTB8v8u8AKLCHTY9KIZ
vPguAyvmY1Z6xEstoAunR9hRF6+/sfxnQOigNlPiL91ppDCuTXoedPKmupxavx17
VKkWMKKDbZ5s09C5rABtqOrQKyQWyjNHzArd8wn7VwTkSwVH/4nrIDa+a5w6L+JO
dxLsQDh9pjVL2bEH26jURiSO0Fn3oQOyOdCiJIOIdYmeB4FiZQ+C92ojwy95CTv4
rn6Ha53olI/n35q+gZmX7i7PM7/qJWrMgSFEQthYOVcWdRe8XXuL1s5udyFWXr+E
jRWSVmZdDkSv34aW0+2J4ZJjXZ6CCYQzBIDKxtt57Q3wxJbp8E6/7EFxni5NOQPm
ILXKCqO3YMHJJOY6OF5BAPvnhm7m+KvkoTFescHLj18d6etTN5tQ9Ckw+qqL5hes
Or26kmDRnFaaFEJE7EhhJYpF7LJxaVebZE+CFDSpfxf6/lwRs+mABegmF2qe3TiG
KuSDGjnhzrmJeBfRcXmSxBaxMlH9jVMdhghpvc9gJKaOD4NEU7cZXUQoAm3/FjPn
DzRZkDZlepfOffX2mOud8Ez2/jKWAa+wnkBmzFGmdYumI3BscgVvRVMUpinPuGUV
VThBEXRrEZxREJH9NOB1K5yXuHyO8l+gz3MYoXa8wVKDhSGzE3rk7tWJdXfyZqkN
MIpiBU2RDRkFa2WNNwQGoz86ZwwIdXhJxTlZfD7hWbUO/jA6x8HPCBimT8vZLN8M
iZ15vokckeffcRVaoX2IA8y0pTqO2/wcHZoVu/fIM312SmJtvzM9S1DD0mpMJZfJ
7UmFvVkImJjH+pe0/NPh0gLU6rYZyhHR0nCQgtVhwahtggZb3NxSfjMkw0kb6GT3
hheWixMlnCdtNM+HC54DTWnOXuHeit0HCYkC1Hb4cXM9oYm/RRfIm9f8psHBXL31
4n4dlkxA+G+e8oolrkYfwDRz6im/VlEORn6fmJ5qttz4gfMgjfs3UjC0pSphflCq
feEobIrOGqCL8+Qt/FuTI/DzYvNHw+xVjR9MlrgAnj9vTyuEmRklEmop8IffzzqF
m3Ka06VBVSk+CzY2iPi5udmRv+Kus2fAyBqDCLuMbOiZxG1OsvIdNkoZEax08Ucy
ftdtaI1Hqls+A9WTh5ZheW6TTnLv4gdtT0i1SBDow44CkHSaDExnDAi0mePiBUSm
yjCwCIn/3i/mnZ9WuenrQ1hw+C1m5FsL6VAdJwvOJZsfxgS/g2Y6NapuYSGOHt8j
QyDi8TDgwsv36sGtNlqw2Fo3SfmGF6n9zm00lYaQkY61vE3xCqjJgqhqgOn7uH4V
VIsQqXYnCeknbMNEnCbzZD1lX+hcjvhdS5UGF8WF6E59ICEWrGeimdAHan6SvLrE
nDxaJld6OyIvrrXiLsL6WlZd71sIfNUV06aN2JWhX2aibWWNu8Nx4WvlbhIF9oGs
GzcBjYx07TwqPo5tAqh0OWuuBFsvHyGshTvvtBRPnnuOOHBgqwkFZdKaR8DdJQyx
eQGwzA4VpZcP1mQAyQTXqbUwaWiJf82LHCk3zihKkU3e9YT0uYJyt9vuExtndxyG
lSaS7NiMPBPPkB4GFeRlXEhXkA1U8tVxDbuIGkkw3bnNvbgXYiPMOeRjviXtLCyG
NtLicpquHs9pKNxJPSmXr7Z/f7aHIX/LAZEUSYLPd4BzJw4lsvnM87kTZyIitEjh
0F+YCLd3lwZqWlZXOOdj4Ben5qKVpjOCYb2EyIkuGLbwpF8+94kR2Ihbz0mFNJr/
xel4/i0ulHG2grrlG/DNe58GgmfftIgPmkLSPMObpCXRsmqP3WBwAY6ZbrvN+H0/
qTzlPkY4G2JIxxz9rmbiD1tdHxcuqUd0o9V6X5jYHjeEzznVZaJMAQ6BoTbFa6EI
9wRhWFKGK2vPbs7JHJDyhS0XruKYohcNZhFiXOSgssCO0/rQvPEYHaYcFwlTucVt
OoKJNvmfSEXqFIxt4xYA5/vMapzuXjmL1rHvL7UGxu8xnxmmDyjGyMG2KuVCrqGk
gXPNCq+pgR0fFO+7vszHW05trBZDcLzv6gs2jIEARRJ7DvyWIhXcqBUF0jiX63Iv
NHqO9ZlTRP0VZzQPlwqK3MkQzcfF1b2DBEeF8mW0bawR+V94A4t8K3eqQ9AgKyKX
btsUh53yzqo/zxkRWvD81nZD8+GkSXqkWxH6LVUvRHciL7h4yZS1tyZlRXTLcgbL
1NwMsCPkkqzGz/zl55hWWD7BmmHJi/oMw2sLL3EZgO8sbVa548e2IprcsoTJBQMK
kAKGWXAKbYdmnH1UstwtIcasFq7JB8CM/QpKm1bfUVYTNUZLgtG75ePU9JbE2O33
1KhDNZ56Cox92JdMVzdsZ88whaOt25gPNwGZaATlQmS+3ZM2tZfYFCGYTc1XwVNe
Cf+RiTRCmPvqv8r32RzqERDDyOUuXxpCZHcC+lodtwUNCNBTreedFBALlmDDJjbt
37BZg1jW5lUFAgeXJJGwH51Sye62DpX4P7AAGK5K6PY1Ombf4eIl7EPCz0sg0LxJ
5hPc08PQBGicU+DzK3WGH//K9iabgf0Gi7P5eZQfEpfl8nabT+hkOY6icps3e18R
mWEE72Tbm9f+uzp0kDtUSYYDZxEZBRHhwcrWSm8OdEGoDMf/mfGi02g4dOaDlVPw
IG0uoLLUJtTxB+CJg50i9i4yiCS/d9GyTE2/2Oj0XLWR1evqY09iYKKXi3oxglS/
vm1OzKCJsGH72yKSGlPF7v0sJEakUJrIyo+S4tDkMoVDVVjkjCMXjeGUAxdadPZ/
rD/Q+qAkPW/HPYlC5iLr+vzMKNbOdsI6Mr8xMiDm6W3zXSs95E6XbGGqjuL16kB4
iOZSVi26zdqI1z5TRwrU55Frcf/osnlOPS9do7ROVQ6ZWXOMeY4mboRjw0ueaf8H
xKdlGSkBniWsOSC4odJzaQxIzNans11ssvNHS7lhaVXPPpHsoqv4TZrLeihi5oEf
mKCZgEc3XTkIzNRTBxgZs1snlU82gV6EAdtyuLQSylN4W6yQJhbaJYscQjIYo/0y
7wFI5gbBu2M0G2qIIxhfXIVqDgc9fQ90X2pCews0ozmDeEGG3MfgUrS8G5/sDzo6
u04UsrRiebUGXdP+N42LFwzs1MLNrUUSNVglYzKbjPApCJtEaMVEOLUeF0ImPjMa
EhufNqueHUVhxhsUu000MKo+4pGlGG3uZe9M9l43d0OqumOThZjNXOKug2T4mtEW
o+klYKt3kZPBCutvOvY/u20WDZzTIHp3C8D66vuUU4tM5jfZzZogXF8+BwnGpQYe
JJX9YQEKKB/DZdI/Ka9fnSP4BSU2MzX3fQJYtbI8/OdPKW84ntsunfrMdB0yTCNf
8Vl0Egzu2h4C9To05LxNbJeqRyICCE4hu7Z64Qc4czsTAthq5g7JdvijSYjcg4NZ
Sz/XI7j3zI6aHCrFmqaMg9mQG4HDi3szndK/Tvo8g8auBXhGa9fWBf5JlhvfxtVQ
qaO0HsM5FyGKJzNI+tHW9/z5WkLjOXMA8xbM67HLq38bnHnYXaZ1qNLIFWhzkwKK
FxwkBE9ZwemPqPazXet5hzPgYJAbr/1WnNNg2ShtiF1qeGFPj+X4t1S5jbJncYdF
tNXM6t/2Hp+TckkRYTMFRTqtlDkFeAT4dJK8MiWRrFWxreYYrPxBEN4SYmEE3og0
DlHI7VLZBDxaWFqN1oKh/j71hBrby7pOHC7pSkruuu+WN/uV6HiQu9y9TxW3goPh
98zaMWQlV/H1FL3Tf/RF9e5ntvfH3MH3QgXoOwptXisnTp/3k7z/Z8MudHZC02Rg
vsQ9u1MW+ZF4OTGGlbuE4KTVeRXV5TuMNwVV7Noud3hYvl/tQGTaWJMR8LeiNMSA
PSuMHEzrDikWmPmkuH066VvIstpXF5vM8blgTd/NQXl2TiX9WpgipMXAisPj5Ah/
rhTnpCE4BqgMqRWOPrGDs+QCyVkKMdFYbUU+CtLrxUyx1cDVE2tD3NoyBSauxU+C
n6MSlYOMFJZbZyEoECQox+3kx/l6CZzFHiseWmNO533RNjxds3/ftclbQS7sq3nQ
bvbTO8djb0HQ2PlqEaQcsV7Ldcm2B3DTff0X+Icm0KlvNUMVwp+2yQEvhYYSXieT
20UFCNnmwwQBcWs6CKFhTHc3cQejNc3i42HPBOLpb52DxYbPXWMWSVRLVLC7/A2j
w+nngC3lELqFcCSKbwsr4zeMr2iYuqcfbPWkpdypW8SbLsIffc1gPugf5YQr6hsw
tKuktlUyI80fnhBh52pJzOAFtYOiIBxsdXA365w9RTbOWTfVPnuDcJwIorQjUugL
DaHu1T2YD0cetI1tT81kkMOLP5A8f/Mg50yDjmTmn3FqBoMdCI+nFN+kWDzY5/Ym
yWHUyK5TqZkvaYvFtquVsBM8O6FhuVH8i6BDMhRAIry/UzACwcdPqlcnawXGWFXn
zVmh3UD74lvnqqmPcJ+ylMU/cRN/qr6Tdj1QG2LW7aVNlI38XHMu0tyicNKzVA7I
ko2Y0ZQnwlrIrrjew5F8/uj3IC/g3fAurrVVpmn9Exz3ioiyZaaF4zAaWMWyY0gk
BtB/zJj5nSi5eH4A9eDKFKIO12TUctnEOk2tMctElWpg5TgtmZ1gOraKklp5aE/g
R0SsorvaZYG4CCifAq4n/zqk2StNCnlmQcAz9Jek+jwvf9Bm1+2w1Qca6KlO0pns
tCbNfi3UxvePXTQl1ok7ijLpnWFRmIDUHSTEGcmIO2TjkuIjcjJ+AN1FhTK3CCQ5
gXS8GGMTISySv60XMX/WXj7boBV+Un6YjjG+ZfZvzdeYxT1jIDlGewZIq5jAHlOP
ls00yKT5ibQdwnt1gtFGQBh/+Yj8UUOclinKhoYbl0GOm+Ue9E1laqSi+hMqI6a4
SOX20zh8Ngwzpq1xE+/RaOoHZ5NCvLbDuOMsWIypelFO4DdplYyJfiX+xg6EcjTg
v9W0vnGnfUurvro4oGysSoj37Ycvr/svlTTU8o6K6VJWzculZuQtH3Z/aiVFjKw/
OAbwlpg3xqoT9Xiu9QNOobxEvXGBlm5Wa4E/H12lYewIHt0He1eQmcOdzFPJjI7B
HdXFvosgZ74CP1rGwFdO/TFxDZXK5KL3vEmeUq80G0orNDHi+awOuPK2rWwQshpE
dlDhooPG0dTaJgylbrwc+p4adnq8ZX4+p+Tgajh4XPS3bLllQ3bPZ0mCJp6smXrL
EzC5qJ/Y9P9zsXQsBD5dmVl/hDmq71aqYx/RZTuHv2qAFfqPbNnI+HLU72eJpXNF
dSE3BYuYTMve+pZFp8hLd1g+SBgcOrnrDEyWJYcmIK5cIpfuEpkMPGtaSL5C0wUX
RhaYI5likgKt1KXBQ88v2NT5HWaDHde0CDzb3pzmngZWhrxmVxFzTg5KswXkno1p
A/uhIpFGOEdVXIEjWZ3YC/6jxehZdWCVEt2eRU2cJirIueOJDVGfGJjRuCSZNhwU
DBZ/JPAj3T4BeDmA3/LcpNPQQWP7A44thdTS+dtmWwEfRmGw90MgClN3fzGfo1Ls
F2OG1ssAdlEt4nRxGnzwZfHXw0kCnNAmpMGENuOhGmgEonYNxKU9D5AOtWTG62mi
dIbF1QUp3Kpb43vbiI818Fn+yfZ9dTpu0O0VCPmYXH2Hg1KXp9ZnWaW8GKJHOljO
2G7myW9/ut7t58K+nwBdu6v8nuCx49jbmeQtpNV5mJyUWW7Ti4ax4PQcpnnteH3/
WLqGbUYB6N8ekaoBy6sEUBflFfTGpBqN4j779If6nJs35hWKyTax2PE0ueRdKAvr
FRFx4YINDlwed1IQPQ6BJzhArv84CZ/xkEUBEy0cBHkqPUzBrDdJUnHaJUEtsSDx
pLY6r2DKM6iHIau+uWd/GjgvQxZg1dQJg9Cn3O8R+gNoCcS4rLIW3/2uRO98psF/
sZ2wFVoT17EGEG1I2Z8AmZdbgLXeDMF364br9Br4OeKwiB7n4gRIR0VQjHdSIHJa
WbeVvdQybgxl2fxwxJyu9SXskP/CHJtG5s63wVJl5mHMLAD2TUGsFuF7hfIxtc7v
tVIu4LP6eI8zKR8Ceqg6IpYJfSCm9/QBeXAvDxiWBWD4tLJbqGmpQcc8/z7bOmnt
MFGhbzix50LkQD6j0hxMyu5CAKWes8CC0W44a7+GxsPa81v5SmMkELLVD4unXT0Y
KAv3XtHhctdjicig4A1yoeLqBcnICNnMGKEpN0nQjyXPjY2zgr+Hped89TTRemrW
CKCtsfQTDkOioX2NcU4Rim9CrhlpzyWlno60XIRX6DVzjMf8frfND/n1L6xLhtXC
9DPsQOzalThmPE5x7OUYKeLN3YfLuYFrg7Ss7taeB+0I5mnVN5jvYlkC5LPMGr2w
VMg4ca+dwtKs2L+EAD1ynAyWUIaUlZMMX2PXpPdUU8MmjZRSVSZQxv/5zd6d3eV1
f4pvRL+C8QnpNSxFFfEtm5NjQjGlJXK1f2NtP22yvER4+91Cy9MyUb4t/kIgAQpS
uwsFqyaJUxUYVlPeKIvQeBNryi/KNOp5EDGxnc2ad4onNHkKVG7yaYxv4U2pZ+So
zEEKuftVOJ4lI+6qap80g3hCDEs4GcmaFPz+9DWnAx6O0V4NHGUsC8FHE8Bx7BX1
YdKS+abRFc8EmaXUTTX+B5GT4HMWM3S3evLqIjG1WTemSiVmNgQt69CAxzPBZS37
wHYG+PbcCEW9Jdq5pE/xoNaR3evhVFdpsvWaG7nHQAMFniMDHPH/AGNSyNNNNodl
3stnsXuVIeNy92WWj6jnofNHp0VrFbCrxHiyKp87q+P395iTDN7S9FVIQDWgbpaz
Xtbzgt+yrWxsmvKBxYBh9vs5TpPSFBLhUMy+M3v0ox8kS5FqLHkMube8t1KaVFzK
EDlAWIcoyU2Uy3cGydW8gMhJclUU0mM9ESo+XAuKV32hxj7Fv1yI0q+c7cYQW0HC
JGvlWvLMZXsAdipUcrK7QKzrCfC6PbM7Mlbu0liCiK8KhmA+h07e5oSfih3jsykE
uZ3k6IomSXA52/ds2juwAjY+bbHf2DgnNDhlUtTRW83iVqvO2RatC6t2eDA5bjKp
u5QZtK5KbHiMUpBlBp+a6IO5hqMswTpBbSpKPvKQvOOyabtYoBydQdVCrqjbsCc3
aO3hL8Xv3l74j3Wet83iTrhw6uajZxQbl6oueiBa/5ygZ3oCFond88yg69zdXXQs
w5Oc34ezthW0N+AvJo7uRlM15CPD7SXoFKPRzvQiAQQLjRy1rJJ7LeSVMCm91MJf
u4n0ygusAp9WzPyOp1Mv2fLhH43zsH+lYyOp1Tkbi+jtPcP9itidiGkvFiBMKV+J
pgX2sAldhOvRR4xUT5VOGFflTF3pQev9S+c/pqQrdvz46XgG2OmZCLUlFf/MKTF/
tpw3A7s8cp3Z6XXnFzT+M+bXlm0XaA5Nx5mf947L+97du7H4OLLCnQq/hJ/FHfUO
rDyRAbyCrkGGW6a6Fbb6fSW6WLLmYhoVgiXFLROvB7xCAOjjsc74jjqOLB7y/YLl
NTU0aqC3EzlVYNfJJCcpoL/06NlmsWlxyBiQSkos1giq2Vry2JHWQ9FVxNNHumML
gYsxDGKOih0AtBuFye+4K8vgYMvJYxo0b5eVuwuYA6mBugyJrd7UzB6fRi36xYKU
DXsZTZ1rxA/DqSWEMw/svajwdEgrhsr/z7iPs9e3LzsEFzC9LJQDNL2xsu3RdaqR
PdBj1z+D85fbqgpttESKNrO+jVWWputSEc6MEgeQb2EQNpDD+eGN/McNh85AW+Sl
thEJ4wOIeHWEm5FBaSVl/f9J2Ip7Av/nd/sl5YMXgYSzS85MdPrBCjAwAlD4XK3F
8k5gCq9yhLoERa2thu6g9XsjUZUlE3vd9P7xfOpa0MMrys1g6kX3jXlquqAY8bYu
kI0BZNlFrgz0CS4a6iBmELFgRR+zW/lQ4A2fS0t56QbCaCquFxJcTwO0mQcliZS0
qnijXXOdNcOv1agaZIzEwO71WZKP680B3ZwgpaU7VRw+9CChnXfObKSaLbPE+KzE
mWgfzz7adu6+uI4EbC9IFnzD2lcNMNBWSTszX3tpx9OVnuFCKw/3rv7KtRcn7URF
azBw68KD1UAjf7nQJKEBUgAsy67AQqLb7TOlxI6m/D56dWwJDWURZN0yWJm4048B
o+eCAfAxqX+a982Yjr9i5LGp4/5ODF2bpcepcYDXoOjiIbSSnIShbQdsAEn7NGIg
9R9D/GgWrtaBiOXD05Wv92fE3I0ABDd6K5gRmQrj2vCgnxHvU9YQ+lfzA4yWUJXG
mf6cXZ46M2YZQe5Z5nrGPSDxjLx6Q5Xcv2ppNuq7ZDhwgCq1lnzv5SUr1it3d9uN
mi0PTI6qehXjp0jTCwSJ+zZUBEm7tOaBCUdLplCCkYtOPf7ru/M7O2LX4rNHYiBX
8zZ41huZpQuTmTQEUEbNT5Ed2ew2XVvLVAQuqubBkzCV83lchso2j5aJytwHsxm8
HxmvBDc4t2ctOh9z+GmlHemFxv9BGyj6C4UaNrmWFJkPAdolxoxvGw8FR7xjy+P/
Rh5Jbp63jnz5WUpG+Ig0KacgABo3wr+GZzEYt6jy0ppzWJUhN7x8z7x6DdSCEISL
GHP3DgvLnN3Ccn4JYkra+dPz0hL/RzucIL+joqUOf36GhBPJtwn0oSsROJjeHxJK
Podd0Dt+tP7F4EWFS6iuDeo/dp8oQbgivZx7xQf708ShxcphQ4q2HfOTpT1c2yEb
yma59Q1/NR1Lz35Vt7uShB9BpxcvVxDvqHn3e2Een9EcjtdS5q6m6dzOpZX2kQ5A
I/PM45cjTj0XPh3WQjPrXIiBB76L0EnbuwHx2ct488k6/ALweXoX12YuYLtOdfhn
Q1owAFFPuZ2zesoIulxP7c4sMPkh21kqT2NqP3zP2RxV8r0cSXd3cop1crgYvIOo
HFWAMjgqTyf+JY4deBTlJ7PSnDOTkDOAXJb/eOXJ0pM+7Y0a53b40OU0a4i2rgUl
RRqHuFR+fTTXP+triGS/kprlAJreQXdA6e6u5sW6jHPy55PkhjkBUCrAYZSWm3fZ
u7GtTPf0VYh9lX6soEC+1QADrQxXAW9epVbcwgZ16TDiZyuFO+WsfLdBMB9NdYRm
2psg/+Is4x9rfKhupPVR+ARAGO75k/s4f44wufMiaI+07OiagbdDrtqdRrw2y0+o
3wEdv5B1DZNr7K8mujb2q6+t6SfXm8RdYuRSERTLkCUUZd9AY/j3mi8jzTcazhtm
Off5hT0IFrOie/hQ6egY9KKYO+BFf6UqWP8pVvRUpw8jMe9uqoJJI3imbrc+bBm1
sR42FlJ+cS4QYEaHxSYGeIg51RlNRerNAoGT+EEQYLjD5WPKr/f+BUPkH2cj7wd3
agW7GvInCkanLZdb44HSrMKbQUckGuehG4trh0Sd1QCq8xWLXrXIWtRkDwyH0BmW
tf6WWy55OeH/FarcSeXXEHdtNGkXOMrXoHe6OHNyLGJvImu+YLTQwywEBOXNNpXZ
H18uu5GNbTKiL2aKs4hZg4hxt6x224D8jkv/GhZF27H/7Nt4F7dURHAZK4jTzYWh
E3Sgvm0TmBfXgUVunmXKae0Yxul3JJ/8qEHlBnRDhrX3F+J+jACOopQUi2j63esp
sXKz9tOYLQnbGwHHdYStjkyTjOdrJPVkoSagamOzioI/quTJObo6bs7avSVtVZgg
nzyxyo974YDOn8ZW7dr98T5DUT3slNTYkHg2Pv9rRZ85ADLCH8Cxvvwf8R6Ppv7Q
rWSWrPtbds5dfcpq8E349Fxlav0Cw2itMhhPqYy7VfAFXIDRa+lFzWyhFiaj3Vda
tkX6oFVwWGzou1V7FAXZdZNILiJH3PCNNkAbgy77AR1QbQFvV4DJwpVOId/ls9jY
L0LOfdKftd7nM/haFS98NUZjII4x0YIfu5kXnxWR5gcyB/Tmqut0owsJKee98FI1
4we0FEms6J+0N51dUXA16dySipSunS9vZQ/coka6yzhIcVDg4tqjyc1cJi1zp5rJ
wzzbZaetgoNaJdjNMPoxfPiMc6TrS8iIT8vcKMle9Q/wSBH7UPGrN3DDCQ1/Bo0W
FsEVRkcSIgxTvAEaFxTLSsYaJ3b0klDuegy5RrRe2fIN2a30klEyYZjiAKFUAlFa
t1TWAJM02GlBvuve+mZ0QzX9TJFwWQqTMhqa1rAJgJw8pdoTEB60tP38rVno4pXG
r2jtq5APKB5qqqxIbQl1cg8TrlQ4yyy/SQTVv+8VC56u6EMbZLUCr/Q2ngAZzGZp
P994rf4B+7zJCIwRg8XhhXRRAS1aWD3XGd6xMD87EXcSkA2UIdt+YsbcXc/ZQdTZ
Ew5DZwC/btM+/9Ywa59DrXRzB8KuVRpHjHBozGdJwg63Pw8Kn0d5c7FQRXEznCV2
XzUescAmGqDNmXrOeLAPFtlIzp6L6DV5rXTvKAUnwzslqaBU830fAEGbzlqEmORB
QTCNgvNksBH1pGKKrwxidteUdR8/gHmA60gLOhkrHrRVxVcW9H4NPgnoo8ODmagn
tS5KADa/8Ic2Ua2L3ZUakcogh3x7uM3HbdHOnwtgPff/pKR1+7o/DkJCpl1PVCul
5da8p5Zj1MUYvOWuYpIb1HqokHMk+K9VN4qlOPUmZZCpEqz7LK2pbFjz14M+wybI
5Eh/2deVq61vOMcYV39L0hH3+NKrnV6VXwVtzmB9hHMtXMeVz1EMDz988q7OP9pc
d9q7bJD1RFkRhkf7/LAUepRRseNu7yGYiN3ckmYcLECP5kzpbGQJyAbGWBtwiJR1
LNIBnc/7ZqQlvyL30tKb0YNA43MOlAmIq8/t6GS05Fn+n7Qc0MoChKI4VgRroqXG
D1KrDa4YZjJhJQxcYlVb1Lwvjab1EQgKv2i1Ldm04ZgzCDrD1jY5e0dLfVBiE/3B
V9JWr4+IHTlqvLtRUVjZuqn5+zR08ltAqBe7UFluDIKCaIF0NWyGWF07U+JoXLRy
Li9pFMiarDPM22EelPS7c2UcyCyaYhQSLShaXlko025VtmDUb8qDaV0OFBuu74ot
AtjKUq1580nO0R29doReNuRxMlH0KkvtHFE/KMslUKkmCQjKljr0+pbcbutH5eC9
C0scQ2RO23k6JxS92KFol6fdJ846aDoNuibn2Gn0l0Uvu1UVahblqtTvINNHECxy
VggD5zvmHiD07B+5hkKn2exRp4GodB+QFG07yCftTtEaeSGiq1VMetSnGsA/ySWF
Zt1vvsvvfT6XsUMcBPrp1B/yTH2HeyKOsYvFrPgZ/mMygZjs4/pv3RW56Xjtqj+O
VwNGCZmUZpUsoYtZUJ4fdOXuOiSqodviciBnG8aW3/9SmG0eEb35q93FDbAx8xDp
9gvaxBM3sLq0b84BV51uRCnUpFQeB/41+n3EqUUzTcNpspDpVw6ECc54Imv8V748
g9J0T2DOIuAUI9R1OpW1IBAOATauqFty+hRcgZzr7spVHWNynaW2+zPJlBFrxphr
IR+8xMOWjQHZEtmYVYxNSutu2hKj6bVIrv7TiTRdBlgqbCQY4irx7olw5Zho4fNw
vj+o1ZGWAjBJzX60/hwuSqsy1JjbgNxJS56Jdi7OI8rax/wLLeqiMx7EQZCmpJ1C
pRK8i/6ZJb3U2V3L1xJXHDzqB844gxN8CrGq32p1ZpGrtrzCjU16kDemWfFvWnYy
wR9zrpPh9+NM08PsRljtU9WbKI0BOPSq9bDYP8C6KjFhjF+wNgvJtvX4Nx8k1PHg
U81m3heuWLNArIB+YI3mBBLL5Saz4+bP6dp4tsQia3vTtAO3zzvoNgRywB104JOP
GEj513oUQ+dTowcCR914HOHlFKxxBISdFTYpZ6K7UN3G6gxel3bZ8UsmGON5KF22
r1wUjVpWBLqnsXaF7rQcTEaWAzZeP1MDUAwqebrVCl03EO1jI7PCS7eLrEgbqV2p
OvoYFGfxyZVKouf/cIeL0ZqFNdCYFMWGWRnwQLdbiEpgx4J93SsxVHQjsSw8Sbx3
fqokNovAF7rA5AaHJKdBTJPaKebxerker1BcgkoPZTfgE/07LGKjdTJY6L5ovLms
A03woQY6VnIPHqJifGRDYDjAAv/cgPQw6Hv+cUqIR/artcX4vyhxkpSzcNJRhXIJ
IetGQ103u8NC5IWUewWPvbmbX9mb0ci0awBD2I2z+hn7sa0vY2kZ/5QzICe8ci6u
ye6rAaP9nnozjIc+zuC117dCmi4JNQgYOMLZqfZpnorrooATg/HcETSJyH/M1pJX
jGumuXqAgCr6eGWwBfiGhjuVEtZdcjj5wRj2hEvnVA8oQxtRh4FFq1Dif/r5A03A
00hCQYt7ERbe93S+Y2qpywXZmLk/+sM4KsdVmbkMug9aW6aX60sLQGQR+1fFA1EJ
E2RrpjOicfHXMODWoDATyVhBEzhNdw/0CiYOGEM+nXN8n5yCxngw1GBj1tQVfGu6
Aa1xRuWc15iaSAQLRIA0SsiIv8s3oOIsi6PxH2u8Gvhhsy6freWw3xjzZEobM7t6
NBRd+Y1D2S0K51iHZH01ghG6gj7Ji4s6m29obqoriMmruuX5x+MSpW/Y7WXFDLpY
ibIz55VJvgNrIyY3qWG/PWZj6Qvew4LGzfkPgvzBXU+N9HPZIR8n0LuTzu3BolTj
deDQuPqXMtLXRuesWZJmeLd2Vys5+mbazgTWvAi/cy4EPhnCESRJ6xIzmvj617+M
fzdxheSlG9j5M412n0gMOLAsVMLOZNvnwnjzLRnRFR9IDBbv1HFKDCDGjsiLA+NT
i0eF4ZGmtxJqqajTZZfC7ufgXXa5sBbq8lRNjx8wWta7eZuC7guVRtMPR6OdD0Y5
QQBETMRsbPXQWnICU1InXBlZk45thIhCID8ydgMVbl/8bPLUHyGzsk6AaQJUAaT1
UQn5pmpijiy5ZB095EZSpgETw0Be2bSQoJYbnCDwi+W0Op8QToC7IV+i92zL5hga
hJ4KzN5TseQ3xC2nnHHD3uUWpy2+QU4rMNcgvmolEnopdp1kZ6psFcYj2jRRiH8L
mN0K1U/ykzQbpK/iV19TrXqnhN/QVJWfO+lArLIhzCAp3Mnwo12ViFcx2xnjVZt8
hTCQVlwG9Dk64LrEL1yEJ619C2LneE+0Gt/ganqXXADW1mVP97Xp2ZXGPwmPXKQB
He9nk5ER/yB0ROjGBwb9Yt7K7SWbbdMZrb7plgQv844YUbGFn4k1mL3pOZymBQdz
w/pTQ1AZzKo2iAwk+Po091dsYnIbseK4JJpNp+nJpKIXFddVExQtHrJ0Idad4Wtg
YDjU3EyArb4OfNHuVcnLPpYlgKtSeUUkO7Zn/YaoFRZOJFDZNW58lYWHcBT0uRpX
PjsSZiErePPhMUgmLjjanEulkLoRmqALG9sWM62zuglR6wcl+lLLDrEyvvpzr2mL
XydvvP4GRHhNUi9/ffJKW8nHgByeRY8O43fgD/fjFobtpxZUuwgj4qhnVziSJwn5
WG+usU90bpCs8fWcmTILTfVqWKH6Xv5mwxravoKASL4zFXSsXrwIjnoutLPeBkxS
xKE+lypfKNv/FtNKBvxOH5Lw4nIHSRMI9ton7YTD3uBTtNtfkna9/V0DFsYFLBdj
lovm65uslLm5gC18VNLr7YcZRO3NaCSZINcvWa/KtvCD4nQklXC1V4KaZ0LQruTF
Xr82K76LbXvVT9Kllv6RmGNbw9W18IL8NELCCdKx4td943PCsRjihS/Nv5FMTCQ0
9+NY77es4sYCJD6d1MzeRl1iKfy+RBr5FfegXwNO0606Wnf54kI12mHOd/WnRAzv
R/I7//Cm++IQW839l07zn0+G+SgJz9XD7PvG6gS/ucfFcXipv8XPSElFy2UrTh7T
vPaQeSh45IrxIvk1lkDvEoR7sWbhRJeT4Td41kI/GWW4WV3ApeRqqs+sTuZThBcD
054GO3FYEyNfPD36qZE07mVDfenSk+fDBQec+aGd1XdDxEg3/o/TfiEIG/+OH/oL
+9JXgpiW9X/tZD3nxqcHMUsVe8Ql31l1raMZ15Okdlr83cF4Fftb0t2O4pDgsI0Y
/m4QKp46B3eysq8QBhIFG9lyyyBydiko5nj07lKFp+RCspzOg8FO8TPYZcqFWFC+
MQTWJAsBIlgmPoNKZidswZK2ygvTAbNU2n0qXLZoOhJUUOBKMWumh9h5oqQoC21c
GjK3Ykn8Vje8jeT54pUsAzf0m2KtILdfjf4mp+xKhePy8qE3VyoIDgltQA1uGF+Q
7rLrF3qdq98HNoAzrxXLad9sUXtopOFy9TGcMJg4ivB7CuDlwsCyQkhM7gIGIsZg
koChHfBQJM3v47YpBWBp7U5iVN+vXuhhD2w4nD/HNPLHvSetWjopsjsn/lO1sXDQ
oW+EOYa75H6gMlYnsj3s0qW8ruWlErSzT+vbEnYdQMzBDjzCeV+GbWcOr41kRfe2
bjwHqrucH/hvfNKuPdcBNJtsMM5SqRYyz6lGrao6o0PN/6fCvlVqVn+yaSRR3Fcl
misRg3Fd5v2KcHAYPIVoht1X7i8pqihxQ5IPWCSAw9cb8KHnFhXPbmNwlc1k9atD
amuLNHRMo6US6mF5cot1Qq1FdECliDzU/R6tq2Dqc3ugjc7nHqrZNyp2OqliiKBJ
A5hnPH2F345mDAfZLcRplEkSPLyjSDWmAYDff/Tn9ofL3IE16maqPIex3NWNOF+G
XUVh81vR/CbfY2shKzXSTRk4YWqSFH33/z0mPiCnKC5Xu2/CxazaKPDt764fZ4Wx
f+slzMPJm6rW8TSGJH8p7SGbDi8QUSaDyIipSr54XXbtLPE96bhOkVFYPIrCReaT
Jkm8eG1BJ8dNurb1OPiYChoWG4rh2T2r+e2QaMjvf8nGYM4AVMEclHkh6nVqHX/Q
u6oHUddXIVOpOM2cj2Vrs8w/KN2uStZH2iTaGT6ubAgJM4nxUTpctc3le2H6WtWj
KA9fYmbQiV1kP5XzI9Y0ZQ3Oi6FogID3jLSVkUorQVVaJm5PLqfhvg7p1Yfh/JEW
mH3k1CwPQvJLrFhIV8qV5IAONOdDZG3XDcRfgwZCQ05bycUUQ+vTWuShmxObPyk7
G5J98JgutaVyzLU8iOzDvTq8uDFY3zaZOnmBI7/te3rubC3psk01GQ8nyxHQQD79
YZgrz9gSKoeXKMtwiq0f05xGV6MIAd+OzqJvBe1KLQmNtCR8Ou2NdwDsKUqI06Dr
NsRxm1/5h3dt4aBgdT/BvzEnpP+5c9jeW5saVtfi9kIqAUFRnm5NsFQoYgN4iK+i
FDf/qL8JVUNcXPEht3am/O8uX4o+xzhaAYl6D4BA7uVMFwz2GRqJ3MYKb/B04V/T
4wqsBjryt7t1qYfL1tG3iwNLmqdT9ShbL2mUQrSjd5V9y89XbBbBmNOkRLgpp5XJ
zjzewf+BjKXQ4N5EO6zGb/idBBkw5/FgUkWSTHGspamg3prMN685z1HlOybaWYNJ
T7rc6CERO/EH2MJc4PLdaheAqkhVJb2b8SKKDZC6BeRH4JWMfBF/ssPcXCz5lhg4
H+s9s2wmgAdLSVTvwDInpfmFHw1RqQ6699Z1kvtuF3HvDz5Hd6uCL6mXmvK9NZAT
E88wfn+2lmLV/AWOH8Mix4MhEKki/uWGCOAw5y0acEhXV+b3BHks7hS8ilLxRavC
7xP1khpH+bCMlNYVJuH/2/wNp30EqnpB2RVt1AasB4/aHiFzl5P0p/8uYxoVjjhd
MthC/VWwvtts8mM16o5czwwYN9rl8kzf0vBoePQFudSjConP92OL59bnGfRhr9RH
/JQm2bTcGoX8AMHwv7qD0M9AmfmFHgvzKc0rjG1r6DqLA9zQJqqqnZY7s6gYHrOU
wL0UszYddGvDIzGU5D1eh+0pI37KH8NbsBByo7KaUDeL18OBQxGRbZnssmks4HQQ
PxJs1ra5zx/LFkoEdR3w+q4eCry2nq1E72drt3x6jOF5OU0wKTzPbBLpxBJ2dwjS
k3dmcw2k6RFNcCiLVXW/y8z68VQsuS3kK+GQGQ62UX2lhkjNjvtUApeSo50CJc+X
P2Ox+EwQuSFIZOGUl2k/Lk6LQ9u+5m7Q80XZFHv61RnCtyS2ZZyq1bB0HOOX5BSs
uZpk4yAAsfOMHSllEAiuPW9V7SSpdB0wvlEWZ0+m6wqkv1rLecSJXJxwYoIkLc0v
5URwSJyEznSa8RYE5KQWMFN1kdlfochtbwWS9NuvoUJNe+z/e/lEaamI6WGUp6QK
r6OA5svJIoSXXttMsSrwKTW7eggIzhRtMluL4qSPQhHsojpsQ97duoXuktg4l6ei
7FxHqfDXDVMk5NBT8Z3uBxVThh8cftWCDpXjKSNSlb0rcQrP2eroM5EQkjTSTm2j
6ZnulFeB6KRzCV6/R4VjWgiXeSsYc/Aq5/N8GWtOgXelqffMvwm3DVLZbZdRb6fp
GqqfYxOHcdYOdYWjHpWhjsgOr+bd1lH/zNm01PdU99onzztI4tw6y4sYYfB4UGn8
77M0z8AS1kfhNAmmvJi6hHgqCWxpG2HUFpW0cIE8MShvpLF2/KGSmms0in6C/2jo
yokBNUnwfbFyvSLJYMzIm+VwDUDZ0UIPB9aqFGNeJmKbb7kC+7THOjuv6Udmawn7
yuvbgw7EgWx4iXZF1lCJdi5fIhUPX2aEjBD7Y/1Kwlh7YS06JMc+9Lo+bx9OsQwD
k92wQAfGc54iHIhVd9I8hEk+PFkJr+ZIq4QAVg8mc9BaJdlpVkd42QRuXGawW9n1
uHbRfGg8kvAZgHhy8u5PwFelIblHVqjyGkpeCPpC8LvLNu26w4APwkN5nf7WliQF
k62MKLE2BmN2jNeiKNCqVyKnd/kJbmC8ReiSH/EwV29EYJ0i9MfaHloYmxgsnrba
FkssaC2p+8QqSPie5niSCENp+XDihFWcMQUHn3GTpO2B9ByPEmeYv0EzBPrshQJf
LkTYBJjg92xHx4015UBx3Jh9/3QC9rvzSpvQP5w5hmV2fL5oEuv9oKmg+5dgYueK
NrDaIXTRvMky05L1Bm6iYWIWXvHENnMs7sH1iEbmDoYvsRQ7op32nexmYqQC6Hen
tCPOySk7KdhGQpH9mS4gSmkWTCUBMhG3Tb/hrpflxZYS3T0gfpdjBn6Iy4qmHKXk
i+DNN30ozcKwy7ldal4u++O2cQrwVkhTSdaTzlRRdiTFsWI/EMaN20DTEehufcYm
iKnr5wtkec9uWBW6NHOMpHCu1MVL60r54QZfPbLzp22v0Rx6iKDXLwr9MJty1AET
kSNLZi9BEeObOAOUh2h2OTc4OAWwdh+/qGjFMJ+6z4hk2dpHpsNzQ/qb9NCx5jrZ
z1AdUMzX3j3fZfSsd1XzZyRovoWU+s3iSdSfxeSK2FcDKq+X8DkHGx6xcs7XCmln
WFWTX2Es1g9TAIsvq/ZmfisOXfSQd0/rICRq0qMmWZeACEBUU5ecF9uxv3SUa2H7
VNwcwfYKfnBhX+Qqo2skf1wq/lSdOveTWWsxrJg2yhq7exszPHWR32iAdFwQxiUQ
osGMOxu060xjV/bASz7VAr2kS6oCFMtYfxhw0Ot72JGVqLdPCsRU7xkcumNFuMvQ
tz4AwbQ3snMHRywcnpuwG8gzTvMzsIvc0Sz7O+sXxSdFJCcPqG8v+d2Gj+09xrkr
ZN5RvngSTt0VTM5JAzrWr4359qu8LLKV56Obx6D1VPz7363lx2E4IXnS+8x9ynWM
dp/f02jQ8rsanvpEABj48Jd45sbx+TSdfxAnBcPbElKjXs+Yb/x+kuQAvRbH1+IH
hvlU/n0fIr0EWdtTM7MsdZ6XwnXur7GKxBsGpR7d/SoosPVGOWcGmBpztu4wBSkQ
vC8xmPlQfzAXVKTOez4/KfSxvziSH63H5q6aZa5bD/+eaU/2cs95PljJLrFzNYOF
6OkKzLR6xq/9C69Uq8HOphS1CuG3OZAYi2d0rlsfj7pfwabgMZ4v/xxowB+bY4hO
l+BFm2CHSyaXLvcg8brNn1Xh4Dj2933LmqA/Me3SEIu36Z11zfS9FU7KMp4wzchN
1eJgK0AD+SbjgwN1Z+pcIbrYLOHgrt/VaQhZbqolYWvyzykB1Ez7/IH0er90kHJS
MQxv745ONhT1ICs62BpDD0GqtzSxyR+WKMssu9yjvo6YBUrBlXB1HBnOBmqp/Dp6
UcV0Ke7MOwSZ++oHa9haVJwaPfUUSgKBTiLYJZUoPMgIphxyzz6Ga3xFY4Ef4NDD
PvpWGO3Br6jTGB77viN8gARX3jPhWXfx3BcP1TLcMs57rhja8JAzCWCnCfyVTCz4
XKld5yn0XiNmvUhE3q4tIm4HY7nktfw+Z46SzX0VlAEzR5nhN3b8ltfw8azVKBZl
pbNeNKotB+2zc79AtUEuDwLuNMeJaj+SofITU8K8I9EUs7OqCg2CeQcT59yCbwKe
0Ji8XPTy5k7gWn9wZL3YrDcMWCbGrx5JHO96Vscgvv6h+53RF1TPfRRoN84LXNSg
a51isKSPq2xiHjVYB/Eqc+p1vwk2waLSddyQTbcF5Hu+GNm7UEYo18iOwomavHyo
5KfHG4CEvUzbbZEDWblmwxVmsPC5tSCRd7WLY9KiGPOxypkAdGsIv+hrZmVR/nOd
WnD32maY1wKVqq9kOJ8r79Tcsff7QSqUT2gafh6wURvMh1Yd5/DU/fYWafhv9Ig2
z1T4fZ99etdP/aj+v6r1XmdxgTKdhMwMx3HBEcBl/rrVmnP/bo+5CJZkmHGJvrOa
byw19Eb4xLtf9TzTNsSMSvc3YLGUoNuRAiDoPPjI5ETXmx9pJitMnsYZqQi5bbnf
C1ntBlpPDdt0NWA0l+h/39E9YgcA1JngNR+5InKi10xb9U2lq4p7unlxnNuMjWPf
qhflqx9fdfmNPJkltvDQDI8YXmE4HNbgBvayArwEUEk+ywzDZD7H8Nju0gWPgL7V
BdQniRTlPXKHsARhYL9Rxqy5fWGLRCXjUQ3NlGfrorNM5PNGzybRZLs5o4xmbsQK
Lc1ROdQLxC1DAclql+oKCrdzyNtYlW4fFZKHJc9qsUuBdK0hpXsBS4RRAZ3J/JpR
0ultb8TMD2UUFiiTYos9SE1Rnb697QSW8yzIV+qHCFoPsJvpOmFADMMUpn0ciHps
G/qymC53PzWvT6yZ231xjO38ALnOayJZuh72qCax50NDBRmnxNvfZ+Vf2cM//kx6
hW/fal1Np0hcheVBhQIOASmIVFcoNMTKoR4xaZ8fTtt5OcA6J/2ODaj/chTm9Vdk
mnxX7S+5t7Nx0VSA0YkfiZLaKTjbdSKcReC51aYmLqm78taaQOv/LmxUmltcriiH
t01fGZ1KD2fbVKxpGbJsQGe5YA7m3jx6QCewbcNK5NqNu2g93rr2M2teIy+662Do
g5TJDPTEo1Ku+eJD6X3ljqwElGOKQBLZ09PFUJRQBm6HuPwjh+d3/cUn5f6crh06
wJPcprFGxwkkroKxOHuwhxrhwznMA3StUHsLqVVRue3vLnGgDw9u0wm2D/fs5l0a
Ix33vsACN25g3Mr8B9swwGJUxvQFhgicX5XAm8+Kx+OueHFlyIre/lmwfwmxho3E
D9saWeubbkqFIiKoBUWFUnk7NnYUS91Ir81g+5D0CXE9IL05Gp6ZN3eXN4pYIyEd
JNXRzxZ4w9URZ1dPCF/mKJ6F4L77fvZ6YCIZsePrctlJvRDQYgU48MJ3FeuebrUN
cbMVhCj0sqiywR81f3OS+zOkrdt/FU2cfB49h8AeWzrEywvqNqMujFeAtAXEL5JV
XIONW/foox0QiSDs5Of/3Fkoo3YmTTslc733GBQpH8DFZMHqdyBCef/9jny1SQYQ
DfDnsQaqqG/CRVbeHeXi+DtUXUb+VlzUIibO6aAmY6SCPooqB2k/hItOJsY7a+sZ
dA9SrtKbqaMicWyvORs1usbgvqhS4zKniDujvmJWnI5vh11fd94dVs1EJaPKNsyI
T4yXTyeNGnDq9sKmf5r1ll8jDx7cEZEpjrhTs98NSibd3dbLeixEyg9OV0datC33
khOWewZEK/dVav2TFpsO+cX+T9+HmYMeKZ37S8qbRpSqPme4G59BLJuvpUiVx5AN
S1V6LVzTgTTaeqZuNAf2IuVU6JIH97Bj9jiRP58WlEAIwNlT8zbRYgO6K8B5untw
y5NyA8gPNvr7IEk716eLDtr9HqzJASodWE4HHVDSF7rl1VLXkxOGlt5g7PKM8fE4
MbjsSO7Ed7rMKFr8ydYZL4tFYdKNJOmGKIDZS4svW7wCaBOaMF0dMXrdIObAZ//I
Dat35pBWMYz5itteXCAt8gqgG/DtxpPusd/Eop8OWlF8wlu/SB3owz2qKaNwTMGM
U+3iTk7CkBf7YReIFNPEMXnMNdZ9FVViOYO8i6/fuw8iz+0rz5yf7kK+fbysYyo0
nF/W9q2reoqOls9ryN8FnzO7Sj9iC9l0AYAcK1p97HJjMeP/07utBjhFMMa9MsfZ
Jd42WGBPtR2B3QuCgtHaHHOiQc3BOFW5XRybyHoo443rdyiiuf/C3QEz1JH1H+9I
jgrtKUfotM22n8lbCzJ2tWpS2PAi6CFC4qZfTkSdEYmpMtqUFG+T8iiEWdDu8xT5
Wodd35koCXF+SsDidB6KF1ZrcrvqKWBp9hupgVY5Po8pKv4TRTsIE3qH5yqaBJhP
PgZ1SUD9KGrKQE85Zlm118YwB+VPQXfRz1MLRKVN50svl7X9vBz1f/Xcmc6KHABZ
6Te3UTGHSyHA0u2kFWhcf5rq6RmJdzRm3U1q2TS3hMPo1aCGZr2/MqDe9Aoj4dCH
CaTnvJEjZoLJz65PtFVAv4XHecSSNI//0RoPg48FNO3bZPjcSAj/jS8Eg7dShjlL
JMXVE6/F4lABK9tsBKIZr1LOoADBA48nTIGBD33yvydEayH7tFmAVBR6EeU0B7QL
XfP4b4GPqjiJYuLFXH8Y52sP1tQpWYKpCYDDnAFHdN8ZlcmQMqa9YTEj3YMqs8Zg
n6sfS2ixG6skCaXRhNx9TavcZuW9yaE3Et4XOgADNm8X6bl+eb9ETedqTdJ90BHX
SFO2XCuRRT6aFkff/6rreEaKkWnzQxBhgi1xqw9cF73IM18dS4gAHrCQxSzmo/HS
IyDjmAKkXUJfxnK1nsFK1NRFx28cpMrp4+Ff8B1fjkNPyUrwjO7SZcn2m1+r/zYx
152nwzFZByJEUAqac8y2X0aTJ2WtM+GbCKByXYOUBPCS8N19rNN0A+HWKkMzkCH4
CzWTFUeZNrGahSmq2w6RBNSoVd6cMZ0hAAavmWn61vn7C/z8HuC3TlYGWLb5hcpP
7IuBgoYZXb6vJ34wMrijVJHPq1jkbPNEzXNgp5Npdoqvo6/IuwLGc7N3MhnebyH7
4x4FdaQjdelIPrFLQ1u2WoCVBHrLXtBmHsgspvjVqluYmAfOAmrwbOqm+2DkB66q
am4ufWpGiw2/EUxaIccZkCoj8uzGNDgdh0HgniCjEaecMWnH13j4bldNpJWpsGhh
/Xz0un+/WZawG8U74MVjhvGmpQxgPNWfnF1XLwI6Z7nPgiD/Tct5VK+TsIuZ7P8t
8Auj1IbQ97MNv8KZk69fIw0T7FWSql+/2kwkKtDUDQTILoEfr0q5TB6YDixlYiNe
9UlJ6xI9MmcE85mK6EUEZNStQrpvF8ixgKWcZjb2fOxXHWXQUbfBnhAtdyPSfxsD
ZXz6gphN0s3Klu7SXmKvOuPcljoHzFLrwJiQheoHkxMzJqVe/4EiuXLXyofNL4dM
jbQuaGpPkuw4uCfs0Vik0XcQSAs/eCyThryj8UXV1nvNMJQ9/xXDytJap5YI1Oqd
R2piSQSvmHip8iihdRSjTGfo7v1+mS5cwQ7H3NsRJwX4pDOdDM2tdCJt9+91LxmL
RH5H0+3JIs26vYZ+jBZDYZFLFTIILiCjsRJ7KvF7pJsPKvoof48xAsY65f+ihv8Q
FyL+fmJYneYRKhVYRk7tatOyCV1NCaHXFDfx55X2cyXGay/qw/8EjinIFlYU8YrM
NzSPKb+O0Yq/pXuc1LUjdBDEVTt+URcMr3hCc+Tm72cJO5smPxGqBNHKAdpBO849
HAwzUpvA2iJsU7pXdLrTCNZ8ur8jshfDKoF6wjzT/6It8KJlj83XaNwC6XS5AAga
ffCdxVVAhOmV2KDpKNJ5o1GOBkfk7oqZQRtMEzvp05sOcGMr/a6QPWPC3bXxvHs1
3fEDY5RbNN8jKN8prih6l15qifG5CpmtpD2LcPeCVKOvhDktC7j7+pebJsd+Wvl3
wusFBwuD39dGeaLr8OM0QJBgipHHUOP1n+u4rQJm2MLrIFHuv0vPkjoVEsq5LEmU
RP7tDh/VKH2vpq670yNTPHdKaOhRe/Gnf1Rt8SPyx1WE94idyz+vYpuihfjGcVtW
sUwrv+I7uy6dohCuU+mbIKFBn/zagFpohaJ4523PwBwghGTUXlv4cp46l3qaA+KU
7yE8SKqID5MPTT1J4MzMzMBjONTeVuVsohAb6JPKz0CXnAhV9k3UzQyEk3NWP0AE
VKhMQnusCwB41+KVuyArdSFRSaySZ/rNHEnJL6iFz0QzylKKqhHkJuQpjIO7Cgwu
WIpoZeLaoYBLEVywFFozTgmkTrjZAU96LWAGfmJzj8MEEF8VbQtaqNvZ/b6ldIgQ
twpfhOtmi7NH9Bqb0zg7io0sL5hQ/0HON8G6KyBLiTRmWbHnOSJYS3rEMy7OFNN4
/d2R//UB2KrYBecZXePc9FebiFSU6mhoiBG2tq0sFTDo0qmFkUkVFRRjePabfHP4
09naCVre98k2lli8KKZUsqhKPsFi/vJ+/paNcAdvx7wUKiA7A3qkXtwgTQlskN9l
eH8/XMpGiA8mPr8OlxaK9An6vpkIMSFCix+2PTHRP83W1rjVPPtftOUJablq7oaJ
fveqrNwklgrIPU/7zfhgmAT0LBGUt1ZUsTbe+YyPXRfteOMw7p7WxC+mKpaKyUwc
mHjF6gjBYnJ32zm3LqbYpGtsawxWrCpxCpp5TD0yNsDLg8QL2Rv7EtIn4yCzCH10
p1IoRY4poYiAiCDx4Ox0CHzUdbGdoIX05UYbRG7LbJiUK6E6e/ZJzkoo6PJAHYVp
QhT9ta8GKaQK+4xhO8DJXG1DGjISS6mFrxRmTy8PK+Z83C5aeHX7v/R9raJ+JCAN
km8rm42adDbAVlVsTJXCq5Z3RDCAplZotYOQclEvTkmuqc4uaTUrzgCU3NANEPwB
x2+R2xVJQRaiCWz40VKTECTx9k7MgWJVC2grZxvv+1DwbefM/KuHn2LYgSnK+wm0
EHGiDkgCXSLjoQICBdZfJhPIp2vOHVy5R7gGKP/ojst2roOuwlfh+0ifum79OzgL
e4l65oH3x51pfOzyp2o+YI56auVXwQJhCgnHTxCptw+QgwFNE9uJHk3nEzCLy0zC
EjiJ2gKxosvam7gwS6NMas+duLbqMD13JMilA5I9EE4GzlVlKx7ZwWXm/71vyCHb
4GG7qja9PYvXFA5eDRrfrCba/LyiXAZO4jJA3sl2fsV+OQlnmnGSxDP3jxVknmoe
/OkS2UxPQLj8zfDC29EYqG0noA4AItjDtXc24oF+iQAO8V94OXxoqHopdRgO0dej
59vdavnUhXTDDFRSh1x7Oz09vWQftxaTg2+aARho87ph+1rkWlQuVliDk79fftiY
kmxlNAhnUgC/By19rCMlp6H8jgjYEe8QopT3Yk/vz1s8MB9AkCqoZ7/amEB1KKtz
blXH6Jh+9GNgSCN16GQ4em/4JAxOzZW0jeHpigyairEXGmQijZ/O/r5RCYj9R5yC
RZPPW9OGow6lKW/o1Y6KDf6Kws32xczw4evVBontCenTIMj4Dlt7lP4wJoj/fbtR
964Atsund9+45gq2jPizuEqQDDLxn1wC+T2vyRJvlIlamHq4hPP2nrfVV7pGhPnC
FO65WHCaSgzHAzIBJWKKIFIN0a3Qi3HEm4iOu/DRNdSP8RjuaxaGH8XhtmH5zp45
CCwam9tKlwW9JYTlSzhzLhnkWdP3YbeAsIWnf7qLyigvOSyPqSYEowFPTajG60ro
ubaM1xQ3wC5gOlEoSvQtft0HqyGcg5jsNlYZ4HMJIyB9+Ny6beyVIYh1/u4FjWZC
S3wsuzh2CMFmIBIFlsARva1k+rzhov6rCgAe5DV60IiHtF05tlrC4VZfCqxYKpKR
StEpT5h/Um2DBYnr6MIZWwoMma4lY/tciFlnLgyVnhut7dkpCWCpW9p8iq6vLgL3
+zRDv2nTaXohvwM0v8aZQNtYriGudhsTm3pd7mzMf4NMf5fyaCVeZtKiwEMADQxe
6Ak+A7qo5VMgwO+pqVo0EwJpuaB8EB96LuWqWzZk6gTqJK9u2uKqBMqer5RsAbIX
yyrwIZr45oTPbknt6Tziyddw5TYReO2rua0OQv65PQZzLFQUjzLkLxq6XxMF1lhn
NxljUDvGGIZ4PWD8NBDZgjW7ROKtYP5AeoXLZoeMqaSANFJl5x3R+upiGLHFNllw
EufHS7EZCSX4iMgPwEHKJa/dKxaj4YxaEGpGHoXWY9JLeUDbSiDjLgB6TPo6LtNS
d9unC3uceDPBwKkG59hwPMVP9zUlEQRk4Th+9EJt6hhvK7TrxrlsQBJNfF6hZoIF
Qs5+rl4CtEpS5eUdtjwOyZlcIAF1up1bFWYsy0EhILSwM7u+hLaKGd0KWQQIrDrT
DF0+hcV1Y3uAKPVOUSF5DEwwkrhN/wTRV9qPT389MuOizR8rKj/qrBAf5j/TJK8D
KQc5sA4pihwL5pvFM9W5JBhvMK12cjj9lnhqRokASO2aopOeOuiR6B/YUwKMmaM3
HdOWDZQq9UlIzFYOpNUYYZ5eiA80y0pfMT7ZW7Aj9oM6PAYMI6K784Q5CLmYnnpw
8K0w2IQJPq2+2cNU/qfRQ3X2dlQGFpqj/i6UebOrsUdH9OelKW3RsPGRnI+EfTzr
3fzWqPQSKnN6mFNSS16YEa2GfZA4grKGtbzCN+4GBfORquvb98ydBIbgxHDlJDeO
Aa56MPok2XKKCABEq3atwHNtuaTu7THzNsm1G9OUVD/V+27PvhEM+67j6T1aJjGb
aWP4kWNqKOLpCEtf3wuTU/sZe8xvLovQtki85ZI0ov9NhjHLoQImUjugNd0sQ5Uw
ZWVx7yFgfWcWW212Gaw0RxNvzyrjN6hnQJp9p1yd1ncNzITT15JOB4nJ4Vacz+6B
9ZsBDr4JJpz/oN8z42gnBZzdC3wYz7/GNmIb1DuPzKIibMVEhjlks0AvSBo2ljdj
qstqSXJf2NyvdeGTF6bwBNDYGcLa716pcIMqK8cJV7ltgBGK11IY0wxNyS3f6Fmj
EtnUqsuqU97BUJ8tYUE07wOarYjdZWHcrcgKgK9lpYspo/EOkwqykzesXOeFvKEP
dUcs8IUq4NOPgnhKjnizyMzGhTNoKjJsDzRV9E0cwOxsLsGJtQykOorYpb4XGYgA
JDgzAKuYJnjFOBLPgkbGK6KmM7xQyszHf1ncUox/44PebJKqsgz3+OItgY3IxLr0
c/mTvtC0WCb6dF0+uexiT0ugexVBPsAMsBeLPt6rJytLcatLnOpk//ZM+KqCFd0W
Ab24vl7r3dx1yeQTP08cWroWesn6zIS7xJDX8G4Ns53jIpiHmfA/J5KSANJZQNHJ
HgJlzri3VTiDUhauZG6X6chfiKbc32WQvy1nW6cH0WYcUW6ilOV2RlxTB0f9eOW2
2xxmhBjcBsjQohImbD/nwGypvGVzVmLmErKLJIBuwtD7TtahGS9QURr9vDEvWDBy
S4XdkhD6QDlUCYRrU5mP3ryuNt0LVC5gf40x/bp14adpfkV00UjVByikiWex3IGt
zmH20EA2KazYfeBvvUoLYAD6um5ZvEQ3KlMi2gBz/O3fE4QJjac2NNL1p3lqDO44
FdjzyBQcxPRtZTLwNLG/N0sqS/YFUVxkynKMwQ4oyhHWpuXqWQSwDQ2yvfOqVE5i
6J5CAXvbqVdZSHF2ML0C0PqyTAUNIPu/P6bmiCwR48JT0ZMo3tfb3oseJ8cXltx/
xE5Mhg3fAHNPaaiHQNn8C7dCcyLzmjN5Ucvbp/y5XMsdDZZFR5OGj21oGol1s/GD
kyBBW0WyXWD4t55KWrJ/lGkqP0VrRpxOFB0OdfqYSenWibmijfWcVSXHWMMBTKy2
6nl/tcRi0mh5Y0tB6l8Ed/AD6Ri/BO4Rrw0c5H9IC+yhz1sBLSf1AbVIb+l779+S
jBBvPWQUDQizUc6udCQUcF4u8026N/xf51FBU8+46QDRiGbUOA9x8yLJfRi4NFtU
/4hc8eebtWoH1Zn3Nu77R921Ugd9RDDDc1O7cg+1uvopb4bDfKMK3a6GuPw4snEL
W2APc/skXrp9qz9CldVA1X4cn9C6lkOXrw+mVZc8EFyBwJW/sbDO+Sq0CeeWz0XT
jXq2OwkHdSduUNgt6jFsblshZ5UszEjuA9T4zNeEnJ5u49U2ArCQHBC9ouNWpwMI
/YrwkUPFhEosILQ6KEcEpBGKW7aRhPkxlITK3Y+Ed9c54sVc+5EAeCpZbdrbdSHZ
EQwQvC2/zhZKaC9FwCuMAHXz2hblZVUn43wHg8tY5zkDjXH/NIvUil6fM1MdkKU/
nRtC347uze/+Aj0DLhmWH8YcBwOD06q22uUPKefBITcLrV9Qtri3jhhpLtGioSSQ
4aIzROSJtxOG9Owy+amYYW2KYp5Da3tlCacW2HBiZ2sNC1oYmzugnUYlpprGoVh7
6OmJrQdKkIXf2jSeyXTJL6QncFYuNYFxdHHdKd8PvKch4ItE4XIixVp3oXz2rmbM
PMoRkaMaTNz9cUuiCr2k6+Ec9K59mIx3ED0NK4gkk8LXmxM6ZQMIiwk2qHwfSzt/
VXOWuZ3wVUuwKM3DFr6IeBCGspBMlHZRhRJa+euqNG0fS0rJ173DML6oYI8aTOMF
YM718E8kpz2irNdvRm1QDnnGNLxfG8tSqFkmUJIrVLnl1gh8bGsbI0TFGeY7fsra
Gevw+/jzeFd8yq3ngqemuh7Eck9txC8sBkHxBxf0B+cuU+Os3NkWL907yT5zxMKW
qypK8gfXnoy5F3ZeKVygkoJYTZCThTOs+R0/pFghGycjB1j7a3Etufe2VojOtudL
6glYLbaXF/tYDn8x1OpwULtw4yEZrrD4yS6RHkwf8en+5JlLBRnxaGkjHBjEiLdr
m720TWfTtLPzEGNBPOIzkEFzTjJQE6+TDwwqwVsR3yu2TQG9Z882sF90KLw0KiIq
YEoOYcvFteaARbnJc+Yr8tdaj3/GlNIYe1/XEk8PALKWiIanMloPuP8lV/YsrEJZ
aFj2Q48gb27Csqrn16j4UtfPAU1XmTBtp5Ybf3bSkjyQ4S/dNpLG2eRAaIaezZUV
hurox/PounXuPNQ7k6ubnMCNanLGEb1iwGh9MxnHQQfQjgWjqClFoTj0eCh9WMJB
PH/HELUH4WaU0kFFRdqInVHcdD7/GGb1ABGLMqtnF2j282LIFKAUXO6f5x0GsXB2
kKfODbX/qSJwoD20HvkPPy+/UcVKuf5UrtdUDCUZeNg7DfcBDYyHbTc3UwI3E2JW
wFAOFQXyJjYZeG76HugWlCkGibyMt5bUsr04N4PiNw3+L5Jd8/xXbeh5Nga+a/jN
4wqErZ9GPOKKQwXHnM2EpEjVp0jiSyW/IgnKwV91MGZvk4SXey9EgQf/eMUmECqR
SV9Pa4xZTP2bHxjPERD6WK4BOLjN8si4/Eo3VVTwD6F1acsPeMStyc1gDj1DmJia
E/lrKPMErz+iDowIWwVMXZCIq/0gO40VgHPJ4X4yEDZI3sLX2fW9N978/FINYxL1
bBhONt/B/gMi8Nb9sBQCbehRnv/2Sqfg4RSAZzaimZiFj73Ba/venAUUfkozkmgM
WJYugnCMB1W8On0K1ydth9FNKFD+neiGscgJbSylKkVPZ7oc+DD5QWqw8FSasPpQ
DIZsmI4EhV7Zs5uqE6GVia4MbT91ynDkziPZ066IVr676R8aBZj9yYkzc+c7NjKR
mIy7ZbKUmrq3rrfDDnYInSAWpyvj1+Uaz1vU9M/ZFOiyfvAkIH9AWFzKyiq3h6UL
ghkTdp0Z2pisJxRcoT7siTLRA0R+9P5o+O5ezsjN7OwyF9EwwSzXmrO3HDt8kKXS
LOq+T36BWF6cUv8u8NfIMldS/q8OINMcymW9ysSSD7JkwPrBxVgPv1hDcESs3BgL
V2F1XinVoIKUGWsOWqbshXqZ3xWHQe4FoVwkKnNIJoNGiN+8+c6qckCFYhUPwHZK
xcmGQMClybTbwxJZe78Yjfwiw3g57AaQJHkC0dEO2JfGggquwq4dhMPWXKU5rRQh
Yp03l3s8Kg1qI5IflTudIMn7yLi3S46ewsmoghO6xcCT3/DESQ139M7k18zeAb0Z
d818jPRselGUYBQVPbcmemeUNvn6mTrYN6lcuCDGU40yOrmgE2kIsThH9f4W7Jw5
dG8v31GSKnST+xsuAoM6KP5SCPix95o5qk9E/s2yD90LaWynZZJTDRykQFO+9inG
6ioxAeav3FhHUrBV7o9WDqoELTQNrajF9YM16oOPdmSTBQaHLki1nWe+68Xg3BDs
WNOXwaqs2gbpCNEYJJGiVV43E0bAvCwpFuYoBBpqTe85hpI1K+6ZMEFvw51/H1yJ
fcxbB8kkavFIA2EtWr/eLvmAQ2tfQ3l9pcvciOMkBfS4pioA8wHF1HnCAn74AfMb
Q7o5jDrv87aE4OrTNfDBx1pEoCfDiYDjZu0oT81MCZvSdx7pO5qcPMwtZiLRuz1k
QzcEZWS2v7ikp0NMJ+CMc/pB/A9C1e1aRUDet4QdDk7WrQB/KxBpomeSVjVuQDft
PImJvOpfYfuhfnPvV9OE4EilwoRatcPZ/fA5WZqTGqbrVlSFNHw+RhWWghrLsxDO
JsHojKYBZPBQrY5gYoLLWNqcVZnaIWVMOGxbnkSYUV/jYwxS0pyiaeDqYCBiUk+v
hRDyBLXwPjqsBC10zXkKm8dqqyNKmQXiBXk3nwxqQ1+30Sul4QHtUs1EMmiXNnNg
GQ8MVgU/O1BRjZaMMOGQAofDBI75WCC0jfORDrGts1cNEWUweus7J2cWBSWiz2ci
vJ7pZ39YbW9rDUvjSVGFjBUFgUEiqYnA1+uD528wBRDeEYdwQQ6aPbjSwv2QjObE
fM8cdtGIkAnP0B+6NH1Z+6y3Fs56ZWse1MXtcQMo1FjoJZq5+6sxYCB5xajWodbf
V+yf2B+wrPKbYEwGp8MXzTKjJHoQ1FwwjlmfYivclG4bvryc44KSEotTEhV6+loN
Vkc6n+8G+tFgfXua9Vnk0y4agnuU3ujksr4YuaymT7dRY+Bs5saHH+5ydKIC826h
EJJ2hK6ppzY1ROgEissGirh50j/LC2OFYl7IWn/4pcvvWtseGS14B7RBonERfsW/
BJN4RIuCsUcAKowrHWv57e0dBRr1Qjmzg1x3is5kLkicTXNKiu3KNREyAd3vuSvi
qJWLVVUHbSQeP5is4fguNCxBCoseHcFqdSVViUn+UuKZbhqFNhu50mi07LQGXso9
uI32chXNXb0u3yY9dQam0eEf3KwV/F70192FJt4jdCoijPw2cXtlAsLmDiQ34jBY
oGaolgqajB6Nmp8LTdX3bCJOgEcjYAUb2v38buUX3vIsjOY2aZKycogg1yOaxqMd
QzNGNSn93jfkOq6ey2LD4jae1MgPmNP4Y+Ab5Ls1f6usox9CQWiS/K0A1jvo7yL2
i9lcSvCtslBlhKTdgtg1SAoDHSKboroyWIxuP9j8QOW5yIJLDHRZMP7MAr6jyTSu
Alm/d+VTqCil9uzY/usVhO/WdgEJk4C4KdsIAi1STI8fBn6J7B3siPSJLJErOCoa
AaLK+6JX0DFKur9tDqaM4KPGarK10Ec+4pjPEU1r2OE5akjXn3TN4pRm4wOUuEDt
upUwQWcZf3f/2/rds+kfIptHDuxoATGppCBUd+wBYuW/AbllHnhP5OSsr0WHWdb0
3VcyQaiJIu+5M+4tY/HVZEPH83/kh6V3QI9QgWY8wp5gPjlSl/Z/avAXQ9KWv0vh
+PFGPi1uRys4X8fIGRFsUgcLnJCAwF/dbQTuyOv97IXfBHTngxVoVclm9OJvWk1i
cvUPmBwHPlhb0VQ8ohADq7QlcWqIt881hlknsa5MR9ZaxI52MAunH8krXr9guBGo
6WdgCkCG/U/mUHTt+HA/Udh4qxB0Nh7iDDmwX/FtwGk340AiDk4dBbhvnsPhzfsf
znbFnTp/leHqbgPZq70liY5/R9FQuHvSVSEofVthPXrwtpLFJ7GL3HdwgZmHxYU0
47A8DveCaLpGapCPMeOSf70Ma343QsDt3/C66GCxwnzU81j/XkuUTrh90qz7gETx
hsecSdZxz6eE5pYjjmGqDy+sAkkKbt03CtksNNgDluMewtpdHhhFLNJAFEIvAEOo
T9BFc+WZ2LTl53SZbjzO4a6olkCIAr3Z8q/+w0Hs1wkUzN90Y9dakKn7unVvJ2/D
cnHBDArZVRNfQ5a4zNhMgq9HVMjmSGQm64ANtPOYvMKB6XBC0t5oWYWN5NHsW8M3
0TM8XvGCVLypugC6rCG4g7Q+Z5+bQ62PIeUblvDENhB+rw7hKf6LILOD+2IcCwGw
zz3CigwYz6OSI3KGaMy5y7sk1/Loae85WuVZJMaAvb4ipAjDFwYxtAONBv5yXJK5
CC0cm1l5eFdFM06MdAIaCEcMaErQ/XBPbbFAFxZ2ZFe1hIBgB5Letk+IVvXNTEnS
Ebg07+JWPYFperGpgDYLdG3LxAAm2FZQ+tikIarSzOURXX2tGX/r63vGgMBTwDgp
pJE3BrMHqrq51vQ6iyMoFXZXGJafyX/ALIoFxfee/dMMxuj8W2m/X+2wQFq6tT1p
d58rMgX2qP1wfdzAy5RpsohFEaeGHpMudgJqgbQtg+rhR3tR8s4tz+Qui08wJXC/
6oD68Lb/X6niAxMGOL/Db/ldOblmyAxWZLvJCZdYlD2IhRafSaIn1iXsphXd2qBv
TCt463nhQ9l0+KIBmCMoVF2R5OyLlKO+Mw27DZqFQoF23I33WlCp3OgnNcRpQLcq
cuGTqPvM4/DvxUTZaSayQrPHI49X4dt+GnsIMAJZEGSZtw9B3rDttkJL4+SD8ufW
ohQ+HqsV9hYWuHf7S8EHqjgZkb+Ap/oThLj/Ha2ak7FDQozIW/J2DtzXyPZCjFVh
v2MgciOTmz1GQ2p+TzR202PhlCAqlIubkfmm4esuDvAMGEaYuh2zOIWIM4cazCVU
eRrG4BXj/6KkOWPblppA6yMrRFFgJDbOBGv5Tf3m+BTI7SRI3ysPiyO0FicOmYka
pPQaMLU+9jb87aYQwBJ6rs1QijMUvjFHaJv2Vp2yJT9SjU+/PkZqLeQRHEpQt2cY
YV1rtrpsXzI24ZJN9lZC01/hSOvdmmyYrNS4nFeWOGwqi95SI67nMrgsNVyYuvT7
66hFFoKyZrvUacP4asTemzKTcqptOY+lU44G72/HxsFl2N0+OMoUKstdAv3X/Qvf
pqS0Rn5kYXIqYMSC8RJNESkxSFv3z1jGGEHTKIj0iS/VWeYp5odsidMN4Wf5lmzx
4Q9yoRqqXtQJ1yWcWKFTtUOLzLtoH22tPWfl3ui1xnMjBDwb1wTc8AWrri6ls+u8
77ApuTVJcIwc4cDohAb69Jzy0Qv6Fsm0CvIFoBnq1wDsWjjtzWnIUeJ1yl91BL2N
XDqb++wPSopcZ7KrQ8aIe8ibkuV8URrViwc4IIdYnClxaTqbCWozxrD2Ogh1V/Ab
2XmyKFXJXIa6osDvCG8T5OCDD4IHGEOuWl1XugLGM8h1j5SrbNoUF2wi8jLdrZJS
P9CQDVBwhX7de5m9HTplDldk5xRWvBQChVWJrihJquaT5RlejlajTrbsr2Yu9zFF
yVYmr/74Un1Zo4z84/QKzUmfhbt8vrEilmXT+bFoBzSi/iUfmUVKtyZm5TjU4FXc
MjptZclyLJeqGX/+3Fjea82ZL4+uCaDaY+afUBhjmqyq3+pbDEMl2eTyWmWo7jUe
gvds1yeFD/M5qzY/hznvdJLQmYjG/QICGVSOPlMYu2LeMRhEMQfK4pw038bOjN+P
clMrX6VOBWF11uExJ5Dt+j8C+Fzjbdx+JmTQ3IDtV51pl91Gs7JOI8O7QXWiEcuO
A0054UCIH8N+JfKC0hXFWimqqTc8gXBrBUwQwTh6kKjdemqcaQFCA08TRh8wE1N/
+ejKgQauXm1KvP/Zgjne3zXhsuwGXWiFZNJ6fIMMSDANe9H4Qk7kA6Ws9FyHfoIC
0AwmJkxQn7ZX3KFsUIpXNjsWf1bFa18s9HLfj7WjEFwWqsoKYH9BNGQhd0QH6Ksp
7spx09vGHdon3gEFod5VhhvqYhev/bluBKzMOzLHzaX0xMxI+6k2+DAfx0/WsmP7
SARSnDGA4+CwJjIqyuuhP/11TgnRSOAobcSlFLUkwYrM45JYm7FJsS/xnvvanfiU
zow5Iu/e+3ZlN8mJWuIEvaqUMMB74CJGU370IhMwpdMwdiGDHmCNBebABvEdwjZ6
O0SaEVogKMx8hijAB/dsDetQmtV9Nq6qooe12cCM56f5A2umTnCSuMXrgh1AMAp2
CaWqTheb0FYDfMSIl2YxPvm/NG9DOgxL6PWD9AL7DFKvKh+XTMiUI0AK1pQEHvZh
QX38AxLQ3T6GEdOmnS+pcpjH6z2OHiM6dDl+Vp85x/wKw7S+HFXFO1YYhqwGazsN
kMBTuZyZoaW4tkAE2uwO3dHhPReYzsJ6mQMRlpCgwoufHK8apca5qOSGRQq9E5mc
Z1biPs9iAd5P1byUErmy0nE/oAqed93GncqLoAl2oc8t6HaqPaC1c9QZKnPd82Om
OPSdMnSZG5VjRqXkHZDeRyYHfmr2msz3xT6+3OsZELJNc8Czn0Pama5Uy0vd6JUg
8BbxfnZS4ZYMSDpVQiRIyNuBVwr0WC0zh+04FtoGtA16nHx2hRR3x0bYkkuBEObR
eSPrfKB9LcWGGgpKPOsyXNUrEg4FuXC6FvMG7FK2Ac7nn7dAXfb9+X/JfCAuvlvM
2A6cVRoQJ2JenS/v22KtuoYypTJt9HHbz6D5CJr62B0rnIZzQxlC5MTXBwfJ8+yW
3aWJ2UjkFx5wT2CANIY5w7bmzpZm0gxzOtFtAlywcq4+4qlSALXASTcFgb67/89C
JG7ZLHwkL7lOGnMEvI+ceMt+MVnYw8URYme934rLzd6LJjENZfn3P1yxYAvy/85j
6gSz4Aui0GIH0AUGgzukbeziAJR6O5nGgeIguUF+6OSkEYy6kRaMYYiZkXHCGYUt
ZjClpFtDcuLwUqnz8FLHqS6Cil6Ks39vj0rUp/+bVXm2CcRgc7BTZOfPqn1AOgXJ
7SBOldNJmqtFhURZHA29HCQXMH1HXHoepUj6uc+UVj/XvmEV0+yZI5zPLrL9YuLS
NzMb/dwc/A0MOy1vUSXQzPV3pr/tx/T1+rl4Uip6B9JjOSgvbXHwleeamTy37P1Q
yroGLxbhWAkH7Qs39EqnIcBuLEi7vElzyx2sOrrenTrj+hR4FR68urXeWHWB15Wk
ryy/1FqzpfDYJRx3dfb0jCAJqLwwNri8GuGO2EjZc2cn2vwV4WF9A5SUb/US0B6i
5T66pvlGjPQWR2v3sjRK6L+P3aVU/SeKEqkn+B6P8KRt4teaHtCrIndpT1q3BkH/
8RuzwVqL875snGdRUsP912PHucSiKQNWYPLiOO4L/Xnp86I3CB4bYX/U7AWVIBtU
McmhGF2j9PJiZzfnRqfxmlDAk7d7vHc99uJlEoRWgZX1GKZQozLzS05w73Pn+2P4
m6HKgW6rpNFajwP7vdqOnPslmJrTNiOwRSodJz2iu5uy8KBpz7GV2R3BcdgFuq2Z
T3Xbv5FBSuEHGrKmRJ0Ovbbu103lPF+2xDxixduE79e+KwxKotduNRt7cxtLUUZF
gb04riJWQrOmPWntjzueoXYMDaNjaurWp1qCMre7r2alEhvvxRqEKmvolEhll5P5
1GonLuMwttOYDMgQbIojc5xiCqE8ED55s9owfPtX2sLz+5IYSd8FvUM96tDmBlZX
Lvjmx1PMuxbzQWKsg8d0wUPg19Ykai3uAWEq7dQyCF3EZclepJXQvjooY4L8Klc0
D1aVsYcRoL0TWjQq+gHwI43+bNzdeGsiURZHDftcAzwaOaFlGwjerbWYr4kxPmDL
u62rnt2VP9sbxb09W1d2lK5e8N2oaMBqHbqxrCeorfms4vCa5K+4M0acdNBKZs2X
wPwaoXbh7KcGyDPunKvXK3cGxWU14TyE/jFAyqLkwXWMfqVe0TR7xa8zAhWKKali
onSCCdhrQrSlKcRaTqoIociajPffkzKP80KPQgD9L5sYKYIq3sp520Oz9QL/Gpib
td+6eGpRKmQMqpc8j1D9vwfJDdQPYUn6MrDeIKF6YYTwtgXQshsrPwvPPPwvQHSY
uW+061GR0+KWQ5bAQYAhE542ZbyPqCzGOBEqb/6HpUzcxAQzw9U+DPAs1UrhNmP4
t+g/IavE7X2raocoH2fAYkLqOsDITjFtTmyOmHK+Ky7voAI68DvbmQFGgqIDrphI
ToGri/5j47JcYptPu4pW2vsxzsUA2YF9dz300diwomIsj7G5F7eS9I6tjOmNuCNo
EKbswIJtfwV1TO6+FK0+ACODKI/XrbfkyW1z8rJ/7F8Lc9l/jne/lU59IT+7u/g2
xbft2hpLghBNdxv156f0BptCO2zatnVgWaKeMhUqGcSjDriulgKSc4Lk02fVZtSf
OcFf4Z0eYDoKe4c60+vM9HQIOsQbEFtw7FbyPZ9o8KaWml6V8b6NDcbqjWFX9ztt
0MCzi9wI5eD/Br5LO8vQfpQpcq/ezFebOnlCwz+OdEKFBRNdpG79z5/beOK9zQEn
Cw2nI0suEffyH5sMIOMELrrltqT4Jrmkws8APjlkQHM2KqhyQ7Zc8QqAUGEyUjjS
7qJLiFd7ZuhPB9NVu9umfUDAULdFpjZO0JsDPrWLibpKuC6WI2RfFmuTg/4dRFmu
FsY3QOwvrtZdCFLIGvq3BYoHYzQjAxuOjBGlEE+p37CvS/xNhNhP+/JXopk0fkRj
YJ2UahqxBlHQ3lE1VO9OG60N3V6L/HHSZhhKIBGAhyggWLlAgcA4WyrtT9N0NAsh
9fTjENbzex72atuD9Oz8+cFuACm+2Pfdb9tcPKflULhO9SzpMtL5KE4kjeGLjVYn
fMOM4Z2UDWgFF6tkqy4h0rWBTvWYDs/rYhhUHNwoLysr4FiqLP9WvebH2yfe7yfu
Izm+qjdbVRj2VczP5M+iS43Q7FoILmFZFL20jppJIgX87UN/Z3/TKqhe+nOD18D2
bzAdSEO/paM/h99Dx8qUzcT17bi4GIwORuVFn2Puat1vcOuVJYy55MhDuNDaeF9j
OqEo9OK1dY6XC8GOhZDlHfxJpOiRdnMMLdRf3V4awqIi4jH8jh9HAPbuuzIhpML1
EgFTon/8GzV7vUf2mcRnv5cMfgvGp+hJm9ExNCmPu4UzKrfBYcssgasEKLgCHf8B
OPUI0ZUc8R1u5ih6jeuSawz8eWItB58c2nUhU+pNun9Ah1Tz0mO5iCwsU2Zvr2FW
YgNEdl52AD0cEOsJu23xvHENZAiwaXbURjC7VuTT/6yKbC1Jcy8W0oGD6A4WAfpy
UWdy2j7YbIv0L06kGxEDWeYfDVVx18v1j8ycdULJ9hS7yHCO2IZj+4SohK81WGqO
NEttFhRI+XToIREWS4DkAmCuLOXZj1d1zu/qAF/ZdeVj5ctL9mccsJtMEvizTr+y
VsUCWjUaGFXS3sp0rah1auFAQCCnXIxOBQERgDZhKWBr6udbDUz6pD3Id4QGOgJi
zhxApDaUudYBLpywioPIO9eq0NoPC7datGYEbd6v0qcK6NRgdlK5PiAIFWhLdOlc
7gdXhz/8ufvbCj7LxJ06Xgv8uSVU6Rt+JmA+CM431w6rXxyk/fnumQ/ODxhtqzGR
6HrT96BJ/LG+7jJahC4CsibTIibdRO51CxYPlDvJzvfmG44ZGZQi9o7gNaodnF7M
K9aTChDd0tjXD0LROvDO6j8hpBbKOwoG/5UnGpO9EgfSb4gt6bjet0VDi4uownz7
5dcV4Ts/ikE+gkryEHodn+gDin6PSTZEoAcTuk6GVH7JYQZXzeGLIEdxyEV9sc6z
uUpxp5+D/JaNtuvNavXn3RPJclnNYmh5VM7l3Lf123CJ+4iroKpLlEyb9qdi+ixa
OFN6jdIFoldU5tlJ7jKZtvEBfh39pee/n0AYLYQ5K2xl1hcKpCRyxNPSyX4l6dlt
JdAzxpq7hEGHW5sFAOyWkSqsY1mdVxp+L4aW9vKqLrGFlgV7pHitaTFekKdjZW07
TJk+xhawL3OTX6la/+lj1wY0HVxJE0iCKzSYEL1Rwca4+Ji3+slJ8eq2Y0T9OeV1
E+sYCnlSgfht8PYXFCfjGnxjlt6q2tWhwWuE5M0m0OOSn2q3wvDqW8xCh0J12gB3
h5H5putkPcNJ53Lmd6BhSOsstrxAhH/WM7XPCILzy6A4IpqJQbUlQ2AiO6wc5GSa
hTpd9dHtnzSJlGNQ2zR9EEoLOo9yZThzffob7vAfnppfeK2qap8HUF6FyzP7rlPh
8ykqjfk15hf8wX7LkDHIxoVKvNhpsBlemBMoXnwlFRKEccCggsGSjRzUX8SM3Pk7
FZbnKu86CYcS0tATCMLDF0WfFM0GaqTsi870GWtpg1DD4JVPVhcLbHmYolyPLsSG
j1OjrODg0VkB2rgVMc6V9sXQOveNL9js9LRyOI7T7AfKQV/rctBuHbJdLskdj/bf
13CapB6HfzOKKW8Xx2rnJaq8CLAmszbeIklzALrHsnxBwWCQzTTxh3DAg6wUOtrP
XuCxBdO5D1w20HepzBNSrkpy6MG8u1odSpoy6dwprCUYCuuSkHyIOT8q13bRI6E7
0evFiU9MQAHdOW3MvcxEe+kqA0BDh6mqWkMJyrFulJbXBP7JPlIOjRVFOWqDj5Qi
KGrHeXNG40yrBvP863uzla7QOF/LsKXEbLw7yfgPsD6yUJpvnbGNYCNHZJ/bfefy
jgqkgWVqMPMQh6JRztLFlNpcmJEBR8CKMttnbCWc7LsEbmd8c9jHgUItDjcXsrLx
mewgMAAEq/5jU8IjkxOsl6/MK0+fahy9hc5QfDdqwAxHB0TqK31Y7Yr216wiwD/M
ZyoqCtyubgzEXbiNpaq3Bgl5N8igB+ZMT+QObvy5yaK6QH3X1s9XUSIQCrkN9wkZ
9m0hfr2V7yUnqsAys87B+qC5gbhs1XYLPVWsDwlGZs8PmvGPv+ZMFMRqtxgKDxRb
o/K6F1alVNaihEGTxpT31hbAgk5e/cKr6ripW6AbypqXkZkmCvncZPfxZM5KaFis
AtpXoeSFXHiGoND2N6QTfCY1S+UemmR+2XAZHTfLZPAHMgU1JhFkrvAVwIl0Sk/+
IAEgCm9BZMxchZtNU+l+9aLXQkKY4ArX6txyslZtxBzUXOpCwAlGfBUKnH981LqL
TAzufmTE287e8yxgrPtVibFBMPBBwC8JPEmGUuoLyQiucpF94/Y+vNwFdAPOTxNy
kxgurFN7toPArNP2OGVFnWLtkcJujhYzM1jBlMalqyxTzlSXSiY/OGrDq3ePfGvq
AZNf0I9uWgUVGjNOuJUpmY1J0imNSvVhV6M8dAzfyXclC+aNsv+CTsTZpz9IYq1K
LllIjNrMaBNf7XN7drJtGuGC9Nk4tTKb3imNX/9aSBWMAIt7euBOTT07ceY94LlY
P+7Flh2eyvtGGlrpzw3sw1TPslZdiXjzpxJCf6eTRt6bglMF7zdZBtLUFZAGCV76
Os2ZNEc8HkRyBsffbzBnVnEXUShat+E/UC/Z1U0B4V8A+l4av9tPEeoeZyAO1Omu
ybsGtZO/U56BOBXxFdfIg4VQ2AO52WXGb+XJXDRGwWXX6ApSbMyWoyH6u9TAdDcs
Mr/bKHXlhFRMMDjnSuPft8KKiyaDkpl1rfF7/7SzC29qqiNh5EZoERpVEBSlcg2A
AmRjMYlTrUtFspYZLC3u6852cQ2oJFesIBMfXhZCFcmbmZ//o6+Y6WNCbLct88D9
aHoetVncN+nfXYfSVvmf1G9sWav7Kkj5LuvrzTpvE843ukM98sHJ+Dp7XZHptBcX
5735qyAKV1Axql1/+dUe3X9tEOAHPYLlQ7Mn8IL1+oM0uW3KaMMoGY79wZOpUf4v
naRGbILT2xeFYExWD3VaSUn7k60Qhud/d1aRGg6+RYI4StQ35QfZQeufcih4xetj
ShbbSVsxXFLB91OmMaKWFQ1vR/gs+czD2MOpaYipS/5/vl5QWTHBzTMy5wo+hpXM
geI5j2Sgo3WbI5tpb4C4VaY0rtKXMTwkKULrhGr9+lFTW8NiBBMt56p2CaAR6NU7
JdeNbiiEgiQlhtRCOsnourpwfa6fGAXHKyL++ac+JaDKL2wFxrAa3g9EVAA7bh/k
1rUNmPf3hoylDROWfaK+HCZ3CsGRccedAA9yAmF/f5J9tIDptEw1Vf3G8YA6LcCM
D1WWI9Y7c1a/5QPCXaC2/wJIaFYHLsBNBGREulW17JjpaTLRUs/tpW3yZasd6xxV
oFnWC/3vb8x926WMtKe6Nl2evxgq46C/CuCj5W0VkJUovAGXX42PYGAuqOW5vL4u
WjaAUV/F2WN6tpCTv7fDPAHPsEvM62PXtd1jACDmsid6evJUFC6NtMAYrgg+6MQU
YPrE0HoodPG6ei2vHcd/YZbn20xAaunZ5aXfu06ZN7PzH31NbhrdAjmRabdnHegP
be6lJhQvRmb3w1MTQHcT65EnEembSfIHz/Y+Zmf3lNPADFGsCGPxTpeCPPZP6Yps
h87+wvRa/NxRD+xTcclIB/0hBst1z34wg4/HzSHAJA6PvEq258o+MbXgTrBcdSbc
KQHl/Q1pUuth+5/WXCLHZkyx3NTrfQ+ZwADvy2gnf4wr9OZF0mDKf+idFZ436ZH5
h1eQ8/DmG54y9B7HVE4LwvvEBJMvna5+lGJzuDczWg4oPOKFhaJVukisVe+1CX/B
JfQQPI+D68HTGeU+rqUJiIzOWC94xrPD3wsL5DYQ9vrohRkyw9HxXezVhw1dPQ9h
0UEAAAekXnM+CFqCYDFwao49dA5Q7Gf+gyqycAL6H470QySaYIgX9F0uEqG7vFLG
ngI/YdXeRBAhwzs5x9dVuubeyFlbbCIILwHqEec8gSh1QNjAewKJ6D5UEMlXyX7B
f8gD9N+jtrsCifbsKm8bZpJiqe/PPV6x+/ZB4x4jaA1i16hFv++3ZLt41YqkT9nC
BocfAgdQs4dEWTbaQj6sl9VeiAbe5a/9BnxGZG4d+b1Z9LC4Xjl+tT7uliFTKGT3
LD1zUDMZvdGzBC0MyqtvK2IyuszZr2jpfBZm02UTzCYjXqWevl1tQugLWkSlNXTr
6tvlVmgdc4PiXGDNJJwj32CsgaKElj6HXXv+Mu1LTymUSh6sgK/Topx5U6/zNaAI
AoYkOQL2lp0wAfV+y7GvORbcOq/OnuCcNG58CQnQhcQqmzh7MbYCX3S6q5o0+D8d
roUOk2slNxxUzlJTzcZ972VBccRoGuhBSBr7jMoR/5yYiAvJXBYbtQNtnguEUwt4
9y+itf8qoGVfbbbwO/9QpO7vQM6dv3qO+HzofsHpgEeGlH2tumeaKdYTiD2N8hFv
SvPk8CCkM0k1eY0tbhspvRbX9cqZspaHa6FGydOALye1jX09nAj79NqbhTwGmOas
AnOWL3/HORHRP2HvP2O2RtxXsNsj6KNqeOVpZsslolhNOtNoEyTtWqzxR4M1tit9
QIezkJu5ErL0MbN2FH4akYqnQobBXhrI8a65F5jg0PeoXa7wD53go/BOd8nlW62B
7z3I3gGdYHQgbPnvgBlGdry5IGSHApl57sPst/3btTjfuCsOYPdiCrbsvvp74Uy3
Ok/eWvHTC/sp3515jWO0XpUiPv2HGDrI+yYh4Aq87GH3dfF7snRUENNWMpaVYYvO
+QLJHFxp0WNLHjkz1kAKLc0tJeE0+myYUoujJ5qh1ZWv5hVKCF1KyIBnMuVprniZ
6U7QWQv3A37tXlb9KNfryRWQanz6VoP86fejchyPZCVB2HjjrxzW3gk1SBAB+sti
jH9X75w3yWxNFFYlQ0jp2wKr/qSStxiLhf7rKTx6xeBRHZRcEnVaszbJHq2P7Ccu
SYIM8Dj5jkKDU4RZUhjpk34zVNFvt9dJqlABLt4ft/9/2q+DvIQuqzUIVd9hiQ/i
JVfp4vtDK9m5tVoQLhj3z1USH5vYMh03FNS4bGEqs4l+6gPEBpJIr+vuuXEFnfQl
KHAlHr9M0iAxgRjP/iIuXMl6r3IidpAAni5hQoBDiPKjHi3+YI8uPuF8b8MOO9Xf
cKfjrJyhW6CuPJV+/jhknrgw0vxQkEoZNYBAqceEo9z1rZ+gjQNr6OPs7Z9bkGRy
Ia8wul+OjuFfSbEKcv1zr2BmyTgtZR0XYDa+qplt1isR6osg457x8Xr3jNlR/FR6
ayxqinrvm1ABXAX/dNb+X40f8kF7PXhavrSVQsVBqdaM6/+yW/YG8PZdSgEwVkgK
HPBl++HlVjhDShu3snQxqDHVHTGNAmr0g9YftTGJ9Qwx02tXFQLpauXwVf45tX3W
bx1jS47h+U1ojPX1/a4BmDJGURIVzSmrgEmO2+OFdLkFukzbAiwsc/+yBuyubzCE
55haX5xAzPpPMzRbWpAuslK/4SXJ70qqfceYMvC5UtqDsXe9hIHD1g+3O4S49VZx
uGW1/ziVu9xFHPVfA/1rbdNGpxZoCUb4wTRlJPDva/kqOEmRI1EAPOPZ0yox6QBw
4dGkp3ctvluPlhW1dJiMWsNc3SBNhxn0WrOUPi2WC3cT4JxPw00wyiYhXkvlyYc6
uLuufCnpzi09usOZwDfzfJXlgSugooZGrKk1QdgddwV4nIkVMBIWj2TFnGFis9cs
JOS2mkBhDTu89jKD+N419h8NMeeqFkx27VMY21/t3/W6aYsym7tZyTMX+IrXb52q
jbekn7C6JEWJIUdUMv/5rprhfVqOjRg+q9hbgsK7WwPX0ia8k/eJo1KWw9gDmqrX
jCLhkUw1cmSj1zx0tnZvZl03nBN5rwdJHs8DyKa3iGAq8JoBfbKHenHSxv/i2OIM
LMO8HSJ1hJzBa92LFTO7/YhrjHLZE24RC1OIvTkA02C2ItUyzS+vMsurrm9iTyYM
csk0VxBb0DE5Enkuw9T/oSPCT1efCYELuatJyKmpZNoVfO/3jUQNWP6ca0JA/2ce
dmbe6GlKlOXtALopLvcSvkjV4TXtbuhm8/sekxGJHdLxpUgvzRxztIGZ37Cug7ZR
llpI7tQxdxuR/ObwgBb2NUyvRhWdYQAt+Pa1nXutWuCdQzbK5vyJuyt1Onvz0Che
Ndk+G3rOy8JuQjYtaQvC2r07pvyTutIvlaEhjDJRjukdVbrZxsxnACzqQRD1jYJK
YHspYdwCERhX6qz7b995JPC/csdrL5HYxUGP1LveiepsMvP1SkE62To6WNSAnkVj
9nHkTu3TzvLWnL7GZyMMKQ0fRHpfLGqpBkHVV54Ff4YY3HAqa1jy1i24L2j+87wV
n03t+OBLtN7TCTgqNavBP4CoJHAqIXfWlV7OLL0YGj25g31ZO9HPlmLUOxeY60WC
HU2Y8HLJafERd3PQoF1GG+5GFXCDxOwXJwxVIs2XTBJG1ZJyfzOm4vly1NsbNKye
2gHVBJX4n08KnCNkvusRPyJrnXjvIu8wG9u7QoMBtWM+hLc3GYqqC6WZruvthtpD
w0sK/yRe5vQ/qklms5uxDiNASjiN2yv8Dk3UFCTQ0Cx9c3wlzfXadQZa3IzL4Fl+
JBC3LjRzmYOZlqfLeAlz7DnHJD0H13LwknzlWjcYye67XTbJJS9crXZYmu2hCvDO
l719nSdY3nNbXk/5djq/5e9AKV8qkEjjOrNrkIHDt5GznmhDm/LIeV8Lge0g2kWq
x8fp73pa3+2+gDAJkj++eaYbYIboSCsA6KcaGoSwqnH/lbuBsF4AkO6N4OE5i9vT
a4evhofkK8EQHEPo7gZJ668/vk87vxKl6b921quRiKrc7v40mGv2fN4RI1MprQ7X
edIjkZTLyEyUFWY0DJ4SqxWYwnp6tS4F6XnmnH6NJJfIkwbqPPVQ4bjFWdUW/RaC
oL2siYvFU4FJuZAQ1RaBVjIAewADxpDOIhRKr7jPVkrbQ+jXzXUF0xl3WOhcu1rq
N1t5RrZQ1oEjOivptZi2K0LNoAxHErSMpVb+T381K6eiSST5GaiykugGNXnmJn05
Nb5Ykj/DkBGkLtto+BE1jFZAD54lhMJPcXl5xCg1QV6EGVgzZn9u7F0K6c+MxLdZ
xDQqwdddf7h/Om4tWb8++Zt1/ZeHWdXEsKu/84cTGP/uP6mNSUNk4wVE0vcbPzp9
PEtifn0p02uAzlnMDbHBEw7BIsciqJ/oggL1tIjvI+Ml22hHrdZoApUTA0py9QOm
cqaroCLVE5YqVSOLX4EFu3WlXXtqpvKAyYDsFBMlFj2UdvkP4zA6wNjBnr0Gjfbl
sgCZ5ozU7v75ZdG3Zhir0s7+snG+Jr/V3VvK0FNv5SCN+vPIjGILMQ5/yazsmTrX
79AOuwxCY9YABr9JuDq28tX/QykSSUWFbWNwfEszJr0EinrKHCk0lhrV7s07MHPN
dvcEOICi5MbTXAxMo4++w9zT//OYoq79SPeuA7kT0NcSk4DBlWAJq271VVV2tqNg
kP8TqkoUSzilBKcy7uR+/YHXMnusvhp/B/tcxNjx8Hb36RKF7/EUTHrlRPjdvHXj
TzBBY8Fs887Go5RDKtQxPqtMfiFbAAwUUjCxF+C1GIQbPRKhNuHZzTCTkJ8EBIOp
BIZFV3AT7/DrK2qEFEPq6XhLPOnj3hFDj4tneh3BIXUPI3i4y5HlLapq8PdEYNPy
p8y5uWWz7yR5+FHsP/cLy5gbXeqNN5efJxXmKmZZuH98ov+oLGOwUeQ99Y2UQNUb
Q0y8NmyTQsIP2/txkC2Pa41X5NENzjHT16QbQ05MhY/zBhcTkZ0wEas+gDnupvW1
RWTDHgk01x5PrVx/3v5qJev+63Z5TqD89YFs2rpXbNFCqhKfD6ClvDhAC+9j9ZyX
nzrXBj5tE6eFDQkP587Pt2X++0UtEi/i82FAeAbWv82XnERqcfOBqFzZnxUEO1qI
A3NztEUayTY7qoUAxwMPmgiFQdPEjQy4ohKSqTDFmq9yft+U2rz+b9E+lyxiiUux
UuUWxquChIrVQWywgIIcWAJGxamkpSHY30N3KSa2KrDrgJmg4or20avpmIo9ORlY
iquEMMmNY0NqL2MvgJzMT3V9VaC9PRm26O6n8vAvaShp7uaO5sT7oCOOlQLFposR
CBtSpuwcbOnhaVIrPjxY+yMZ/2R8Etz3tHB7kV8UZjVLFP0/gqkFOCjeVhKcmgSg
UR+L8F7r4nyrqztE3xr8ZuEg3Pw2U7gtfs8kcYcYuEgPnmFbUL5rC0rDz2+YHrLL
CijuVDLh+65C9NvZp7LmIIxJmzFaDsnp7SFdR5TwYrDXHz2XsgKKdGtfU9UcTZZl
+IB9L6MaGIT4vJJc3qDxwFGVCPVTJmpzsEFLvujCaM2qmvuvNYiI9JnNo73oM09A
8yIG7te35b/Fm1LnEOzv2UWYBoLCelwaJ+HTq4eVtgJiVe7b8/W2ubNGaMhkdpHu
+e1q9Xa50iRrzJSRazJRtum+Zcstdv+iLKpryfo5JXBzERJvzRhLgPCi2Llk6faQ
I6KLA5XWOxt+AezDur86Y0nStEZdLGW7jctEZT//gWNfgMOdWhLFxHygQ/8LF4a7
3O6ozrCEtizZpFNVACxxOfMeyRp14gTWAaSfgcmPGMiuASQA9MQb5pWrzDsNv23l
w7Kc3TIPRKbFfMHLIVl2HATQKRibBDGeguBI0hf6NyggZvj11KRzY428xsOD4YCv
amzjrl6axUeMZn90r7DriZxlPlMYd2SaXOQv0oYFheZ257u67R9lSGwhoQ9L2HeX
iOcuKEQAmEar/gjRGNRcGsLezWkFKB6vMavGGbFTAR5reVTt1K+S0MhvPOCQZj0h
B8nsWa2ac5EFnDxNgQuS3G7+TWO5qiCxmZxhjbyriDnFaSyIiF8YuAv3FLxhdVBN
5E+C+IpnkiuaMTV44pkY9PUVuOvnjnGMjQqAIDvk4ieN4OldP2uWiyrrHrhFzkwe
QTQ6+UBtVx5f5V3xJ8yEo3IQS6Bb6BhJZOtKbIOYqzeGZKGIW62Lu1ZT8hRhSNcv
LZFvlrAO9VeJt3T+DnMVueLACutHHegFXpL5nieoX0cG8eLOh/2ObsqY7ZNtSRGW
qmLxZx6+wHcQUUC0GRPM2c45pnLHlQf4kUDSUehPXRqPtmRsHxHlUNhzoGoOuXeL
Ltf2Q3bcXOTRJQJPKPTTIWm29OM9Grp/jwCBHNpSgei+r/qXN0QbnPCHiOPuMGuR
7o2SlSdh+0HKSmsTFrx32f8EDanCkGwWus0rwXZPFFozokoB+xbrvTDftTWXz36B
XqJZz75Zk3Eru3dQsEx+Fwel6LZMVKIwp85m8lUrMD//lMjGNoDiuq2WvZwFyOpb
5EN4XjqfvKvGt43VbsDfCaWpdmYApXfxkMiVMrQIA/SVbacavlJ4UHmMtFfDhZmj
Yoj+0iWK32QgHlKXOSrT1ZN2ib9sp0Uwc/D6pajwzoj5VLUzU96/S+OQudPJuXhB
g6+a4Ml1Vhd3TST9Taa8b7bFZOM1h1cQHw0aIoWBzOPxhco7cG/GZh8DVuUQA2hr
P93sPh8vbsKpuMAjXoAYW1L7QRAld5KcLXWuhakDBh+nw12admNssx3wV1vzfbXS
lIl9fRkr6epTIDvjBJYb6PStpI9ol7nmIZEfroSz3VQ/Z6DEeIQtbct42pGB/p3u
YMT3X4YjBy4vrXJLzi5I87usQgVoXPY4xsbk6dtDUK9mDo4ZP0i0jdhm875o6z0h
lXiFpdo09m0jG9tHFxYC3IH3B7SAR0Tu49tb7aR5EMi6wJKr6q3ox2d1gb2Rg3AN
9jhYVer9dDKe6uuvCSYW547n4UI7EtpBgIEwc25M5Wp6dOW2pWMCZV5JeTqCXk5h
wcfrxnhkeIvmwwbQuiAiLb81q779mi4nLAxyaRPORfAQ8b3UGkuH4cwbA0idnTva
bo0HGp4/nND9rXu2FeDZa3X6WhjTCMAY8ieXzfl5oVQWP/rKTold61QQxkyPtApI
I7Uxg3DI+18Ji+AcygQSDlCUmogzbqAxA+lTlE5wdvMn9Hfl6cg2gVHWVpEAR94Y
o8w6faoZyHKJ2sCa4dmjaO1Oq0Y8MZ6DMEbgNFkApBKDpC6QArmjnmO3FYbMfK7J
ZaKSF+d3xqUMGUGTYHEJ9s9ZceqjOnOlgs/KvOWXkYUjYMHEcuSv0DgFuXvMCoen
eSUXwBi17muCYIP7GtZTzI79r3EM5Y9IW0SSL2byNKDRle4/3PBHflgGNvaKQt+1
+G8mD8zACd1E6Eox5mJtfwlY1xfDEaWr5MEsA1tK3P8YjFa3AwEcjknKFfDafMMU
Yd2P9ZAbMnxNJ7i+zrSGsuKcMIMqcH8zUs3KlZeLiTAN7wzXi2/zWsCIkqqM1OpS
ir1kLeQl2ROvJ/c141HJoRTswhscFNpIlNsVN8jBQxRihTgOIzN9BCQVh+WvufQ2
TVUr7bS7+UFX4XWcpnG4HaEwrAHvQ9flbzr1N5Mo/crHfmipMBC0DDGYG6OBfMUi
6aNsZcfCMjra9OPxniMJ/5Jm9PsAJATF9mQjpIcLQoy28wjO76G3tUHbnsXck0rq
Wx1BiyYCMsmi6zfklIxYR2dlVZuPnq0ekjgwieiFDvWDGC073EURf/MMcnt1BSP3
/9BUNmxsFh3Z4u/Sbc1w03ULnfRlqUk+js78WC6AUdfEWRYrlD/zspvMF8ZsGA0i
m4leBeWO2c5WOBBuipuSfwZWCcizNz6sLJ05H2KfYtdVIFdxvkVIjQgjLnpj4iuY
/nOSTlp2pn//4jYCQ93vQPSkZavdVnnoNb+c9OAoHvO2HCve6ar5+LAh9Az9CeVX
+9tdQsXtjc340Ywh2xPD+akPkizs67TpHFFkYwOzk0poiLZYXyZMsWS6cTaX2WJH
AIup6HBGxGqaYw3ijhDjqfHLERxFjnsP8RZhoN2cJf5EwrQa9l4LS9QQCcakp8Hp
f2T6dq1YHr3/M1xtD0gnfqmRh58T8rywCj/axVo4RjGFOpWqeGou873qVncgVdOb
RLTCzafYfh4mmvhUfdtl15r/OPb3c/eyfqO8gyScIRHF9Z8q47JXfOZxwnyOTe37
yndyfFY8/Uk6MvvxyygtSj4TpoulmJtXjs0yM2ebutqlFTdkLhWLEiFohmlYY93j
O9E/ygHfR3RZDPcsX9VeqBsCp5rE4Q36GFyJs5N8l2R4JcXgjQz0XW9VoqmcCMjv
eN9F7rsduv7gaukoYMyLeIx9H4lLUNkkW7OhRB27Sdgl+B/LdIuSYsmv9YY/33eg
nzVnjRMBRMJal96hKj591yhvJrJiUceJaFbekbc4mEr8/EdvwPU2x3Z9VLURPlhL
D917MFnfpNkan8ti6tLR62MviH003m6WmexYfuntSsG73GrsIdWTvWk0OMIdeDzQ
GSrfxfzkdc/x+O2pvIMWKkLxfQXg3gMIid7ck8UHMq1b4fOQAdz6lW6uz5826mnQ
7xE2SFnPKLR/uB4Uu7MaKvygdP+jxzMoQuf7+0NJofz/dk7hyBS75UvQsMGc2Wa6
nSqd3tXK8Amq26O//mK5JJmdUc4SSTadWx5rA0jG3YAPc9QftfBD3ft4c0za+gGD
cpQAVTZwQTqnz0EFuuGc/dmTn5NVQFmEGwGAAr1yJp5cmyRMmHoeq8suULrChpm7
5yQ0Hpj1mwZXlSRGsU4Y5C5363Vx4WlDohVgGcpWz5DYF2UaITv0wEub+rmTmxTp
4GO0u+2Y0cZ10bedzw4CaMec9GSkaTpAYXQWOHlWwjrMM+AFyL+WULgRX+Q5iomQ
1EpImku8T5cG08pv+Xa4NVPPVQXwdGSSZhsVXAbtgSvGw0p2cCYbjwYnYcoNxAii
N/RN93L34cVvst5XXFhtmP/YYxZNA2z8Xv2Br4zrya238ukEzZTSR3hnr9SzCYAt
r7lInewnpRYSrkmkyHX3NZWkxVIZ0Skic2+SInzKn59s5ohXDdi2g4ARE/5AwuLf
UHrcZwU6wCD3H95ziseWSc27t6DQ7Fpq/42yLMihhQnLTTZyoyMhlwI6g1Qln0Pg
DipPjhiLB6tqM4W/8lejboThsODH4eOGJzAQ1gYyrzmyv1l1ZPMZuhUE9BIGmH7I
SCbkcxFXFYAAKtAHP4fioqAfIRmOz2hTOhhxiK9Ol7WW/oV6XFOn2isM+m7qCk/z
cqP7HDAVB2tOwC99KB7UPNmttfkEfFnDzK346UotDkQhhKzVIeNJpv55Vct/7rhE
CU1KPYCIuw+/85vcY79/m8bDlhNGBa7PAJQHv6BmUF2oEkSUPIzhPBJUoKj3kv7l
3x+0W86fqbrbjeXpPN5H/sbAwDRNrG73K5lHmGPQz2zfCc5IQHipzDBz60zmle+w
GrxmU3yKv6ZEdv6ZOu3mygO/0KNGtVZqQCpY+cLN3nQ9/LuJY/f818QrDvUa33WJ
mR34TnfgXHfYaalt5CHKlzaCYthVn1YyypePlWanVh2cd7NitZQtc9rNvNNohkzf
BI4DIQFgQoIeng+3guuDOmBjLP2MtozRtaOn5sthcFwayCekJ0fBJX16JCyrBHfD
MdkKg7BbjL0iijpcNuTZ08Ls5AEGPKIhCxsnz5d/iH9qMhOLWpQiHYtDleszLZYk
5gJt6bJyGcN/mF7sl1wj413YBkA2ah9PGNAj0ljKHAACmm41JlsEOc+3YbFfzfiB
E0nvJzKcw0PraYcwV8cX2lGlYRD3ThAGqA2Wl51QsYQazlU2VyXXqI/9m0BPbu3o
XtdncnrP0xUT9UN6O1fBVfnSkWjYsFlUKAQTn2P/uiPae3lRNiLVW/PFvVpSvw3F
y4dufDp/Nq/0btvAUjomxeGOUCPkUaOuHha1Juswv++4TKV3aRfUxrIw1WT3aq9H
d2cxQ49IB3gL/sqmyUYLwX164VyiL4OrIyojEXcTJx5Nmqya0nnewrluNdxz4uwD
SK+OKw8Nuw2GLEUrCOvIHElTxhBv1MXDshaSxGssIQG/srz0Om6a12iYH+IHOsJ7
nkYLjt+OatUlr2opjpvX03LM3aXbR2zkZNQuJr+C5mXovdZsg9+zxBl+4oIYqwK9
3xHGWUIq74eOWtAqzDMR+F6hlIJ6StXaKXj78AtXSNkf/0oGdnh/AaI67fZ+vexf
jv+8JnAtcsTN8O/9+f+NJVAnwmr5dedebWpeoM18ebNXt88Q5phgkViYmwAQ9xde
XUu4vlSN/mBoxvsI+a8grAVNYvsNCl5r+R3GmZ2dhqL6052BnYxALxcTNNY24RqD
x5D6QerKW1hVjZYiDqhgDD5N1xz76hNbmc0hUbX1r5AWhEodk/X9lKj4ru4mFgSI
iqrq/gYmqu27Ygyd1MuZNC6AV9yjW+kykBGFlEanmSd5suOalUadcdyZsyRO4NvK
qJmpstzGW7I6AN3QIsVNT+8oTQ/Hl8BStxd04IlUApX0hOvkIkTtk9PTKI2v13sy
bDOMLL7cTUQYBWiLONfvH6wHlHWHUTdN25oZoYz+U9BqZqDKeomT2UbYNExX+f79
1cvLDa9cUONXSCOkel7nTb/a8O+SpYFf4N9osaKU5u84Nkw1aZAyQAv3KAk4xAj2
XfTkbxgql8LFWoYSD19fzT85jq37ZvbH0Z78jis/Hr7LVNgNjyDysoZ46EXTHjFT
AsxSWAct0kbvO/UZHjZxuCkxhPCUSXfKtepuOFRbo0kkoHqyi2DZ7bUJHI6C6Jir
ss78Q7a45CKSSRVgjxkSsUH/8trPjNyUhj0AEh0bApQ4p6QNPWQoaqt0JtK+O/fL
mG0RTmqYWDxbJeUU/ZL9d7BSFZCfrePtyCs/TDOGNNqMJVkrVRUjJSGBQrINL7fP
2U0oi3N+rn5c01bZ0LwJtw0GMBVC46vaEjI+h6ytcg7NqS4r2Tas6pMlHyU9Aocn
/TG5gL0kQ9Ja9sFddRoQAUhqTh6bA73VAmEBnB79pMhbSl1YzOaP3Qn07U5ciVGC
hwmhd9YuoRCYjh8fjW6i3HZ/zsVZZUjASJ0e1vlKr4s4HVnII4hpF+8VQ8FdPvs8
jW+hZ4Ut7k9sBI0DQ4EBc0vYPsXN9jXjliLoWO09+gMLV8oD+7LgYAJRzp5w9bHQ
B19EcAaZwrnQ8CFRFM2Im/Uj/iY6ef1FVe812/QKO58OJnsrejnIAr+/4LaRC4AK
BIKs7BTTfpX7BoDDimOd7GncQTYlHxU5QkcVM6qXq9eXQfbSvHNYJzS/GrhGOg8c
6s3U5ly0H8wxnAdFp461KgHVr2FyqvKEd16E7bccftq5l5hXeIxej/EgFrB6QlY9
hBwQyzVsSMp8/k9jJqxPZ2DU1YPfMaxaFc2t7a5ZPNw3uxbGH13kojnbMgzXiDSC
VmBnxrElNtyDhQhs3dY4XiIuIyAh131RP5XUmhD4ia0uFuCpW9Rs/Njxq/kpE/rG
vJ6fICNjYdbmyVLCNLGcoyRcgmrw6gd+UC0JOTnk/gIyTsdGG3UV9BJ6lFM0hqyl
tJqJBj755hWt5xRyTKreBM2Z/Og3Jut9VCL4Z/aDJqGm7npzAXyusOxKcaWzEsiC
3fyBCW2DJW08MTikJ6ho5WUN8zs2l9ZKmMs6DVVTUgNhBzTc/l86kBzaSsFeTPRY
aGIN08wNwtoLx1EroN/0OWMYCdbm9ne1aCBy6J+vvoeLUlq3ZjZztKin3xH6KWxp
kiN0jt82dqaz0f63I+IhLTZmF0e8p3FcL8er1xQW+jXl3ksJgUr16aHG1wy5yf+p
xcUzv41EdmgcnBqeQS8WsRzFjSesw+MTi9yxlPg0/UbsNZodT842c78RMVXWY62P
oLNjkLC9PkO+NTgQqf/u+rBtonb3X+0xbzy8igSZV4mnzoFMxxDiAfKYmf7uA1KA
rPwB+rVrIGXzVjdJ26clZansDxySiBAWWrGcEado7UPJIpT/MH/qPtHqWXOlT8IT
+96s7BMQnWuL3+3lwy9jo5c/WkQ2l6EtScCidm5KA5TN/8VOE5CwWDgu72E0GpaD
cmXhODgRsvheumGStQag2czelltCabryGck1xQ4OIaYvUMljqFUwjzEr4v7exdfA
BoBUK5T44RRwzZlFMD/1jaop+eZ3fNFI+GT5gQ2f96/Uv3q/nemrETtncLiaoDAy
Bp8ZbfCRI90SgjZN/kTXfvJLH2ncOpyDz7juyipU9jscdY6XM5jM7T8sMVv+4kqD
uF9AHzkE9pQ03QMQDXKJbuDUtP49rv5z9nMDDUrwxh9ghNuyeJenU55QddKeuFJl
YEOC5RCVig4a8JC8jrsDpfV/laauFg/UjQg1mqdDdmz1pkqQJA9UYqMyL6T3UvAY
rk+gwWhy1T02w1O8rvyza55et48hIiDgiIQiLnWH5cx9LUZ+dXV62nvJ+N+ulsEQ
s7VjM0HJwWx9msznbC9VuhG9g6g7hjbrlkE4oxzcyF+MjTSQnBKM306qVqc20UXC
vn9vnRfzSfzXRUlspAUOVMBB5IlYhsYbEZiby4IJiH1zcrgbZmgD2AM1sVFoX2fQ
XXHCz0vLqc6laoi7oMTbdSmxmdRTtPiIwYidcGX8SsqiRxyjoe3cmYqS8W/Hd4kE
95/K1zs4xXyE7T8cQKc9j1cQeLRuCNwPfBduKFAHkPs9odo4hckpXn6koy5p6iC9
fxmaAXr9rSgOSPyMUTeBdCdYlUq+BSuz82vTgAiNAcOcqS3L38QamKJvcQcHFJ6f
UsIoWiVy8lWdjZsXOffemK/UYhNjuDVXcxx9vVYuDQkPrqw/pOqqpDEh/hvPCVKo
TARRHcsdvDbU6B7YaFrpnOFZA8ldz/F6by7CscuoZ4PFASJY6z2pgkkNr91YTW2Z
nqfOhxWjycdaM0Mvl9HatYYQSr9fdYrmM1UoRd+u2n0DKWQaz5dLHxJHtYqld7YA
0tUVsrT3ID+WGmWgVikCgVHb3YjTNw0mXvgIxITLhZm1/RKlANIMRWjjilw04j94
awUUxFwg3SVsRozMsFMVOw3O2z0VrNcJeRe5pprQCOiWcCOYMKqWtiSNI/YQXW7i
GDZzqOadGe8ufh1AP+TpykgonpPGq35ISV7sYd6P+k71oDNrhd5y2Xqibfxp0OPm
nHGuxKnmKGFyWNTJgCAjuA8pACi8z5FlSU2cirfZwiG5heJB20bE5uen+H/dUbS6
rAHtGMDoaQaNCmteq2KGR1cvG7sIHMo3CTrs5GdxGfM93UTpBPvq+YkSH6OKwyXD
smFqduVvxogcoC9xd7WCpdukrd3e9H/xB8qZiiynh/MdKf8MbjwZnCO28Nm9rgWZ
G5S7gsQCjLsutux315XIjrcMXLQC7KCiuQLXc5DXQZGs55VkIbt29187RLlYmZTR
zMLfk9HlHa+R6QoMLwK8ypDpgrOXi17CKafce5RuhgTOVG9aWaobY86jEnlca2dR
MdFs3PThR71/j/dFYAzgxTpWOJkwbrqnD11rU3wZOVTJ+jcAJWUq8XI/tY5War6Y
sUJXS5R/HYo2mkL249qobz2ZWr5c6OZe0p/GuKBArSDxyw84HGWDhuENzv/0w8Dr
6uFirmHPw38jWwmM6NrilTWsaimxi+zYplnwJhm3P/b3JlXD0PqyL8tRwgEd7gTD
FWED44DED9Y6gstnGQi+MzInu0wEaXmzuAJHJ/c0daLsdJBR5DQymsj0Khef3GzU
gMbB/HObS42oY+zsHFarzRo+laByal7fiotjR2/mZhNhkQ+XeJdzyKmX6C+Cb+qL
PCBwEY7Z+aj3+jLfe+QhggHW1HKqOlbugElOL0pMN8rTAa9Csl2d3KEFxzQGVJN9
hfbeIaXUXxRot3BiThR4duARcQqQPqd+DbLBczaSWnN3mYT/5sWzjKOiO6adgyUo
d8+on+xnZz1RVDtCMzRgRiZmvWu1GjN/lC6IE4Va1v2CAXU50HXydhnKrYqdjLWx
pRbu9Z2yadbogzjHeO2V2jDFggyuwUEFEjwaBy2cGG8/+4wTEJVz7Z3V4j2U+py/
7ZXhuv83sKnXLOhfdYrCRUISCzFSze+n4jmHkhQRubJlIKnUCrpJStXKML0w2yzw
VUJs2PeAzC7bThc2G+WZ7fja/oqOJxo5PZ8RK2kyX82UWiQ+G3KBjs2mEC6x05VA
GMAkyHya8CrD8zfr/1tQdCiIumX3DGOUj+v1rS8HKhGOSY6gWeVNqz3GpoOb4zg3
NOW71R1Kp1iXC6Ub2aWsHb92aai3pwRPu6sXwE/qt1gscIEayemB+xueXUCCb4HP
8OuB0nDvgE4kB8B5zWvAvHW4dG+xeO8aJfKTTBwRm/aqGd4IIEDcYALYDq5OZA/8
iLKBI2By4I8lj5kRA05GvVSxeKa5FGa9N5rVq9UFDYJPKNxvSS97vWIyuAUvjdqt
6b+X3A8PxKGnsyAvbCZd+2psTkWEcEjD4Jcp5tIBqVOFEKCPOS12h3lhezjdB9mq
+XKGKUkI9eSGJC+ulHMJq6DCxbnKUxmMeE6+jPdv77JzBxOEwJCc9AuOVLC6ptdf
Q71K2Iuly8d5eagVLO1sS0hz4IFCsM/vL2bapHimL7jKId8TgjnSZrxJ4WOYfBXC
YGVZjtvRxe4MxyOsDZtZhb4DpcH2UjzcW3h3rAMbqZ/0tgTK0LCyTbZcbvKYUbXE
wrjgKZzowAD1VqNcUC4HDXpbD+BikR64sx2JLHvFDhL7+sgH4Py9qCT33TKaX7Fj
xogkpMsz0YXz+Yo1bbtqVtofZhhF7MZA3qunTZxGC4cXV5D4g1fttLjOhM3Dz0MI
Ug3N1YyuYPk8anJoflhZ4/yakN9J1i0J3+GPG0iYlDe8J3c9rsFKTYn8m81UpqCl
CRPITGVXEDRYLZUYu8JMK+9fOKfPTm4b7em8p9oGsAnLsgncdNLH/0vxJf9hqpX6
lpOF2j5cWkHzMBMo6/OvdKAf9scjixE03W2DFNKUvBTBcXmJlWK2ar6Wi5mEpjDu
tQG3iAbBRMEyh1GywfLdjx9N7HsVtwiFD4xGjl3eep/SKa/05JqLb3uKQtQ8XDul
0oA1zsVbA8umnxTsD8cVyMWAHh7lB41lye5Rg1bQ1Ovf1ECw/uXF0NmuOLFRsja6
a82tJQJKGhoLl6U1+NY/NkhqBBkBmWEywLjNcCC4+lIeVB3XXdd5taVIXJkK4SFy
Xe+1Wx/zwSj2aemFSkoJUp5lowH4UGQBRzz+lidPG92iv1SHuGIVLFzqmoJqJuEB
j5CtZFgCp7D4AFcjdNklnKLFvnT3oqVKp4MBoL/WJiMtoVA8tnj6zU5l/nLMJ7Pg
2vDPjTZI4hgR/ElLLgOhW8o8SCB5QZYWdzJ94FaZ8xWU1Wo3smBXTDZaHuPB4NtW
PDnMqF8NML34QxCNXwOfPY8nPnJk3EyXYT8f32zMVXbNpGtSo/620PnbtpTY4jjd
Rfj/3golmWwhnkEJZdED4k4UMQ3T6zPmtW8JWt60Fr3oPh7amCoosNp6yRtNbmTO
gstasgWo7NIjZNZmhNd3RhpP4rCpK1NmfONY4TXYir9I7NTDCWcWJ9eu2KIF6aVw
SHq1/NaRF7O6hs51jLasDWZ5zA7SB6SBegUyS9YGC9Hu9WQFBNI8X11I4oDzl01j
ixUOxkJN5HPGLymyKKAzPn5zskyaT22HXsV7GDCbhP6h+HXm8QJJL24C+5whAwlB
6WD5MW5tUJcegYgFc+AKbRywcsFgw7XiucqsNugsMJhoUsWg/lCLaY+dm9KbOp5X
/3Qga6zwTtwCgosDCDTxeU79yzOYRY9Bs3EQDBu2W0Q6K55/hl7Z4oN3XUZG5utN
VjaELIkn5FiN4O8iPreNOj0WDDr703bmLGs6gquZo91elXcWrkjws9g1j7R/UOrR
4KP+oQkIjDK8fWgiDAVcNqZc9AIm/he4U8AT8mgrYeotgfKAXNPkXKuBKqYLLbIt
OvGps5+fb0cx5t2ci1Ika9DVmRthZPjGuc0mouOfex5QAhfLW9jU5x3RKgb1XHxe
a+m605z0SsRHFO+6sf5HX7LiF74eZrliQRStxHJ7RkUpygWUbp6U2GQeKuLutCd6
48mDAEjcpLpQlOtzTVaUW6Ypf1xVqZlY0mvz1/a0beSe0BoxxgyXjoZWixbgh0ld
wizlmBLUlTrO7dzI86UrmQ9mKEEBCbNiGUwaSNAsxU3b0uUk4iVhK7tzNcEb7Y/i
iStW9Iyxgw9BqKJN4jXQFIJAOPZsSOWEB7ZY5Vy3kSmAXLNfqW5Gc8KYoM4RsuZP
BBFdJy2Ky69Br8aCxg5koXpgAc1rBojL3LDF5kVHKyMjrsmS3b7PRqg3Z5bpb1zK
qkCELMzs4FLVeBJE5Bq48VwkOguambAiMRXJQVfR+UfVtYjfnFu2QdJAHqF6UlXh
zRuc7fP1uavf+N0FFrOioUQdHVOO1Ae6AmXQGCl5TYaabulcrUGMJWG7HH9wp8e7
l2+yunTNl0tqyOXFZpX5WZQoNOh2zRJQi4Q99flS7Hpoiz0HzMf09DBGIy8X/2kR
xuuwLMZop6H5gpcRVeq9ucxs5+vEOAO90iAqeN59i3B59Adz2Ds6DibvSRM8pxO/
RzeFKzKzolICfJQFwLoPRD0e0Lan8xakOCdi9ry9RPZlZ3yW6izFG7cLYPdj1B5s
adFV3lco4THe3/KOLCH8sedmuEl83LrScZZ0F1RQyIWZkQRDmuOGVwghzGkyHSDb
lu8TOMNVoR6onhfzaTxlFFwwiiCr6fQvwEBRxHxEo4QEMwS0R0L3pMA7IUJ9cx9+
r+32WvmUB7Xceg65cCwgMd5mXk7nuAhc3AhpuDrJisYuNYWl0RM5U8Yh6EI5FFCp
1E9IcB8fxr02lGonyQmwYNCo3iGt8M1BU8f45y5Bh9/vce4hgLQrFSk0kDONvqv6
SvbVQd2je0N2v9DlXrrE4J6dzoHvUjdac/CVDL2l729NwkxpPbXoQXooL6iPw/4f
iZXFRv1mJMCu5oi+cuxRmdzjFvWKyMRY70HWZJ1KsS2YngGISxV70USuh0TZfRfl
S2SHQ+q+iIUueKINcgNDi5Plm3wDrl4ndoFY4lmG1EEycq2O3gUh/0X4Rc6ZUXwi
qANeMU/Ma/1Rf+dVUXJj6FBYKNLoWU+FHTuW0uJ4nfI/yhQl1xOyfaqNutG/3iyd
Xodfxl4wWdgD1s3QxI+xHlZpOhrJvp7pmEp/sTfm3PuFulVzqHrLbO4blvxeoTxI
2BEW2/If4+Vw+Eiqv7oC8UyXCPeUdWIRHf4FZ3c+gv8JVVq/XD3rT0/GfagCch8S
BnX/k1ctJpxb7lJ2M7+2BHIB+eQPhEDCiMrY09UBZ79Y5jGp4Nt8yOC+4tShoxlP
2OeieFmzaou1mK4rE1WXgWI5hbNX1gD4GaIokvKLg6i6TYAFiOy1drL307IdY5qc
3r04m+uqCbEu70wFVGtSeYJ0WKF3YbPJCgYcN0PXPcDHVQp9zPACjN1GuprvHOh/
kRg7yQ5Z9b/6COQXKmiSe9ixTdVNKBh9z/M4qEwqVzS/nDmtuHHUcEoWpzuUZ9ZO
MHAuUcnIAN0NSW/KkyYxZ3wI016l9S4YdNsZl5+RhzrGgKoKlHR3XpMUhHGW+5yl
cELKlkn5XnmaQ9OEaclYiJVm40YBCtUeT4AGSLcI5i/1T65atMTHH67o4JOB0Me8
uxMX2QKTwO+30unogVF2dEcySp7OdHHKkzZc9vEEy9Dq58IhNIwrP1C68CLUiMdt
azYL+aAxaflW4Ec/6OQlBVBM187Z+f0Mff0YKuyUvpR1SP1ODOGkWrZxH4iQ+E21
ZXuH9rTtTSBa6vRsVBQijSPkZYSlarsRJovo72xMwqGmL7fq4CZzPm2MA7GPaemw
eIY20+2uFBc2uKbP6DxE9D+LMF5HxPnK7uHPKGu8XnoCxvcY3Td+Ot5Px1gDv11Q
j6lLuz5IDDcxJFwOflis/d+v0XKYMhLFhs4mGNHzbwmU5jSAHDyMMBZhJh58Aw6c
HbLHwf05DihwZEMyG15uZJn7jBBnaHRh8HKpakPean3StXpz+hdu+cV70tPeQaT9
rS0kMKw0tjD0UlKs4jk/C0YP1J95U8UQy2MscJfaaJS/9TlvcE+q2QbkmCWiMx1h
K8iCl2+uVr6Re1MF7AvtNZjXrIkTW6yWdASvQ3/c+KtQJJ/jncmW2er9LiBr2KhG
wpXgYKBLdlbn8yDremNe9osSOw6mL1gjeUjKhTt+phvPipfHYCJJo/hml7luBQp8
JNbk6QRcbLE25wdSW0kWnKzvk6A40u6QHyij4lFq5RMuP4kToXKAon7i+doCUykp
CX5/OoPAsKfip3vjQjYoP74OqpwMoK6mtQXtaGMiaKcAj2EI6npLSL97eVpSCHpr
FExtvVSU7aJFSFOHEqY8Li8r/o9MpGvaFqmijt0tVfNRBe6zEHZULihPRYGpG0Ee
XWBqNqtCgY4xF+ya+T5s+w2uLm40NckurfSuk0Rn6rRCLo4G+HlYwomOPjtPaJ0B
Sz0ZpgBXP3PG8jOrS8QfpEIAUgAxU6jWTLKRz/gnYpWzn/N/rJlDMszpYpTalk+W
eH+hwXNF1WMn2lLjP1hVlKEM4qsYsSEjrvcl0g2gtc6asPk1PFewKTWcFo0x3H04
A1f4fhC4zIkdE5XGk62AWHlcZFwHFgDpb4+ToL6mU+PEg9MEpwTtpQ3WHU4TBhdY
u/5HLRe+poYxie4GMa59DrCC+fGzE7IniLmehkjj4B6J666wAufOTSKiuXl16iXs
jzdTxCe22NUuPEBKO/7nNEJKMxYSIquDEaA+vYCNR6Bhrcq7Kt8v8kmuYsGcW6S0
SCc8qqwoh/t2NqFqVPKUkuiCjCwfB9n4xDzHSn+rtW8+h0tDTlx/pFR7LxlbJxp9
yk7RXc3uYGNSgIhnxxMIGEo31NO6hPlItArRia+DeLxDBvxkUmdJ168S5CB7aMUx
BnvUysC1AaanFqpiUCmtJphHkKf6b8xRceSXcGHZwQ2Hm2PgRHf3ONpmKotKXiqe
ubNYjluVsLbRD+o8cgaPk7AmmglpA5T7aEu1a2TViXChQrUAHvlbf/HdByMcqZUT
sFo1nmznbmeh6pdO76tN7kFAamJQdAZS856gbaqTjjQOqrzsJ+YdE4TwrBVRlB/4
24Ey4UZXDrFBC6mjyT0iWjG9k2lb2ooyO85vZkZadAXgLzWXWJh2aU1KeZppoCfx
tg2c/CsV4gO4gHxwrq9G87P2ukSL8KIao89E9cCkoL+EBaWkri8zZNiit9xp2hLK
+gndDV4O+5xRMCUYKCBoo4vhh95/Rlu2Lkq/B3gemDC0ON0Xp7naR/7yzFSLYmo4
eyF2aq0E6DveJ3/r8L6VBqt0HRHsxpZNpbl5Xlu4zaBok5vH/m24uCoSwDytwcHe
ORmMnpCLkwobqt+RXSfBssjXbx7Ni8UYp7xqlm5ODvfD+nFMA8Yz5ecAmSo9SeBg
aEXYg+WSgNQyi0AqoWV4lzBPs2KiJKwRe6L3dWxle3VpAR/4PBIgzFQ67iVUqOqo
TIFP7e1WxU8XsVeYHXnoQFVbWzSHXa3EKxta6YQqT9a/CYm4Dy9+xkqzd9Gnxe0S
BedFZBBTChfPMmCvL4BotqmXxZIWHkdWg7/bI3EvVB5q6FWWvr7p1bFhAWGuOUqb
mpw0i/Sc83D2f2zqtVjdaRVjsxIwj38lWVhf9UwjAHjBYKT0GyzEX6VoUQDI4eBM
Cy2G0EUGSEjs8+0D6QPhr8Jyu4X/iGRIgYW5NzAIU+MJH1wsNpXmBDrVij7U/wgs
jg5gg/uwO7n2hySMD85qx57AqFT7txkdC5boiNjb4WXOPpDFQuaAhxjDJFzKl5tr
TEfZZ+Xr8yE/CgHY/zj7t5694oEVTQKHknXVGus6lSTm+gfrki67DqG+cvknAY51
J/Jah1SAtEqUfXOzJDbKDwtP8DidBCqICkRL50QnFNv4BdL6ziWyEy2WllmQJjy2
PVD6v2l9HpiTIUmlhq6/ZLQrNk/r5xKhRAZLx1nBHF3sGM94HjsWwn+IQjQjNUmy
29JEIdYOTEL9Vnvvwqnqlbrapa6XLUSDh5qXmnsRKuOYLXaciRn96k9jgLjjN559
E9PkJ4sxYsOYqCxjTMCgHf8i8Ho3YV09XN9H00mDAjxlc5QMC+RY5crKNQ1lqvZs
Kteuk4494iMaEV9klNTNjRpBfHcL+4Ue/X0DBxKyZrRyseuD6JD0Stouiw4t9q0+
CFTW1JJSOSpU5xdJtpfpAf3nUxd34pUW8wPYjRD18cHQKeoPdEpn2UzKHoN8BpPp
h0NzBoEzHr+kQIkLhiUXafbO04whJNW/2zRtYh0cyImyAUTZfX49OZi8bVJTYRsf
CsEQwbaDFoP0+UVsZKTpu3fHYXq/wmJCzYQeBE51EtEcX9ZtZGZzHVKndz6ZE53l
rR87EMQaqSRGWKzh/QSf4oUyj4ezeFx4UMBF7RKTTe6ydwlaIm2Zkh/+L+AdvWr8
nx6luaaLoean4w+MrOf1HE6q2+SLkOJdbRtTWqmjy3v8+QDZFZtJ4bcz1AB24JDh
YEuReScOljp9bbsbhgCkHQLSRMwcDMDeoaTk9CJ0PPXK47R25Qmi2CFF2zROTXX6
injpSEKtrG7R9VQndNElx5stG+NAGvsqjKk8RjGBvzkzoTa37UMLUl8+n2NHdeVq
+HiAwMZw4xnh/oxjbimPdybNlAwVskMH5g/fZqAwMqnorLZhtct39rEY+O9bqIno
+Ah+hUi9JcGBqungswYV/Tv7IQHuOqLY9B0kyxHTOgr3l+RDLGXSZMRmLd+n6P5H
o9BE70WniplBmGSZx+a8elnC+xIWZPpxym/PYHEkOjPnF2zT5anow9geVzsM22Dj
TBYvxg+BVlxUvZ6b8iUGevdA4hGoOyiQ7vyK5MpJllvdhX8XQc9vXcoCWHif1tYA
SVzauTd+to9wZPBY/SsnmvwTHOcpxhSRhphbPJMN6gljIYSnNYu36/mVyCeEDg7w
Z43VXD7IK1HVJGD6UVKguWQQyMY0Mmcfhc2xW6eXMybW/ux6h2prMmTYxMICQeZA
ea//aUqAiz2sBO6YcB/RNI877bxCopa/WBj+0S6rp6s7vYz5LGAqw2FjVBGYieiW
6ZRoRIwjdVSINgcriXJCZKUICkQjAIVtKgNJn5qbNCdCkBhDB1Hf8Re6KvA0g+hx
nJPq4xpZ40l0fh/JCJb4mjzi/LuFhXjHVqCFZGWYLXi2B/gO7CoVwuXX4BA6WQAa
6nbAf6P79FmSMv4fHky1Nm5Bi0w+1oZuKYj6O/UucPOZpRYyeb3ZvtBZIlmzIkpD
wOHM/ZIGf9HbW8G8rzu8ChlvVC/IW24GNVdMHSLpWEeS6ataFsAcdwzFDAQB/E6c
tJ4ApK19lSSfCw3Cx8UItiXmR1wmGh+3RwaYO7Iq801Cr2cMN7ZBrf3JNJusy/Hl
K0286eNNyF4VBLiwE2D24P3HysjAJQLG5glGoutGlgRyaGtSBQaxwVsP4hClkJHr
1TrGqTE1frS8dR8Qo1OTyn6l141VE4K6N6u5KVY7TE7Y5FJ+9OFkBgYHzHLbocCp
AuxKF3GXmOErHs9BuxE9QjFygB/bG4Y++7I0HZ7Kp6JBfjdnmN8UkRuSjtFSE7xf
FaSS0SrmxD7pE1J9aSzd2h9MPtlwUM0am3f1K/UgjccAqtP8BOfsZ8ONfapTaiqw
dJQ6v4J7n2PzuZEuNNiX27wfi7b++LraRFwnAEQQW91Ad8S3m0+EgBpOnajgouBs
FvCYVMDd1hYrNT5tfyf014PPAEVv7Rk54UL4wrZ+fR1Y42cxE7gJefyBNnhenFJF
lkhgwwVJxVxn8EuW7HAl5g7vs/Dvr8O0FJfENiQcXci9I2LrSvSy78Ciwpl0Y0+7
zh/SZIPKYiv4TchnlXVpk74M5Undqr1+5a6iM8Evmf0reA/gEIcKTOIY36RezvMe
zpa+LqgRTnyaS2/181K09HQnzbZXo6lU/tLxcE1LQ2Y9C4Dt4waoHSsis6Or6U6y
DKKeGoG0dpyzu4z+I4lFi+Xg5hOVB/U0s1DR+8CpxRuXgbSxoTZMmM6/bC2tBvUH
7+96SrnlNXxeNXDAr0wvUe9o1OVaExzkmgp6eRfzTYyxUsfmdiXs3NVYVoZFnxQw
q6t5FqSD4qSk2kNBqX8sA88oCJBclTC5qKrHLmcsoo/sMAfcpC5mtRoQ1TxHJiJT
DbYNU17VA7a2K56A7fcBrdOTTQA47LwJgFdaSAdOYK1/4EX6839/lWV2qA6w+XE8
9oHvwu/f4VEF8gyPHaos2uwiilUvrsm+SmDhoCqVzEu+ddOkahCPCjFKaEkLdVt9
dSfcR4UZpIJtQNC3fN8Ae/WA0M0MNVHT8uwI3q0Bfdi0IZD0o8OZTyz9jQwJRdAb
6CT3yDm3uTK2fdxUFlfupzaUqqJAYQgVGaAP39vQiSZD0mZ2jqieTmG1j8E9ziu4
CNPNnIsoR5FMe85bUsGcOhM+m/gvE8ibXQZfNM3qLEsQTpceiSiIYG9r9ahgyA00
L0Oj3jfcKQ507FJnrEHszv+sHneQqcZu1MVImkNiqgIJe6NK9OqHQYoj2xIaQxdN
3m+bfEb2D6e0lPvM7CJ2HhKFhzKxnm4dqRKxreymBXJ2jAxB0Lpyyk/gp+J/cz4M
Zp4cka3xWRjTCXHsBB9LrFfeLnSqQpa3hMoMhGL4vEu/qEgMcL7fFMJJBqL6/Lm7
hxvLipExXS2DcSOIM0jIlRuR9ZG03KDWdQFSIjXmfZnbu0aECfCrVyXrE3Jh6szd
QJ+S3XBAdBXFfIgwv6/Rgt7fUcAmdrVjF2LIyk7gZdC4+MoGJE9c0BqJyxzVpvHY
UB+n8ro1yCMgsYsmdU0MCbufPKNHN5YUOyzO5uId+oMBwAQ5w2ZHHJ5DN1aX3g2H
gKasAM3UNVKmYSzsbRJpbCBEGYcyV0QZgB4ECQRTfl/GrQDOvGF9pvbxWTo+/FHn
Gchh73wrg/gFagoc7zeOx4wHyHxhZZTwH64FCGc7bUVrhGxjOqxhqYqZEB1G/8sd
MmgkiaRh7fxPwBhoWD9o4lXDXLbGjTJeqjRxmDdjgxCjpbA2jsT/W1Ee5rLjBerj
dpL6Fjf8TMW2ktKPjgGGtov7ha3vE3TY5sPJLMGQHVcVC0UACPIX5r+vdkHRDgFF
faTD/3X+87Tr3zid97ZnnFiA9n+/G56oUJeJuvnAU06nMC6PtGzenQ9yFo1lRN/C
TycvhJcpEJpe3RFoTE5xSa2huijRw60FoKJlBDZf2nLjPP7VRY/8aCt7LgOAwxor
n568//PSm1aKo4ExknGJCGCWCzqyINB6o3+nIg8fFmkE9XtQTDtDTzW8gbN4IVTz
p1+D4OnFtp1oGC30DpnyvkatM8e96Z2v1Mb78QXFK55LOBvkZjiFmI3ilcYaoeyW
Xv69za+wq4pD7nHCP2ZVJLu2MjPG3A9WdtkW24vz5V9OAt1I8y2DK5NrjC5sRzaM
Sw+Wk+2yhyBVTiq1uqyGh/PK6Wv7aJlAWqR8aDlFjVlAfv2+n3mIuPuAUX63aceu
QN7hH200c9cYtg6oreRE9uz3KrGUXT6vdKE6UDYT6ItBGiv+245B4voUXPpHkcGA
mWiGsO4m4EAuEuCxXhjn6Gi7yVGph2YZg3JzaYqber8srkNjZeGPaPw+LJz4vnN2
pZwo7cYeHlQ1spEibRHNw8Q99/u2mSd5z0WS1oqJFfIAW2aEkOAj2ib1UJCVpGDX
L6kz2vygRTs8tn+vnbjHS2wurHUUt1m75DdrLhUUEL5zZaCW6KgtMbXTyaDjPNSl
1QaoLKY5fbguWY8NXu+5a4DzQu+Z6kkGQSVnHBLqstHRBeSfTpGZKiMmj2dugnHW
Inn9Bpm0pKWbpmngXXENQZ2G99HfT044A3pLWpfV50Oi+MymcXB53zxzrYec3tAa
8y8C58d7L0hhBaLqCajriuINtiPb0np8viFn2S89EsP2oAcUoiOVW2/mbaTcbwej
sJTkuFe/LSBnLXZCu05tQl46a9LXAbvAjhYKNqBPmSwTNiOSehIX5SSYK2ilE0vr
43nI/Yu7GUcwvpNT6ICGWVZgePb36cR5tR8crXHZqiLWuNZ/j11HpBOMWPosMa+W
Y+95M6QKHB7LeoxfNfgAI7GhqBKQFHh11c2EddCuUnU5Ci4bfwX2cGWIi4+/PNSI
asVaJvIuuxrDuKfn5LEjft+vwlL2PdSpG9hDp7Qu/jmA5xr3OIdGASm2yk37mZCo
z4jh8jH//nbCfYR5P8N4Vg95z6HtgtBhBnvBqTFwt24c4UYe3SNfcYK7RfJeJ2nh
uVeBeTotsJPOffbtpCHCLTgKJsb6U1SumOk9tjBdD68tIsvg4jOgJFxmne/POSlA
CIL9hy8lWcvSuWAnlc20raveX5HLGBAH78R7861PEBbvBoyiK4TzDdB8X2dd4BNZ
NilkqLUnrIeVaW7tkBYJ9HV+omEB2mf9hqBX/WKdQr7bP8tp8cSFLGt7e7TaCTPh
WQlOIX7Gk3imNiVohIYcEXL0rgphdM9EBXIZq3D3uspN04+Ly488BVXaW+JAYEEk
cEwP7W27u999fb7KUpW6xNU5/4gYYXTz6c+rXz7Cezn2KSXlRM13VswazRe3wbUh
rnT2m+adcuiLWu4F7UEaiKXVjXiBLtRU+ioJmygeURAE97O/xnuMQlS5o5YogWcY
5XM75WNBkuokThJB1h7oj/2RDhICeyKJm+poRHcY+1chBR0CYscWUcpGdcyci8wQ
cnKYEVIawG/T0xCvxMirRuJyZmts5ojCj47FYsQCRKkeSK2YEz44Y3l2wA9eTwTf
xE0C61a1FVdU7c10gbAReGURqkm0G1pIZsr+i8aICGg1n1lKMk99CY6VhN6W+xFn
inYO7VMbKoewod9AmlWnOb0ts58IqvBDJBt2Jjso99I0Q/eDyOOq1pCj4Lir7qUv
3xu/XMcFY0Hixmd+qeqBS46SfJBawHolR70IAryjEYQDwCLsK+HbzZsm4F7uRaPF
maZRh5KM1WGYbEIXd8tD5WTE40uQmZMf2JX9L9xvYv/VsA9RKwBCEzGQaZGSmHHN
gxgjmTVmFZdFKs6p/lCmJF5rYxDDaCWEsxgcIwZ3bV/Oq+ArPzeXY/bNKDcgqtMc
DvwA+Vx5jmcM30YQihGp/F95cAOfRW1D8GsSA/h7magnjwlfaiF1zgocvlykHldj
znhnAOyoLHbBvVp4/wd4RD2lSQeYDTizeFgMjOBH5Ts/8OGwT8FSw4IDUxO8r3B3
5rDLlbiWBfZ/kTTQm4sA+0ngGUIQHnvPJ1st6uJjAgmATYs6KMq2dMmh9BSyyYcM
9iMY+M7DZKKvan1Ud6BlE9XFyi+r8lKXCxkcICLwPO3exxOg5xyCypSdGYNmMgZN
yazzOQi0FZ/HYIGLSPH6G2B+W2NzodOon3nA5Iyn59qtjY+BuPFFlxKbuAhSkhWT
MoLUSMI8xMi6fh9SDHKINNNOlrG1CQq66w+FLtXjejvQaiWkPVbc9SfHrze0njky
SqpeAKn1+Nce3j0UNUhOlQ/UH0bGLoTRWNiQFPZHBm2HlcqEphkhSTgvYYgyLP8L
JIhox+kPaLQVGBCH2Adu/WvhnOtkW9Ml6U80anevXBsVZw7mwZTgE203OOF56QWv
ot2zO/wduy5KWJC5JoG2EsY2B2Hkv4CB8mv+QapxKyoCKxx8RdQkIAfFtIvg+Lp9
0AbMmNUAcagwS/jfCWTlZFtF2hHYSkd6qTW+YopaoZiO1UWzOvQTowM1r2Jw+gY5
XsUpEdR36CSZ1f9QQL1AD2ScVh8cin4kJTIzUq2DV/Tp2mVlVW17oME91z883wI1
rDfy3gNBsugkgPa5MMOwF9er2EPiy9OnU0Yfhr7ubL76CzH53Lqghq4B5U0KhIZi
QhvZv6wAkG61HdsKLqdCwfrje5KMpxbskqc5Z3Sc3heQuAAkEu2ilrT9+ptcepF2
JSm69h61dAozod0rSJ5X6T4Jky8BpT/TmghMphYdrDuIZV+nMXkPBRdS+5kTEDnk
Y0HtWe2N1VADe33F2sAfQt+yOfOWOy8atLovBn8T24Y0BkKu904Ni46XXUobHdaF
7FHSXMDfIQSeSV4ht4qMxgedLz8Cp1cp/SGgnnOWB55sn81Y39escjIQMzpwFYxY
Xk7ceQ0sT+BGOBaGWAz6T6cz+CwvGv+g2XydY7PystvyeHXF8kC/W7wJiK1W5v7l
HZDx7krxhMiDKT068UnGqR9EU1t84AljWXhI6UScdxUbKrXnXtFWZ8oxKf/0RQXk
0jAXe+h+eZ2MRDfPCYoZn0zM8ah0fog4KYkEsiWa22msDFb6qVlEAinVP2UsPFq+
O0o0GzOGNFJES18EXjuJnT7TRT0PGSocfsT0/BW6tUOEHO9gRplps8wMvNpfWd3n
kmb/uz++gzDhQdmFcBgWEspspPDOZV2Lwmmujv/9p2L4dfE9pp+uvqijuzacNPx4
vY7GZA24lKqgcQYFm4m6lFl9bDG1M6rLx9r78U7ehEE/QvZFRAvmrKGe8kpheYUL
Ud5hUu3ITgFaGaVTIHPwUQrvDAp1xALub0RYfu7iOlwnEgoNqh9zgcy1VHH1rYnN
0UFlnjNGu1ZWqXaQK/bFmN7XNG1CD02KrMgeiJgVIpcdUe378k4OZICkS/ovtv+d
EgrblBrLvzHz4ontX8rt98q+yVUI3HihAJBD5itJCIX/s/HKdsPy8QYAieN/b1jr
YQXCwu4oqEc0Syvea9ToDQNBisO6kTapUWKeOqH5I7du3rjgUUI2epcJIM7QbaNo
uDZk9ntovvIXpS18SE9hQ4sqTK93t7gHWTkFj4P2in/FefFZqTdGAU2wNGKBigJc
Mc5HaoCY/y3ufvXmIECrespiLmhNM7ALUBOC5RmqgacKnGjhyzSy2AO9b7+0F1EZ
pIemIG79/si/LRGbN0lFLHZxqnq8b666lk+qzKPLlnbpMBwK9SJElYsOvgT0CVTv
dZXlawhlFkFNNgjMghaLS449CyRc0np9tzG/TeO4MbvbNdbnsapW3JqxgLI132gM
Q9SlBN6LLMXpMemiOV+fpVab0joMvWS+aTWXGZ1dLqPFtwnGEy8YiEULkDSM0g2O
IGKlgAsoEKZJyzysJmFUwM51evMG/MFnN4YzVI/EZWGsHwnwLvyD0iGJtvL9k3m2
vK3fKtBvaGsoEHd73N1AanimCHalNrmjOFLmoAA08ShgHyYn+VmAR9VdIA3m4IRQ
xzVqkig1q88q8eaN56na93sH8VPqFHBzjQBYO2jYTF2f8TPpeCtxjUNZ54tygQ+s
g1n+lZ2nMYMhl5wW/Z7JUAg5+lfz8XGbG8uOll2J/G2VefYnxcOcEFimOS4FiIhO
raOaOEuIHLiOw8xunMUcQz7R/w4a2lFCbA7U/x8mVoBungS+X4R8aDaAG7qlqm1L
/gPxCJGsqxBTLJSakGpsnWcwrKgyBKqqBhkksVe2up/4iarKl8mDesHkf/Zjq4Vv
6ma9Z7moovbV+r8FfOeLZWGLNZmHZVqDhJ19jk+ourye3UglaImIIKIBKT9kxLu6
yudyAP7F8pYGhgdAnPiwu5wdRhnCdoz0bTonW9Q5RJ5m8K+yEkPNDRxWcSbUcdWD
o5mWzRDm2hNXmIwDTOogwqst/buEDT/qSj0ejy4RVvQW87aposwFxerBUo2T9Wmb
MS4fFU1rPJ8abro8C4xsUQb8xF65zscFTcDaUiQ/QU3CFogIKTtHQ9E9EAF3gdLH
W5cgnZFLlbKZ/IbiwtRSKkaWkSviKXsCo8I1zAG+rzupPYHuustDeO8YETm6Wy/r
9s0P0IND12uu093+4/oGjCLq8/n2nADKWhwb4UCwQSU3qegbhLmLHxjK/K1+BG/V
EhmVcyagSh3/kAiYcEGUmNlm+0ZJXpWHm+gOluqk4ltcqshfl1LpM2yv1vqg2HgQ
9z+NJoONhzEEmGct7VV3RlaYtq+6v5p7WRZhVIL1WRdGHzFkbc2QitIx1LRYlNmo
qihOjHQKjhdaeRR10yUEIF/x+Ih20MqeGPqrSLzR/GIsv4htnEmXfSlEPg8q0sAL
z9O0WgoJxT/oX9FD876z55+j8f5UcwV+11QkY9FvKHfxTiuDZogI3n14B6A1Y3SJ
XQDYldnraCYE/4BPuPgdllJR3w/pIBmKfQ2pd8HwvwJ5eOeiviD2ZUEpsOi5FaFb
yc0ezyL6vVW00hgr3UOYoRxCstpd3GzxGCl1BJ3OmCw23q+1G0IXLaqbIkBf9h60
FlSXHiT2gaYv2wCzkKc4lTgLKWs0911KH4l/PPBKpPqf8EEUdiU92oPOJvGxghxe
MMra3ssZy6bH0mxBGuhtywZ2XVjRodtntZBe2KU4OsGZqPVnrLFUqEIgYXO0DALJ
u6vfH8/GmOHo03XSxxu8u8PXilsAYT9nF4OHN8C51LNQukOR5YNSt6I5yjIihGNu
UrNly01ec1Ycq1kChWsOkVb4L+za0UAilLJdXCk2qNUT0hoXR2EeKRG6F81UJy1x
R3yY3RC59FHRxUTqSQ2eZTKwzsmXj0w+/6l0nquM9FDtOyLipkBb71utkDBtMWm3
+CYHQQBPhEI5yWMRT9rnNoP3g7Ipexhyz8qfvjbdvlRYUCB+Odym4q43PHujdoDs
RztYlnm1Dq7v/W3lFOpdqsJa19p9MPop0JZ2OpfZ5LzOVTPhhrpt7rMaXLv1rUX1
ucEUuaWrqdNz1oOBLiSL9VMKBpx8SkjSx6OGQCW6iT+ZlhciGwOJTRF4BzY5+Y5K
knlpvKGtV3nYd9lGoMzxQY/aQRpwuEs9loEK2XiraYo+jhQKlOo1647rsnEt9ksB
OEYA6SRhV0ABeMsjFIkUahZUCagOG+mvmqGP1a7ZQlQ4VJWrmgCetoRj9M20QBTA
36pzizzQ6N5f6tgZKNk36OQOvjL4bMNU+C+eVANGbzN+GStiIp96dDKXpt1cIspG
G66JDgFudfPH51Wo1YE3EP/ligkpXbQSPN5wK1dDjsQMrvjNwAeA9Al1IzSRzVaE
H1T5t/HLJ35OXzsqaSAYKcZHPLqnSf7eZ6jC1vb6u2Bk0whpQQuHRM8NYYgkaDd7
SbfVkfzXutnpwq5+UIGx8ORJHj4smSdK1AX79hX4hR2vOYiWGAwip/Xt1idFXuZM
da4PQDNoH5bfAmz1XQUJgT6foswSEUZU2YMNfvtHPkHKZ+eMgxUFpzncCj3ixjj7
RoAacT2LhNkU8x9YVq4yaWJP5tVrxxQMi5PNyFUQgnyrku/rIrdQej2ANlJ7swmJ
qpWWiB2zEK59XEoeFiKa4qctk1l2bxS9oC3iCCCvDgEEorP+IAYp07Bk2yJiFiFJ
1Wo2eiU8fzQmJrM3zr0x4o+CqKgxHW3BZTpmRky94ED3g4Ixvhg+8XLsng9cNwhR
NVcJOJDAuT67ZVfXRTfKqYYPzQZWq9uOoxR/c6DQD6wcak+QTiwYtguXCezh4Enr
qf9goft2vVDYHdQEtQTEoMLMg7eKlOMWN7Unh1LUTj44oSzO84rms25O0fTLZJNE
gjy1OJodDU+3fc3eOKecrkzjmiIxmO1XqJkUxzAy4jT2L5KLD7C/XIUiCgiX4Pkx
TjAiTIXYONf62x1mO5cUdN4N3k2GvZln1DYWCfVKe/ZnnIkeUOx4ICVvnxAoOOrj
dInfG4XhPJUzNnXW0IxxtBQsx/UKr3dwBBy6BAmrDwJ4YFgtC7xl2mcpmkwWUCS6
idKGbG6/jB1k4tfhG0EOXlU6JHqp4DhCO6FtymR3DQupHGBpxVGTEPrPcj9HuixS
ZfKgwyj7WhP2sQOyh8+gDdcCIm3D/81U2XyqvZTkc3dy1z5A7a8l8CPBjFiVBkqf
TlXyIBC9jzFfVDcxYeQ61ntIwwhgDHMXSQH2dTCeiO1Y4NcO/3vEQH8ukjAuIlvL
Om6eJfGWOR61DBr3bBVkpPFlR0GGJ/q9zCmXhT5im6uAq2RsSaCdifpHR7yKcK0g
cc+KYtTlu9CbGcMzRKpH8Ikiaf571QuqCR5QfaosfswK7PTWSaypHWkO9PM3FSCa
yY2xPpidWYaTBGBVhciR9Tsx/T5QPiQF+RZ3eu74MCRI1gODomDIV66MjZEAiI/t
Tag1lDtOsaIkdxGiqBb3whjRAZUe56Y7vEm8J1sJnysac+dObJthhK2qm9f9qyAr
ZZZUtAJQ5isJHj/Nw6kFzyyDwioUTNS3x6bYmN7nF5Bp+hEox36dutA8U0zbjas4
1ZvEjS7v98LIKv+0rj8Ailk4Amqojs9frERn39khGO9oYFJrk3+0h4ZrEpSVtLiv
BP8+8OwomO0+ilpXD7bo9Q8rSpbkimVTLuK+1C2636a7vkIaaT++HjN2aGci852u
AwIj3FYVGxBtTw6qxv1rddpS9TTy3yUepIyMmjgfzhJXWpFGfimxXfEcNqyQVqFd
H2Y14I2jOcFUzIWmDlYNPd4tibvjRGyRSxR1tA/2f2h/xY3m0W1u1jvwMtN8pVKS
Qbt07nt7fm5j8JEQh7chVNve+WsLlXHTX7CpKjo4MIYj772JmmQFJoQnFXc5lgV8
WtPtvLQdgNSTgfdqebaosWGGiLby1LOXfmn7QhYp1ecOqx4jhMq8qqwBi89gB9Gt
WLQAI1zkXsWxTAzsWX/kO3lOorbAZ8hc8/pK/Yfq3o6qzMbvch4mi6sY79VifsjX
d+KjoN49ifZkMJKbKEMxi9HJusFr0L34JQJQetbTbJP8zul0yJYSag8HBcAcgImW
Cc0yG/shNtfrfBcmhs2CgIZaSS1WWzrEo/2QoJSXBRsjdGT7TWdj49NElLMR6gYP
nKeYxX47HTNGEyb9YuGdqKS9OFpZrVdYFXztsOrWvbYz0pNy5CuV4OtVcuIXWtRx
FooKC77zvgY7Yibk9sCRYL0L+B99CE7eSiwFvBLwx+lN4q1RrCja5vuerRjlEYGo
rzANhDSwo5avEOWfdmcZFTNrsxc/ll5qLTHJI1iYnNqB9d14AwDtj7KaX0dCIQUP
lDU+oJn8190iJSaYoigebms6rUE/H2k9t1aaxqipvGi8xNHCT2YSjvXCsOOp7XoH
Hb+dHiDRNti7ZMo2Dvur49hQs9GHtn6Idc/hSSKVRCuL6LWJkduCA+7D1RE+Ucmq
4itb16re0gYWVAeMxoWPd766qpGqYlHg/N5zUU8XzBiB7NI+FYdr53dEUVW25r4i
0wEk61vLtD7xPon2SZyaK15Xgp/wm7I/rYsjBUgBk2DBdtA6NXV46F20A28kXZg6
hXmHjI8+h4Hn6J+K2AXdsOMgK1aBSG2S5mZyhBXoPnNakyKGjxNh6tT0hz4Ynkk2
0tf/P5Yahfm2ixzfK+LtMaA8m1HdNKeMjUAZ6gvrayqJ3ghIWP49NyfLtdqaPG8U
M366zqiwHLTD0HoMShFfTJxPuJgAucNnG/4U1oB/RcqJTSnGefNnlsfjnoLL1qzq
1EfUXY33ukhCCjPzrZ80nqbfR15xrnm01CI/maXIU/iagSAB3ZHTZiHKgERBTnDu
3YzZ5Tbc33paGLeMT3l6U32D6gYsJRcGgRpBzzZYb8r1IOVvTtRaay22vMtc8Sxg
a8OAMmK+JDjZX5NvW41hjen5DKDwuHrm6PFNuYA+6wvBaaEqHDalWirVNuvPsMB3
ZAVt5NLEwxLKecCyiQvHeSJKHzvHi2OoS/FiQmWS/d/AGi51EDdpAwzp4qIJHy1k
+UHUWwy5PYjTfRaNqk86tklJbKrPifuciI7zimOB0OJcfdfTDlPKesP7i4IbSTDY
UupWSV+8QJNMZYpg1UzEUo/ruddjYJKku+qv5pfdSprmtWIpkKIPNuoYleDbDyuL
DxVai7VFi1okBlLJaBzYp+L30Btfojt7fGfABdU911DetQs159FEbSaWnU1WZNtU
BnPCqEPJlT3HNh2qGofjMYi8vdPj0xtCPtVxQhf241LDHocebZAS38ZYW+pL+i7Y
4RSzFvZ80xgj8q1ntKgWyExjrRtmX8Gukhzs8sHEFr7qFCFHEdaVRlJEnwlDuOTq
HpL9sL7nwLxfbfNxdXXzSypx5W4bOqNxeqfULs3FH8gCZNBLc8YMDnd6PavrfzcQ
zbHpJyu2FRUOXfQCyWBeLVa9+4FmCGS8WQrFSVGZNoc2Gp5qkxr4fwJxjzkVhqUl
yFtdOc2oD8uE0qS9UNfGsSYzf5XQHF+oR/c7vu+iROkFoPuzkZq6fcwfhdPqY2Bs
LOiFY2pvwMwlf7h/LiFg/ljq3k2C3HEGvtnUM/Ch7Z/iKpDvSRUdqy/odQdRPKO8
YwuPC0xcyNq7wcyyCzPZCqZhhXc3l41N2LhrVMTLb5sNCHsGcRH31WHNuStlYh4U
TSHBKkrxVyNqdl50nWu7e0nC+icqbM8F0VOKCuTtBjRAbtb47yVcf9bcbNpFWsC5
bcHayJHZNtwP8gsicukbe2mpq05KO8IAEHjhfLdlmbAjKP/zm7TYt4AYrvCanrmn
hKgv9DhJJJUqmEW4j5FH2fTjKbofLzLysWUc+m9GJUUuPA6vtcexCJlPuSamhEKi
uNySrLUuOyaGrQ/pfD1Tg1WuGpl6TzohuM1yaBDdgiijAI+1SWK1iB2bCEGEWP23
0SaOYskDSTHutoixAQzDqC9mYcG5SC1XEbrXr6jxTs4g2fTHVuklipqKNJ8a2WvK
KaMdptTapRBQP02sIMuDCcqfwLFiGw3yG5kDXiFFUQ05JOwRWlINYHEwaWwBPsAl
Qj3d2Lx6g/e8nPsZA2q2M/4+k9EsjQCPNdGuecY/i5eFXDCeG1mkfaDwtm75ps34
RuOllsBSYzTxsJAnPIUrEppRLE9MyKSadVIjHKg3Jm3GdxSMKpW3W/KaBfhqo9mu
e7ToQLucqlDas+EDuESN602suKguafwotqqjZWeoHZ8GjwmsyBHiRRY7rY88ptng
IFvi6uVaHST6ryfh3eA76OruMo4mYaTxIpfri2iP5aPQKzQANXdJOkCjrF4+a+P8
Pj+fmpf/pOpu95cuNI2RTxraO0bGUE3iqNi6itO6LoEqyyGDktYvhyt5SFPx182J
O8nTTMwq+zLNKkWc6aMXgiWVJ3OMLL+KyzEx/PVwwHsOxQRdE+O/nkCuB5FVah0p
G3YLTjVUkNxioMHJhnvsJd9eWScVK8qOndFTwtRtgTDMtACiq3uEUG8Dl6rXja1y
X1t4qtAg27KlWpwpziYC+WDp4wmit23jSfL9xLu6Vt0RZXSWmRUavOojSUaRw2Rv
0696JbuK/ejtN6q0osWnjNWGeXLeuPqNszspPjTq4wrU9yrp/niU9wFpFbr9LyO1
7u2TSksFTnSYuIQRPgUgijP6yh9s75Hnr1iP2Wpa8IN+hCuq/+sf6fN1b/ChHISr
Bc3RmLXxkDtf4LyNTfPzOlr9RfKpzawAjIHOqq2/S0cUHFc3oxepy3YX0HORf0on
oHE82ARNkX7ev3N9260VjFScnICrSCwryGNNt/asAKRtAYqK1IOOHftU9je8Wymb
UEcdKFZKaog4YGC0yE9yKdxwScGR3gdc6Dd3+i51kCGtGFojjKpXvyYldWF/cS1T
e34ZH5eU0KJyyEV4WDToiTj2IBJwW1A1uWB+GUAgZtaaW5KjLJsDsavZ4ycwcFZy
0cdUujnL0DZfC4iI7a4+W7zcnDEowBbRiGERFzdXgT57jFkUf8GC1IKgl/uvogtO
By7m3hpK3NtMDizd59ZRlUzYrNsxO6Df9RJ0mSHabGVH5VEY5g3hz8xJBE6uwFQo
jJtmw81cRNMEBWJRoCTv4iDMYoATs9cUXEk+j+Ol8+BZGkchd8QbYtc7Egl//s9q
7mL1TPiT0SK/0e9DkljGy0eUv4iFCCCzefyLQt7tMn9DtWhFTOA9/fCb1ct4slfU
Ow5pfiuiJ5yk/4m0LVk31lpIPSfiGvH1hHI833GX1DY+79jJuer7pB1Qm/AybXq8
ueVxsLW5GQK+a8Rfj0FM2oA3skwSGHUl8M2iMlxsKJ/wfFuQ08i7PVhYmHUYUHr3
AAyF9X0XOsm69k2iinTmcL5Zw5+GT48umV0M70WgY+SH8+E3zCkrSOZo+7MVZl36
mJxB4EHIpqCVgqRANxOWDKHZbFItxudfIzoYfGirT5VjlgIwnqDYGgrAaZPbD5PM
PJygeaNoE2vvhdO0biKuvKG18+L4APcmG4p7rO9FclYP1HwOO/Ddhk78PJTxGYVt
6W923FLsFY1j11vWvV+gXdlA9JxcPuyxRqRrnw7PreutzZiZb0/q6WsSWuSDntWV
PHbS0zP9KCdrg/ENx5CIBoXGa9TWgqJapz0VeZ1dI3uKpBvy2MFyiT6rWuQV0bRm
5Y+/b7VP1NcZI3Kfrrmdm9YeXSZRzovOlBfkieCqxZZCsADZtxKLyVy6APAgOcqK
RxBnLE1XpfPL6unoAP+PYEjnfV1gPyk0PAwIAG9bcz+0/YM4u4jgl2U2X3dqza1Z
uWo7CumAhymPpX0IbxmgqEU7oE17lqaS6kR2JXKeLVs2/uq/jDnKbz5YNJDHaBHs
utadnbin/2aDxqVom7aOWek1gfSczBnj8Pg+jXfkeC6EytkA0Y7OzdFcm4Z64Gi7
/meT2ITkOWFHMyUI8T+6CmYhW2eSIqyGUTpVz2RReWiKGkrav2O05MIdbIgHtjNg
HlLt3jP4/IjcOTf6xu9OXOpkYSI0jTgCIHxs66z59F4o2TR6dBJ04YMIBdc4fdgW
SQ3VANYpPAj/6zQwFkLa5cZ2DlVrzBi4y2Gts8XcwD28S4CHBHSmkVhD+q1SQ4ob
cN0pkCExxkdegfJvUsjxjpFed8EUenqOHonJ6RGvYH532GgcVaug1yCqPig4N62O
Fl/yjPzVOdARcXc3K+z1/jHLMGGV0XUyu+KpSMgsMT1ElA/gwA9u2FCcsdZhCdtS
mZQqcNSpkYCDtDa816KXbKdrnF7iwyFZCLQVmf/E1YhnFundhFq96TMnw8ZWPK4K
EZ4vU9lGfOKZQ2+PjwW5SBz0+nALhCsQnS71HA5AouM/xnreXoOD/O18i0gT2bAi
pMPWFUNEwZZlnkDJFDVtyiyQ332f3ciCaKowiHrUKg/whzDledNghm+BfbTAWaGu
4yU/GARQ9XU7G/Vk8fbDSIouJKqnRXsFVOADl1dErmz/bBfWemy/gWLqox3hM0+P
vH5i/a20m0ljwEQiHmD4be53kWO+GQL5y0N5PlKifKWUTMLeqmrED4sL751qGxag
VcAZ0/6BSBXpTD+FvLH6/l6bZZF4N/ZdACHPE37QXrKLhx7Mgep8xgp+1BP8XakZ
WUzo20kjLZBb7rOkcPGAixP0/bY5xM96uhFH/gA2m2c34YDDzC6yLzHOlreTD0uu
pSfAObST3Lvcn8nVe9YWEdES8fR5gDGViWkVcph4dqnpAfcX9nOTw1oJ1sUEDp7d
lhjlPgOEuViqUIkGFjqpvIfDTcTvsFf0To7ahmqdt1/KX0qhreoN2HBXPweFppAm
txQ/brHzuiNItsCrXsB7sVIO5mA6fWmCregYeF/3eDmRvRYbTIn/p1YvkeBLxljE
BPUBkPPxehh3Twwomh6/ukzLH8LXSmNW62eaWZMTkEEF6yeGs+s47i/aWgrcEDdK
BGQsSIWeTBcV7QHvt02fh5a4ZuGvfAMnlqRqH9r2idqIb4nvuobZvIXDMO60IpzM
Wm0YluJQm4yTBTkW4LtSzImlsJLwQfBhrmwFB2lmXLNVocWYZPRn5B391A5bYv5d
tA46cLQzRNQ5vhFoVS49cynMv6GvjP9nJ/gVds6ErQ+myM67yRTfCZqoS45wdyv3
ktU1+QLWeRtkhHLQNbH8ZexHK3rHl7rkG0MB4BNPnEfHMTyG+oVgL+usaxCYtaSp
M0pQSYtw5bEBrYrqLauEa3MD/CpHbaujpecNeREdKKl0H4aib21opHOMtNR5V0x7
3o9A/C61tRrlAbYg1foQhpcXqTB1c7p1hewzJHaO0dOK4V/Nh2ygZHzCVXikzTEj
z5xFww+dTHyqit1cfAldBOtU3uu/Wpke0Kt94kwKGWkjkzxqHs7T2ryUuLnsGcoX
HU2iQS6GM2FCoErCRmePlJ3TjiQJohenthgLAC4zu8l+rX7afcHj4p/swLlUji0p
Oi7ACRzrGpvaP3k243kIt+Et8GilSyAQ4GOg9IcD7ujuhQ/wEW2RdORS5DzCtBhC
fIOLNnxG94s6w8QNpy6+SApcAP6vf8LVhSQRNy8etn8Feve878QU9+bMRr50ESW7
MHk6kWGxOROSgPg3smPA7iZ3fwyuhDv8hwHN8+5osKvzUOov4muI6reBPeRkxLmc
UcmGvOn58S2HBNJSGx1CcyCz3xpacVGPAQXkL6DUdnTDcl3QpWCu2avqm0GyZW3x
S/7kExvncQHsQy4EwZTWro3Imuf9KfUxvJGgKmUAHmmHnCXj3DwrML5JWrfXqmiR
Jhj2GfdHc4TVMpSSBGENaiy09YX5mPAeyLJv6JALtYBrPbmfdeKmTO12eGkyFhY/
ClOncP39r2rXGum1p/VICOTPbVb+ekG2nDV4+AUPnZvqs6vJlV2r6s/0a7u/1d3U
MjIleBjXYAj7ja6QubNfynh0MnESYzKvA9iFLE7N+ebVF1wpXzrRRildmnW97Oqo
VPDu8rH3oKI9irh8l6rnbtUF8wTD9RrlZk7UB5t6rn/3Lxf7XJDROJO501THkj6b
2CdCGyAdUasDXyWsbDHZ1llOlz36/EmBizycpLBLrs15I6T7kVE7ob6IwTo/NXwx
iNVd34lAhV4V4ypa86ZCfG3R7zr0cob0NYCJFQ7Yi0XqUAGI5UaUpzqhBJ6R1CeD
SzziPjXZDvvF6bCOJ5OqTdpj5+XRvlJnQ2ugNmYItZeY67ZvPwWbn+7aGNAq9TNg
h8rig1yidFRmg2UCO7XZ0ehIdv83/iA28F7g9lHTu09DktWXmdRuv/hBzYB8qxyH
cBNcZoJUvklOKMQhNm4L8xFh8ACdG0uQQfmlIA/9pyXEhptcRsbztJij0Yr0PbSm
+nQrBSCGHlq/6JWvZPcgPHXNUVCTVXHxHIYpOaescjRr7y0w25MEOaZ1UU0aM7mT
h3ZgcpL6+kKf03GP1loz+3TA9tqgVyvLUis1O5jr5hCrKBx/SHNE2D2xS32zIywQ
OOu7a/u3MgDAxC6DhYnNLy2oRwnPiw+iONITJkz74mjMgZSQLa6wBLwtr+ksydfy
fjudYUU7LwZKkGcsp5NovFp/m2kRlNJmTD2iY8J7D9wJFOVM+77kMQxVMG7msffN
x3Y4kId41fEhEjhv3cK8RlrOOa1pZxyTiWEhbpo0JsE45iZpKhA8027kTRtVustp
c4NAeqmKI3tCUb7uoli881zLr9XEzmeNs4+y81T63fE0Qd2jg95v1V902O/QzzoR
zI8zd8ui8rT0QYP95amHzntRBq3dcvd+AWOSsdlhHfNA8HJ12f7nMXxXOKtJ8QdN
xBTqYx5pg9+nPsLpL5jBIqMqHsnux1bcBjkOPDOcIcALWNsEiinEzBhT6qGtybAD
fHFTXLmyDzcUOleYpFt0nXYuTVKCu+BglNTxxoldsTd+f4zljVqRRyCU41Wkr00D
UgjJ8yNdiI3Zn7XQZdObhvdNdvZ5Nqs/O1RqmTDGxuh3IL5XMG8CJmncPeN4IPPw
Z/ktBKbJ5p0rRi8U9zxsAzVbqaWt5hxdSXJMhFFGCnCP598h2Zg93aB4OwdbPmmR
v3k81VKfUYUBoB3h7ePD1B/w553+3WstTlRPvcUJxW1z6Cd26WaExtJPQNe35HAm
wqMHsRNwHkgAQhyNu8ZdcDMu895lTtJLavOlFuRHBb5fKVJJ9COaofLmwIsqCGbY
bZ1Fr/jAh0xGZYnwjdasIRFNYykDOS1E/33cVgBjLvHOuwtKJbJOVFOeIHJEZ/q5
a4KVEbWuFSUz17Ydi2N+fxd+E6eIbZJBfT/U7HcxYn/PLezkn01FuzO+ZBfF7kyz
iOJAQ/4H7UJ6OOt7a4JqJMqpwT5Fngf++fJ29NQvEiMZWOcOI8yl23ql+Zcs5x9/
EdvU1vvvdNwcNYjrjw48ZQbhXIfy++ygI9wL6EaqUR9XIQd7Q+SzxN+EK66F4Lbq
j4R/arovCXw2UCBift+bE6Ap/chg6lZyEKsXT2YEHBJZBaNXOs9kV+lr2BokvWC8
qU9nCYoSeAx2JiQw/I5j4Vvrlrbf6JX0F+nzw746QVfzwIo5JaH5djMGGGSpmA9m
nxck0IVGvHLGe0paShwp9X1OtJev/aLzv7xF45ZhHu1swoaSl1Z0QfJBRXWcnE9F
fp+7qzaqY9C87GiS1NqcZNn6Y25PQbP7yn1LFXsOg0xatsnjlMyPWhZfSb1jTe09
aT6+UxvDCwaHEuTqULGYSYn6YV/AKVbCp7/QXheYvWuweG/bjXwdtlc8/ZcistYK
5pSEEG9oUKH4evNM4CSa14EVXeASAMj+t4RHN6L6lfsSQ6qDlwg4mWyOUnuCH1gz
U147rQdH1Lw27vaB3L9NUewadr71JplA3JsvfpQLWuCzGbARdlAuH5Rfi43XDUQT
Oami3f+62s3ffieVQ48hWRgrT4x+y7xkQiMpN82Jue5btGRZZtWMkPEdNHdGl0t3
l14KzynJMNxGIC41H+V9yCbfIFWPW7uCLP/0vXbFcA+lSDRZu7g2PJkC5raFPxt1
mBCrEs4mRL/8eOsK9vXXPYPRNDAwlggm2Ekpsokii6jroZeuWJLW5tMXQWHxjYJG
UMrsWIahKJr6YL2EV9fFvaFOUkPe7G51JUfmtcGwQ9jLPk6QIMfzbxabUvGoWN8q
vHJDJUgywsTGX4lvx6NssWQOe2Kx36NmUL49gazEQucj4VmU4RifrLff5Q3BG/s9
fBvL2fmWVsFHmIyy2lVPDZDMNtKnod3oShK+6mG5YOsacCNnXmgHjveZG+RK/T1i
+BSSxZAjdcE88UubHD3CE3/YiMo2mtQ19Fx+x/HelwCEcmeGKuK/fyIDD7TAqueE
KNj2F7VhodPGlfRzHmLwie7U9FxN0jaAlrWDvaxNN8nv0nrKcJP5Kq7xRwMgUq92
aeOgs8BhraclMMtB+nRgOAUEK1AapHRFeymahL/n5weG32fGVTgrWTwbeGJsaZ9i
QnTVj6z46UquO9sbq37CQfQPNvor+HzEGmB5aFP2a4JYhrb/RE5FkkmOHcPplhMF
lCX1ZreEXYQ6zFW2UHk+T39LMZQGC1B6eTwVB9XeCgUmIRQKb1AR4oo2bx1Pmpo7
ddsGnQS25/VWzNqnxE950+U1VpPOcF5PBfCcF6Zuunl2K/a16wl40Zlx6Rn4ZnEM
hK5TYcohAU74jVYTu3eSoa0/8JWXYJQvsbBGATiBQeuZrNJ2v/kIbkrfKcqKr34D
8WBu1AM5L0vYQEjK6CEvtrjXiZa3G9BTOCXs6DkMUj4K46nhAFn0+pT3ft/h5uTl
VV9yLGSAqDlsfUDnAiZUFZnSG6CeH7rtQkTZjcy6lFUGSF5flMLHB5/uZoPHRFHo
+2l4Y7aRlBfljFuPivyMnA5TEjGm1jTRRRZK7AsqkV+KiilstW/bPc+Htlfn0PZ2
S+AuAr1rkpyc18AbMPcvSh7xP25cSSoWiA0ofK/mFd4ybdQ9HcQEDUhBbxudi5mN
Gklf14m5eMfpmWrYxJTIbDAyfgYGmUnPdubeUOw24PBxXjY5tw1BITUn9jQl1v1z
fepJb+YxttduwNmQg6g29l9E35LjOXk3+IKzbIRge40KmZR4eMX721TCjka11hjE
706gzmq8q36O6MfjG7Ka1pae1yse3dv3zwrx2m7G5Jlmy2xrKm3T8z3wNScP9/n8
RwZxcx20U5wHTgdeOW4Cic5l90B4YRyUGKZKXhoJ6ii1zqH7/ofY3tCt7+wErNv0
AfHf2qrowKOWHSRRoeTTdq8BDwAEFyZf/FXVDju8t2fO9w85DVJNoV0ydvVuCR0d
FPr+Ekl2qBTHarC7TRNxVNDrc4qq9E8MKL4P09d9ClPn3Kg09H7S3MagoVddZxxm
5deSddHaahVuMQEaDFXrtDfc0RNbQwVyE5Yn5HNohl0A6+AoLRWxxUserbbEwiQM
FQLmcWp43T38+Brh41UN1nqYaAWk8XpijsPt3O6g9vMb5b56RT5lRcuuRqOYY3pr
8SWl24kdHpbJDmjIAI6OJlYO4x+sAvQ/9q/rkXxZt9t8HcY1pDmcjzCULVfVPIFj
P6Bo06olJmiFb2JiMKPmeCrIrAayPisekwnco17t7WhhHYJcDq/g3NTptb1m33E2
s6QapM5xERyCSOgAFdz0xBJdllEpplIAmN3xmH4rUScXFBfnJR/mWQDZmqH52Smk
YNHnOpsmgPckIlYdYAhFEU6y2I70cfNxzJPhYxH3hGdsgG1n7Mnh4dR9yWer2I3t
smovLVnOoM105X292PEldvLz3C9kTcgWtme8csJ0nnUVFNm4+uXZQ98U5aG8MUyh
ArVYvgBCI+Y3EkNcwvmvkDWwh8/g0F+5S/dpnwy31YzUxcurqzu/tR4fvvF0OH6J
TvYytc20Cr5mGIuw/HfS5ymZlgOoA53rgAslEumvSgPuO9C04rb1cozqxDLRWQ1U
NpnILE6/KZEFJk/LkzXk0Dq0FiFRsbpiycyQpIYAW6EAaJqI+ooNtQUzo+8N2g1+
+IAWqywdtL3Wz/kIv010ww5mbpp5o/b3iasXPlxlL/u4/kXZO8ULEScyLqCJlTWn
AmduGEvVtB5GrNpbDTuR9tcg8JTNv+t5a9BIbg6V8PsDzaIqsu4iYiMfQayZY0HE
mODuvIES8GY4bLXLG/Y2CdwzeDpUBGa4f41M20lg+daIqp5mcZCB6Dtw5R+3wiwl
T7YQ7PAq/opMQJedHmnsY/zh9Lar+Rez0Jh+p8MmXp9P3jSZdkMyXUdDpSx2tImS
W7G5xDUWZwqnWpbj0ZpPGwXPew/6TgNb+1u0dMuvdZ3pvhlNlHuRkrvBUdX4bbN4
ISikFH1EYMt8Npzd039XqnNEbF0pDRKuTKtiaZN2XaNPzN7VNKu4flXRhXG8yORb
w6HQbgFAWLA8JcNJWtj3YGKuLg4hnU8dbsWDrvPudUok+BIKg5pDTO1N9eInl4fM
XE6YahyA+IQgzwfDkxTgS35WG68Xly3RjB2zTG7V+B3l6mG8pLCmqatDIzpUzU3R
8556y8NDS30dJkl1uyc7K+xHaOeGdtSzytD5Eiy3+dnFNQagwYMAkHiI6KHFxgUx
3MRHTZ6/JZWxojdaXzoVF7XtzOuZpE7uWa5qDtRqAOg/r9i+M39DC6zhSzD7c7X1
yT6XwGSzWdPprqyxfc4FppQdjATLpEfEOHH7AuM0S4GtdQGas4YgyvwJarHQFuUS
OOzR3Chk9iPxT/WvBgcBbhE1pLOc6GkNN77NrlxVmwhSL2ImQr/QcH4t7gimlb+n
xogCBeSmOv4F6CLrTxMpy6RzCS5No+9N0VcA7GSKvJyZkvISWBZDsInhPalwXBcM
gx+v9VFUNwhY4GkcH+eTrpl7HywQXj97gutf12c00bri5cLjMwORnxZPFfOqU2QZ
F6sRKLeDeNBrCU0mrIoWbQ9iypgJDyaVMytkwuD+d4chhXA3SXlcUavmkXQrvLj/
Ua7uqGZspASDYQqutfLKkmN88yYqWL81LydkAIjH5pIFJeVrQEh0XENyHhOsIsfT
mGE3jMIs4rh+LMTNu2k1Pp11EMn5WF/5I+T/N0UpoPpkln4S9Ftzb68PWnaFF6Lv
WCgQIh81GMznmJ+JY93AyaPTW8euCfv+kxZpcALGaUxWCZt7zFKe2tGKkkT3jwKw
5RDmGjmuKdjUsmY2u/KSbbwEga7/Os7K7C12CyrM4b9RdHTm+a6I/mXSkX2WDtuY
k4GS9nmy8UOT1H27k6l5hKgs/rnAdg/JH8HD84t3ue2MHfMfCkCSO9hiGudA5dzc
UE6Tz4jQ5yzssQsTM5RQW+ptbXcp86lhOvDl19TACkl9R1EzAsNeald4VoIKu/o8
g2uUnWAnMRceUfHZvLN5HXOO80TKG0z5UYTyXTYTsbH9/kqFfVePcL1M460RywPr
4ltbo5RMxVBrXFqLjgSQn4y561k6oVrVOGj/AHr/Jm09xuUlmWW5R2gcQtyS13U0
7hfW9WL5p5NdLgm28imPvx5CSmLqgIQdSDKIN89O97zY2fMMbvnDeHXD5TYNgSKa
BmV1F0pJAqiLNC9ZWSkTr4f/lZElqqWwh0Ssg6tliaBv8L/oMnqnXTl9mic8RCQl
yEikPYOEDaZ5tbZ+9UKWshD4egyQqJjY8aA9psL6IT1VBk6U5opc+zsVwQXCX+ZR
5cwrz4gfGes9hPKgEwafeU7H2fdcBo1aVyvj1J0AuVoQIF8ms9jHrqzq46CsEAZQ
iv8UmOVmkGMwQiaroypGvCaMfPfl4p8g0ZT53YEzj/jeKucR22bsikjimRqE/Byi
zL2AfSuB6pBGH/WVik9SbIR6XnVx8+ZuU10EnXu2VsO/Cyx1LHv1uaCv0SV6X357
yHG+BaJe3yIMq24ajEaujA7XZAXyreb7BNZY6kqreR3tKjPPfwHowUQ/IRY90oPI
6vBlgmNPinmGgGCYUI6lcbxqaWZFnrQEYNej+rAGzcPkDm639riIY4QXW5tao4HK
7z402kLGFnILbg/8ECuMoItoJZgXBxV2DFApwe1SqgxeJCEiTercMTYbo8c10PAt
6joEySjP3SW77h5pgtftva0lGiGUwJ7keMCFeoRbG815hvkdEA9Zuk16W19gqtQM
EJOKrve9m0CBDq9himvCehMxNZ+mDRbY8DuKOvtUp6bzL9uAiESmccD2vVHAgRzL
dV/QR6BZJuU6dH/jY7wEY/u7xWp5UFHN35PeuZ0nsygFwoo2hwUFyfPDi94hOf3P
C5bVei5is6s0Ak5tJHRqHRLbbQq8WhmBnW+NdZPnkejlW/9PcNjCX7r4z2wbhc+I
wyA9Sg4TZg6GrMZy3RgvXQCUT88ajFAa/cgEOwxqg/V64QlQegdl4hDNU3vvu1D0
cAzYXLUsQKy3NOmGHcrtvhCZBPK27mwX5hgFBEQmqvch2dVW9M8Sj1O3/uPEje/R
P7LfMZ1QlnATFRxXPrCCvlpzBAtSjmllzuLriNkh5AuzFqd5vu39lZOokuzhhaQh
WAe7RlvGv3dg+7YjpTlhKJ145xts7F6DxIQT6BjgYUqZ22AYRedng3iKdEtZt3Ul
wrpNdCIBR6njT0gbw5iX4ZYM0wTZGhr+T9PjfQNORO2ObnXU5j67ERt2JKWip0IF
CpYrnQ4rxBpxbUFkBDeEJ9pMmFuE8OhHjabM55XrTj/jdjOXoREtIJQt9yftIV04
iRcKP300n9XisZo0OU4t2zNLaUL8cQfbHn9cJ4POVdpOdUs4fRzx+GexT9dd3BKI
b8epJOUHJjuygQ199ElTQTrRSloqGkj3TTe7JoR4ap1H9UGcryxovPTuJT8B8J2P
UDBWr+rfjr29hZHlNsWZ555c8N8M3ixF194ZeWUsGuEo9ny0IraVEbFduPamnz9L
wbNiPb3BwZ3PXQHIXA39uh6CmwWonptmHAj7SX8rQ0u9bcIYJ46gjpJbd3Bb3la+
nGRNriXIJ0XS7FXEKcNPgSZuUTvGedv6W4YD9jPWYK1YVOOJl4LH1BNb8AtZXUEC
qtWmOJTFBWl4Q54RV3MIo9PfCueMGkHcEYNdCnRxQgsPNJVER2PBe28WtRhul0Gn
O0Y3GBGk7sLXRRcarsCcoQ840vEF8lqw4G+cdfsS00/mSubVo8MAag3WaETXbG7w
C3GFUBZqcRiohhkgUz44ONj5uAiXJ+hAdqQydgnw4p4q/wCl1AYFBVpNlBHRiAM5
mGu2FsQf7maD+V0jcH/mNYUZa2Qf25Tx2D2PLypdmEJgwcvrDrcyEIctSFuzxN0h
Xydx4SanWZbT5zUdxIxOjhmRd9NkpT3LmepYkQEDVsREJyqqpALYo61oxmtG+FOY
PpwjuptQZqaWwbnFOI/ep5c9JIWpe184SXkQhaAF8HSR/5xK1KikJVAGVrGppAcf
CquDKZpbaPlfN2d4G4RuKgD2HGn6DsTm/bqoN3z0wP+OPxXwjQoHRhqq5J57jplY
Lfcv7GY19V6IbU4M+LK+GYVDgl0XD/7dOuAuJ8hXqX/wopnZs2Faapc42xdMSlDs
zRkMQhXwzc1DAZmYNgir3SmPPo+9YfOZo4f9qFJJi2SsQ6YxICbtvLzBFXVCCrb6
4dVpEQw5ObASXFUOUDNMw0mSopIbynKJdqJrEOTi4PnMzppdeF88JRnWv0cjE2SO
vtJV1q7brP88GmJ2uLNAOGK/3n6lytacSr6ShjMlnRo98I1Z46jAb8O87edTfd1m
M5QykxwrDuf5onQR7f3gEWMEOq2iSnXhtwODMDgn10CNfBZwmLyq44JctL+5SLl+
73TPxdBysu9dYEbJ11yJU1tgcXuGZdq3+zZai77ItUYo7zffxkr8ZClpd+bOvPf9
R7R2hYREjqzyQlhC4Bk5drlqa6wIbnVrhvGydtTeyTumaGkuddVNY12uuCw/eXjc
swWN8Noy9aqpBd2LYf5U7H9b2YGWo3XLI9F3vOi3teE3iEPDwtzpGV2MJpplysu7
ZI8LzwK/TdNsrC/71qh3XyzQrAtQcmkeQ7P1s5dT1C7RloO/azQ+v11sPY5Ud7qc
4SQ9AciAku6p852l4b8snrvkQ7XCigAWTZ0/SwnCskabrylr1tcvqPen+cw1PrqY
5e+igQ7qV1AKmbbaoTRa+1CELduH2Gc4QeaizwcRMRM3qBFut1asiKkCCjeTcZ+A
i1v/FYz7IljgT7zhC+oP3yBNFk08DNU6Aojm2N6lgx9HNoTEObWFR593vYd/shpo
QpI/CA+2aOy5dW1pswDGm/rXYdo10zQEjBAyRWBhDE5Z1uFJ1yNL0vx9/BIiubsU
efLsYZu/t7usLoLdxhbRkiQFP2lCq6K4ty69Fc09QVAMGqecWYyUQSc25QGkkHzr
+WvNu3OJyESNUhrBUl9B/V7cJHB2DbyiHeXv9Ms2Ot0CaI20xYReqjTrD8L/PI86
qE1qcycBEpgJu1P+y55iLQfTr5TyF3vF/cSrmUQWJMGXrlwamwiOk6C4fNMedzZV
XV9zDPvFrypYVKZuZK/v60AD/iw3ox9HW3YzRKiZIH2cVxUMXmfDDxxVMiDiX20I
oBE0gWrVOId0VuungU9+KX/2kDuap9bJ1RsEdDyOdb9ZBYLtYzxD612ivxhmV4V4
VZ0MvnPgOc80gZwtA366b+y36EHwJnMi/j6IW0/dnLlpI7c4jq7Sc7CMQeMQrxyc
vzDhlhsONny7PCyRHdX8Lp7965SxQKcRQm2uq9jI4/EPVR4c557bC7/hbZty2TUl
OcsX+/t7C6pmvam5d6r3e2llEJmJ7oLubY8YshFDRQDH2PXmURoXns8a/UiVxKAR
beW2e6GVeYjbDpSfna/68L2ZZO5cQcdujKqOWQHluVqVPulGurI/Ka02zsMRWKCK
FJKhZaWSB4x0A6tcpQVyODBls6oGORH8a9YSzTjuNBM5JSytlrVMB6apyO+T7DSr
mCzqZ8+C+/R9sY4hXzGalCbnp8347Ek+0u9p0rcDByEblyVohoix1tZe8nqVjqHp
O0Fc8JO1665jIly/hQrJHxJcnA3OaBpb6lNFA7VJxrwsfSRNbCtkqmJlvsZlK9LW
zOpAsI3xgS7jxv9klpzDBMbLDwYxTnc5KFeS6wj+6NFswz6W1bM42TrF+ptwq5yF
KI7e6J95SsP1bLkH+NUqm+oXjJFFLM0m9977wH2JAREuPzREkGcOY0hGhFy6HsZ8
JjO5nugMPn+gQP30H7g4bpjr55+sjsQU5e4B5/sXR1nydSDXuW/Ocd0NMRdmOxfx
LCCr7FzKQ8TKet1Z0SID8qANDfIz5IHq1UEzxh9kiGvexUA7eNnsdkHJrq41NE5c
mEBWHtFHaBI1V3b7XoYAInSE5EbngD5y9R879TqLZRDMGUMRku3ZvaCE1HMxLC3c
nTZTaDxBq2cItrjlxl7ag6tWStn+Y18pph29itTfkIQsK3aPMxzbVxLK7gl7J7Zd
p8tAQ6mp4JqmsGlYBtD4UoIKMP/bAJqMPahaQYy37Ly5iv9wCZlYi/XtIh9jnnDo
byjqtzq7J9oyjOr04rwNDbstOxLuOBHfhseT9jGUWG4CWQNX71XpwPGaA23L8lra
OvEnFBWcxfAy3FriV7b8W8HmlwVBtJAFvSkXe1HkDCYrAYqid2Msl1XIQ9OWMAld
jbScu9r0291wUuQU+y4E7tcHYPTJ54rlvJEfqlju92Ow6QPz2ut5nLRfV1+LXOS2
GC31aA23zDuUtn7McgcQtcBPm9tbPaPv5C1piqUcwSearoW8ebazACfAzbhTRmiQ
nP1DzmzJ5SlZAf4B7gKbh319BaBM+S23kRNcgL2agn78H56ZSriXn09jsypu7o4G
XKRwkOQ3MZF3wHdy5Pqy882K/g7Vb3Q/bQSitRDR8Wxb+mWjy0JiduZdKrzf+lpn
Bm2xwUm4R6wceUErqAWN/fd4ChtKMKpEj2B/N7myDmERVMxfgGNg81EyQqROIx9i
xruec5JgcCtxnoLSaQp7mZHhLSXXWoyqwl5/Bs2g/juTM01+IO4LEoePaJYkw/Nk
C/nGKGUdASyLgN+HJiksHaMHNtp8VR1m4zlZOWgyFtXgAG4VnvXxUTAFFJtoNTBl
Jq1rv3DAVWamVu8tdbFuuQcXq74udznx/VPXuhIE1Rrvj53wgiQOxgrKAyq6TbZj
9KXuskOJjjlGQH8c6Yq3Gx9PspaB188OlfNKPS4/ZyZETFZgAbErq7jFzt1Zn+4O
YIwbH1o7iWlmiatKS23PWwt6uhe+uXXBBXucS8agpHn+DLYbPTrli1qzSBpQmU9O
BEZYqHuBvm82KmtIczmzHG9chFv0li6CE41bwSp1mTyNS5cw51SFs2hJptMIfacR
oEdPABIbYTs4NYEc2NbzPKU0Hc5Jz4170eWyqQZhUxc1+2Yip5hnkydyhQ/6xG2V
i9lFv++ag/SKXpHXbMw0akrD75Tp1M7MV9UuyYqMfSpNijre1SHeg6I7Ej3dvPfI
BadjzKr6Uq65VGjgOwfdXlEcFwsjn/IIQPtKF5p+OMEJ21TsfMOmMvzHdqElr6Cv
03jE1EN81ds+JxL/aE1DsgVeaPCTkQQt6+h7oG5FgobuSp7BQ6XQrSBbGu1IHlHU
y22kHhnSL/K9X8CZydGc15F0cZFrxqo9qCojsHW8EEV4skJNC4nLfejg1hVp7KG8
xqDwb+22dYgtZTXHN8Fk6mW1jXGsy98jIJitfTP/ukyC2awN5agMg0PitGxV5uCB
WJTc61zbKJ7Ms5nwxwZ0WsjuQ6DscimP4OVEo+NJ+hgD3AGbsctW2t0md0FpfDF2
Vp9tcCCVG1SyJbkHC3lYiKcqM+pq/itR1ofii6eBAJGMoQmNMtPqzU1BJfz0l+4q
ORxgu4lFONHwYBV5SyGm/HPp3s8X01mxigIGuge6MdX6Ul9hxOq2leIX6r3V176g
GTkkbCIaHM2aBiEjy9J5a7owWhDBVgnbRKwchsFQWly7ldxEznyff7IJPSlm2rrJ
ZVY49x2woS8lXJpYmHFcnRW1hc8Wg1fQ5HsJnokAZKzFk70fMGCYsgfzykC+9vcy
lM0J3kVoBn7bvAsiEQ1hCS9CYQ+Vi5/OOJJFccljd0gAgcfQT9mbnQsKBM0YmayK
aX3H0Cp3E3h1obRUwYr/o9JRK7iFSQsOagpmX3vJPlolLwWTeIy8v2Lk1cqMIR5y
23kr6+oZk+NZ1+nF0BM57PYXfGFpvEDIZHR3i42K03Dr7m9zRbXZD7RxSuAQbEpH
mC30hEWLttgO4wGntJxUq/A0gdw09XEgVzQQJWjUSGj38U1kQcEBrfMRjD/oWoGY
yRPTVgnf4QyAbL7OrHACj/3TnrvVwp/Dv4PTwx+Xx9g8dWmc9dgPgMQ77CA/3I3J
yVJNQK0smM3eI+AneCxp84ay7MtNSyzQ3zuEjkgovgJGLktkQBYQV+VEa4CIaNtZ
XQJQE6YBzhrXAfRbtE0dA55wB0fxNas1gZIBR2jgd+XnnQ7Wr3RLro+QRZJ7nphN
knHVMxGlTpd3b/PB7li/YoE7eu41nWw+MOmRLrMz2K3g0o99GdX/u9f4cfSwttl6
36/Ov2j7zXGx1LxpsUXDt3ajNEphu0FiweI3dKuzzGCc2OhBT1zrFxyDTuyLclkO
8b4dvHlh12p/ojAYip6aglp3/ThPTIMqxzPrG7UrsgMJA/wjxGWGrcIu4hGmbHGj
sWS1vJDdf0k3Z3KREy53iOYPQ6s4te96rWXps55Qv5IM5Apf6B04Fjv9c2vrkUW4
4uR4t1tzJvBQnf/WzVI6eVrllupzyvcLT8XOHWoVdlv0J8Z9BrnFBkN4JQLiw9dF
pf9Zdfc/37XloiBLD24tktyfCopQflfaQmTPeLjnzZnWRLim7CXy9R4kU2Oc7ZPR
UloLcT5voRE2q3igEgkX0pWDdyuBpKI5JZoO4ojFvg6nOj78s1pn8TQQ+1iopxhy
qupveB4vezPejUf9XYdB5OhERs/q2oJVbA4g0eNaE3llY6kqH2GL1YsuIm0vQou6
YvkrB3NDzj9IOLI/uir1wOaHJDMBAwXBGTcZjeCALSuqHnHInU2cOO5xf2QHDVXy
RtPeCE/vkmcLsqiZ08pc98ZKW9i+1f6A7AwHZb6SQbSk4Euyq5TLCPIeTLMQa5a+
unbr7WsU+6hDAfoBXOfI0pngRJ+7p3aY6KI11jHQDTYlqRPJzeHgFcj0i2lFWrQx
9MMbExUfga2pUh9EYyjGwzXQMA8ySwz9T/17gcZF35zK7jaUiOOKFpER9r8bz7uK
/ivShKCgdK6O0AyIOnfyVyAEwNLax7TWV2ivXcvcV32fBNFJwjt8a//uKPOtGxYh
kavYtkzE3bIK/okeXgX+Ud7zctDtpSF2JBcyoaee7J3DUXem9aCI0fUYIOoSqbEK
XrpDF6rWvvU13E8BABwT9aK8+52QBZntUlggSi0pYabnWo63/3Byp7qNyZrsRqOM
q39ShtKf3vmsHq/zGEMMv7n3YgveUJBVhDE8A2Gg3kUqQU4zEgTOcmExXT58TGw/
8n0TmO8ZA4/LAtD1nxD4GyAN6FICvmrUY0jYeRBwB53RcrlK/Mf6BDeEmxoDqnba
dtppCcQWkL+ozpWCF4NGEU4Qy0vmvGIPZwpElGczgqEg9i68m0JIdOZxO2ahyOS8
k3hkqRvsmEHU3KldHjJBYfky7Fjx+yybyk0i2ybGgFXNF+baS0qg57vVT4cOKmSp
WYC8JxoDNmSSQ/iCjilKhcvIkP0jbgkwRehOLwv2yeVtLel+vXYZP8W8rqN0WFgq
6Te5jp9+dzEJAyPHtvaWjOCCk59NueElihdfRAEbgDYiDNdmfPMgEWBYz/x8fLp5
AFp/xYDqAkc8E/tdAcimS8SKmRfvxacMz6DQ+ogJd/tafQfkdf4gLpQ6hfFsXDQ+
C9cmIwA6ovwRc2Tfo4Y9IwvNSZ5Jlw1JZe0sWmscnSQvzYIn3W6puCAZDSwBudAk
8mUNxjt/b9E/U9qAgSh6WFRLW90Hac5BMDN951U3e3a6eqgsJ/thX4Oqxk88fJt6
f9g5aqx8bf9BkOm6Do+DADBbQ1Vn5E7UJOJ9WoRWv7yO9A0ZTLVIqnPXtl39j/9k
B7Ijdo2VdNjhBkd6fpUXHa/cew75K63s3KkR6QG9c3AGZINVeAxFOwvZaIFgD4Xs
Agz1/VYPb7ufTl4ja+WDVgMR1fT3dVIKddUkCS1hsOGMv5E96HIDMZAqfjCCSTIm
NHrawE0XK4J2BP+T9+oerabZ699IkCM9f5c08zB0RaeFmwGMzJEwiWosDASkeTXy
oTnxgJlpk3R9KXUGZVyfNsXDLHqK5B5V/nkMDPpyypOOsUKSEyeu6T2vxa7NAY9f
7MRh1wOQfmbtodRY1c0GJGCOX4MKPU13t01eA3CuJzlhsFvtTxUcOJn82Snul5bS
N6JIafuUvC1mD1B9uwfp258nxOh2E9j6yFtvhgl1wq79PVfoKDZaH6uwCnd+vslH
ArLahIqGX0pfB4xdbgRKrkX9nKZsUlQgNV2/H8aHdDHca7PH/Fy3/yufendM4yVl
5Ks7wHAj5U6YvND5X4p83wjjP/uV6dgk3Po56TpoafeS/Wx+nARZ3dD0vwXGMebc
nl8TUrIU5g9CaDlHwkCueio3n3tFuwIq0a5BILlju1v4Ha+6FCOJ3XqKQcLTXMzF
Em5a0cqMJEtEDEUa+lCahVPFXPkapWtubnZXcT4wRaHGBmp1H12fRHhkMOt/ejtz
sBNb/zJp2svVaB60Ds8qPOSYVLcwa5RR0C365KGeRcLuO/54dRvCnsnI4Dj2ZF/r
zUoV7pzASwGGp9XUvOrJtaW47QAlcNTAp1XNFtbRhNcIzdwwMtHh+3g1IXTBvML2
o7S0QfvU7A2R7A/kPoqpOgTsLSAND7LrEkR5FqWzyNhU2H3INBaDbufr+ALgLn64
VXxZm7s6koHFtzMKCrDp1thhQNIrvpo7Cxwyo9gF9LQMximyDQaQVSX+NF7+3FaV
B360pQNR+cpX4xWwxvmaXWHS6wc0zNkwp0MWmZb7IY2e0t36U5WVpl6UkXF4F1Pu
V/uvOmVXTC8t0e95I/i13J6KRercsPG1Eji+vbRHK1YtizzVnjiv+22TJJjVIyoC
SZoJ4ie8Yf9QX0NhoAw58Zqmx9iiTjHbbPmAHRoaeJAu4011u5D00g3z95uFYy5N
2Wz5UGYCV76gcylJbfxrGnTiCwKQuipsLNnhf2ipX/2WQNzKAO2rurYwfipyoyoo
A+qm05Aax8Ic2CSMI3ktDWGE+0uxH4hKE487LNpGDvsZ5JrUIH5potWXjuY5sDLk
ZGcVpW+YsplkcfStrrjL4AGeSCaqwN67Mdr4EXC9Da7mQjxXdsPDZuHFwx/HzNzG
485XiK3pIcPYVorH377hs2nP3rt6jOLXu+WLfVAjUR0x8aYyyBa6rKpWi0KXkQqA
AMRoNWKMZyomItD7/qEYC7EwxPQWNJx8+25YE/3mX0hXROWVXupOY867xtMR0Yks
PInZNirZtKSNEQk6FLyGlXs6LSLbbkUsIBkUL0nGFc37r2u+58xVMwxT8ClQbGDl
8ufi1mNa4eenGUFqTIux+R5SwnKSdN0f9Xu0/ayjTm5BAqeM5QYvMGCNwoYEQZFw
f2N0xmZTypGjBucUkB6rNMEwElgRZi8C52u7lwXXvT6y1M0vU5Tdk2bO/BH/fLgE
xwDO9FsUGJIrbN0MvMZ15LOYN4vCPOuwnQBUz+mNYkkXidj1h4Rfs2umTPT29CvC
B/6MnqrUvjAmkefTBUfb0X1uhvCcAD8KwJ/VXmJmo9veh8sHsyUCM6AYWrGYPcYq
pq8Ik1tk/yMQcrUC4uXo9v5/LIqAS1HUxjkx1A1zBuxVDX7ytPhzYwvej4boqhg8
8PqO/JTKaDBEGyWffxcLBP5M5nld+T3XvE6EFkvOZ2worJpSb+EpiPc3PK0xqpTT
3Xn+kensZP1EP6F9QtRh5lEV87YkXGa0KHb42NQvcfHZqnTVnJily7CwAdg6J8JJ
opfyt7llFqulnnuKb1QwuKDN3onlIB0F69p0RtbUKRvWSxNdDZdcRgo1j1Wgtp6N
sInb6PAJ5At8vR4bu5ywKmqgw9zN+N5NJfBo+9jbpApoeLigU8sClxTbexfLJmBH
B8oNfOjJ8vMBS/4LhHdEvujMKVAmuYWkYFbghNAlC0zgYqe70I8cUjuK2qqVY4QI
6Jv9uVfxZDfYvKQuIX4BW8VGlB6UQFM7ksFKprlkEi/umek5GhiF4wld+lho08m4
U8ZRcUK6oXEvMllTTPxOFIhsnRggQxkomesNL4PXwYqJX4pQ8iUHDAr+i88sbCdj
nKaFn9v6MjMEl+ic8/kZzfe8PSZSac1oqvTNs1FKjr2EUXUy6m9PLyRhBkxrxVIe
M9J3q4aj3d8BKvw4U/rlBl2THJjWvDfYfPt/j82LEmg0WGRLBnTlcMvkpjHwicPo
X/Nt69G7HR+umK5tNO9FyLOwWeA8ilEZnUdREIPZvaECmdYZAp90gACYl0Qp0cRU
1wAfbWaPu2TnKvLx98sCbzm00SIEFe8NhJXBCDiQLCn6if3oj2lQyQyAZCuCD/i7
Dd9BSx6BM6BlIX5dnPjj/SKummIWc6THsDYdIldnD2lfCWPA6cyND5gK+tJp1YrY
269pp/PeezT9pasyoga01UB1+aTVhEhi0eDEeKYHnf7UDD6Lmio+sJ4RU6TdP5QZ
JSodVu3Tc2u1qeRE/aEkRBuJ55TwXSUCKo6QG3kOJGhSL0AqwX5VYmr4kn+CblEY
prxSS7Kw8s6qfdKJFrPLQFnoHKfwvbqEzWKOEzhFwLVcaBVffrzAFioTK/56J+8v
61ZiySMnJoy2ESZdXRb/VlEOjw46oSrzsG9tDyooZ+lb+zNsPaNYEyCNtJJYicd/
d4jewhDBijzdVeQ6/6Q8KaEbgOch1eCi5ZufmYquuRnYoAe3UjRj3PEu75ICxTCt
5PDcacn2860Q7CqM5mhJW0scqpjab/44XMuhcich1qve7IeRPwoCxWjE5K92oOOe
y6k2jCKpI9lCjigblMvcffNlA/xB67bwqHy5uMMfSLyGLgSkR55vLVsZCRpK2FhM
snA37hdxAPCNQIYxfevYA0LEwCzmSwwhrx5esHvl91Pvdr/AqS9mjPmKjkOVFIV+
UrMCoZu8qdlZLysI51/qy+pFY6Qhm+9PEIkU1VmRqXAMQ9fk5uD7pcSqEPiQCkh6
mnIr32vIT/9vPAMhUsgBHaCZOv11oaLOwIT4pncKBxQlBzFHeIyTVBYBl3Lh34LH
D+/8N7DEFWzgj9hQfNTzPFQl9jaYd1OX7nWeJToqZsJ3oAblL7JBqFvZbLFIOv9p
56NUVXk7Ij42RSGfxhcDlPl6Xa2o8VnRehACe+Pi+f85ps8jv6O4a4m2TEwD7KnQ
U3oiMFuhTHUPs/GXgYX/AGrWKJl2NiBNPZ8m43qBiG+PJCZguySvL9jYZOpVW2/c
CAfJkBL2oRpXpcu8tJFv0jmZuCryNrHoZtGTYclPmmqKS3FrSXRNyNDktXm5sxqK
1iBq3YuWKer50QxGfShmJbSa/axqdopfCJZQYFFKmkiGsUGvhjNjK5Ua7cWDh982
Bz5e6N+xhfnn5so/XKAxajlgtN9Kt5IWUnFMDOH1oPeI33swgvzi5pTZ5ayHiujE
LpyrFsvXjx4G5euAnQo+aaAjjqm3zMf4/R55MyEi+xQCaRSSizy7P76enEy3Z6Iu
R82YPYv+fJvMnAtgSwyNrVWDFmsIkRQrghQqa/HtEUQt2iwMOwUvSSVbTm2khIIA
KwxxVn4hq55U4QHd8jvVSbe6Yde76FNGSIO0eJi2KsP2CYpX5Zj3hzU9vLpSE802
e7yZH3gAPCPpUrfPP039m8PFY8OixGSwGVH85T8xUy/FLaAuFoDqsJUe+VYdR5bc
FaHEVe2EOdHN5xKAdqUuaqgGWBzH5UxAYiAoRX9/bzq0OQt6e+2eXVczOaIV7cgZ
+sQrQa+ljlPK6TRnYS485mlaDhY2wRRFylE94bkWACUYa0iAv0bEc4vKvQA/Gncr
O6I5Y+SIWG4ZH8z9xvDMP5IVjWXddV8wsGyo/62j8ouOXMfUmuVKaMoIkqtvgfo7
75yu2yhOmohosxVh19npWXfmIllTrRaeKZFDFiPPlJLpX2qobNe33N1FKrb/R55H
52YpPfD8iSp/eaaAVQb0qMZhFCR762Sl3wkax01UPWvYOcmIT/ypn2A1496tnmA3
HiDpfovhwcHdmh6BHpb+rhm6q/mI1SqMvmiM5ZNsIu44+YhGT5xZNnUEkI1icj+j
h5AaWqYvqP2zY1vlo3xrI5jCafx7DAJeHADxnm2Qwbw/c5tIW+tI992yJw4Or3iN
cX7/77WxsPRmePwyow/s1StHBvkltHnwSjWuZU48zQz2V/WRODmjsOCTOsAkJeMp
aHXdLK2bUPA3QXCvhhHuU7ped28nxclTaNoE4mXVsAYyNfKWPzkB8U7x98BVZRub
2Z2RfgDA/H5/ZIuWHhOdciltb2mE+zEWsMjAfi9IUTT9oG9/p/DXO/I9ZHtErmjH
OFVC3jShkKqj53Xp69pMNnhdK+xmSNRx62+xcTBbNUAfwXFz4WXNXw0bskgsDkN5
dg0xsNpkgtck5O7pxazheGAKabQvMIAOvhbD4htdwuUU+Jgj1b7Pw+dvb/rbE4VS
iro++h/O+prnbgBxryjh58VGIR/7E/RVt2LMeHPjWfwsS3r6hlPV8oeOKrx004O2
Taxi/WAg0Ltq5+k1mmsTTv2ky9qG7DpjtpOF3lPEzQVBj0q/7wWkrSMfHuu+lV+D
uc/wfFdZP8cLzhSZPppPQ5nmz6JnpxB0/Ft2YcfSu7ZPeuyzur26ipxemk4JnnFF
6hp/a6GrxP24nw7tLcEg6dTBxLG769XZaApFvHhLE788jnIh/U6OmgBQlJKskHqW
sNpQz7ryNGGV+vN0hlQS9sKi79iXseP+3eId7hhpkuFbUXB/E3dV6Ka2y6NlwduO
uuBuA4o6wO3jAUHX/9NoLTXGf2LwI/w3RDs+l/dfHKRsbPPBzEqic8g3oXLheN3d
lKHJfkA6/wcxk3OOp108hjvPS/gcALGP1QFlXZ3o+0wg/72DCJB2Uz9zsRjCJ0R+
CVnuzpMAOR8CbZhPBNk5wXa0Z7AKYh8Df8xZUAmX4+hoOZjtpAMV5ujgJGmp1y0i
Ri3svhPm0rabDC20a5SVI71d8GNprP2Cdk+t6hl6HQhQDGRcjHfX6FAHXoRooK6W
W4xFg6IMnPCHUs7sQKpwStyAal5Yx4J7gmA+wbBKH4d3ejbpOI9jr7w5TsezCHcA
9z3/N8vWSqnPCyPm6kLkFaW7JVHSFd8FJlUUHiH+U3BXyKsrm60fP6a92lTQoFcZ
x75+Lo2fbu1XWaBIjOBEk6KrAFal0uvPEm9TFb5+Vniy1og9LlRkOt56r3MPNFcW
zpEX0Oofu8LXcY7/6FRzaCPtZrw3nennxfxpUZ9yWeYKc4P2a+X0/sch+lY+9sLH
rUARpWZpi8H3Tv2rbFg9/cc2gv++2Lbj9j5PLF1cZOP74ahvtNvKUsvufJw0IjdV
ogI+f8sXuoSQGazefgz13khfjKe2kRz+rsSMHyxRiVOve3uoLO219jNDkQSKIjdK
+3hWy4++rghsuFWQSG1dF69868ho/OqT0QLqDPYT8V/2KEfVqw7HuaXlWV/VLPUh
aqhM9MfVthQSdU4vLqkp/oiUwBJiVdU5IuWQQJbVxa7mZZ+MpOdLwxIMRRyZefCj
5fIPxGvyw5CeVptpnOi9H1V5HvKwMwqsEsLPmcAuTAurNaURW4kRfLs9C3PE1TNr
3keFdXXxpvcZSYs0fLsHMy8tx79SHJEIrnPfTYeuByLQTD67QlXwpp3vRLB166rF
rPptXztzkVOD5thVSyNITSvro5K9TJXTreD86uPnEIp/QRUsO5LPMXDKbazKZwU2
W9ENKp5XEZfd10zp1rTulfry7mqpHxFpQedvrDcUS535ctagfoxOPWhP3f5C+3M8
7b5p922FgD5azHTvHF4lasZJEKFf3Q9Ct8b//07aBvoQJXF7LUsieriEqv0b2SiY
EmiNXXLAMc4lMQ+1OyOIfUfvBk+wbN85yoWfA+BYfSLSv3oGJGD/C64Hl/iatAeu
sEnlLWMyRhta7Ne8a05wzk35FC65lIo4Wdeiui7zRhJ/ebB5tFMLN61kTaIf99tA
8Y/5cTRNynsXd85e9B3uPtFgfofpl4VJ4tfy7rh/90f7vLrKh3GduewutwOQB4QA
tNFoAPgSy6jYEgxkoomAIeBcFYO4lRnrCk4Q9KOUuhQqCXMjHn1qxz8kqBlZJgRm
eet2/Qs+Ait7ut20rKgFSACTZMxypMUC78A1AqFOTXVZDtvIfuqo9FRlewDxPJin
RSVc0VxFVM/d7GYDunkt2uicqLaqQHlsPKlVxhI9OtCWHzo3+9IEKJc+F/JDqmty
3V2aTw2mxxZ9bV70svFG3gR+34/n2ofYIB7tgJut7v4bPFuPL+9Gc4TPUH60kZg1
38WBFvhcLc8E35QWbIt6JvjUbNRMNJsGQ3aBRXA+fP9dR5a+KzTDWDW+9xJ8paZm
zeyvybq2NZFC8nubmO9MG1A2YmkvRsUxrX5NU/A4UwJk8Z4jVEi4sdmfts0chIO1
G71QkHa9KoUGp85QHvTNjPad/kfqEErEw9nXSmlcnGFHqiFyWu3ICkjKxeMU2lg9
zdCYffG+hKYzZ04oD//6ysVGo6jIhvMf5qNp4+qlP/sZ24m/6CqIwqCd/ky7Rh7L
c/3pjDzfc4dQUu7lXqOEbdhpgDuEYMcYebc3dokK43wzY2IM7EG9Ay/upu2yGalP
up2ck4UepPSu7TK3jNyu+7+nTE6xmu5Iikl4IgiQhDOQhVKVCE7jngSUdNk33R4H
tafMV3U+AYcL20D1FtAs4ROeioT+BiKWFvgRVa0QcekK35ZLIcPBJ3wthA9ISuIX
pHGehKb4PyPwp7pSqBFLylS0RHsJTHvjDZ8sl+c8DLvSOY8ksYP9u0yftfLuo7Za
mmrpAzxkn+3VA/UHSSotkMoVkpbMt7aIcz0L4cLpQqzuhB0guXOWrtgoExzBROUr
PvLgvuwtqLgDqJJVG9dITII5wIsn3DxfZqK7cvmjhL0kyar6FPIiUiK1OOk13sbT
M+0+IKjcEKoCqj9zAtVtzDyUCJsHzdeAcudDw32W6sedswOKYvlywo7Yx88uybUA
lgILYbE1Z8Q8RSTq2xzF6Jq1Nv+ZS8N1RIoUZMlWXt9qpf07jtjdB1a6C7ocg/Bq
itwONOHGyS8Ozq6/PyFXLNigoDvE8U0RN6y0wtmDnR2MDl4534XnXn4taR/awXPU
Gx0LBsP6ly5BbLWkhDmIB5W6CE2Of0x5WOyFvJimJIe12fJBF94ROJKQMzy4QYS/
eFKQqSdTp44wIIPieX8oBs+iiebF9NsfDlIrIYyDk/n2CksTZnpxxTncnN6gTGj8
Q8QnDKRpt5P6COa/mBGfURy9YiDEPL1MGW5i+Dnseue2Twt8MKfonxsRuim00aqE
QVuXGqB0qH4C9ZdYWH9qHDIj6F6heKg7lYtDdMnIW0GKYACvi+9HBtPc2QMmEQ/e
ooi5UiYOVZZKeRvZs8koLJTXA5W32DpJr1t7bIgZp2EsF2caM2QCYYvnDxsNLnUm
6BNNe0fl8hiiKYAd6AWMrV6wx00mw0JQbMtRGEFdxYy7s5e6fkUIfjtFNICl0Qxi
BVbhltmCl5U8b5OVwIFnJUexZssxDiyIT5iYb5G4LElHhRB0DDshM5qMf2tKnnbD
lUr9MWGwKFpE+RMnl68kvzAXUp4fP5P/aq6jJcwSKIfKddZKSXMziVEzPBf1bjYF
do/BWTvXte+yT6po31tupCVlg2XSWySNuftH9MibVPl9TX1rTTaCNOUyHnEHHdsa
43raf0xaLWw5ScMJkKFItyslP7rl691c0r08t1gNIBO0DL2eIf910TZPvyCP35My
kwKzB39PbVUC9yfuO/Ly5xtF1AD6QtBD/iyJ5589fjmw/a8DsR6FlZwyKb+C+RTI
04/YtVcYJBXo4Jl3WHpEf4c0WGsSEEtzvhYpbZupXEcZKcTM5/V2IL9FM41iVxsl
clzeoeRsgak+uVzWi/6VKAFPXD4RWz5FT+mlm7TUMCjLzsWKW4mYbufim8QudqZG
f4HPx0iqv7SOgBgKOOo/VEpm6jR0/4mrwXoEtjMQxYdsGhTCYlAQzCyBqxKzz2Cf
4N4VL5qN3uqdV6G21fua+upcTZo302Z6mkCO5QTv2RznvlAKuALGPMIAGvtcDBy0
SkXkxXqWVkRwFjtSbO20taoKU17Q1Q/K8UEI6yXd2aIwmBO4G30Z+ef17QgqNubx
JpYR3UTr5+7RqBWCQ+qOpGluvq82/YPwM+B/k7EZWyWBQe5Zd/VdcX7l8IcVg602
8hxiCqMOCLVJvPPt8d7fWXOrmXOuQph0Q0+bCX/U6KNjJlUQ1wsrPxox/AdPkjSV
vqOpWFb0I5Lxy8WmwdMHbJnbZQW60SjG1W8CQUViiiaksjrFt5gbjILcR7nbhtLz
EdSyKnk4J8Xj39t4aZnE1PMi3TNK4CRUeTL5eu9nRVfaUnz4ikRW19Y0heElPTI2
i8ySS/R8F+grZINWG8fj0kKWYH+fzDa5z9IAl2zAplTCxXhMMlCjJHN2cb3vlr4R
s7UTIQy1NopwDV5jsHloUBU1KnLEUs4wmfUBnbVAanBcW+egW4Mex3fQsqwmDWVC
pkdcpaBnVv+YlUDXjnLjG+ND087cdH/3PS1ClDA6Bar2RH7Ny5Em5Xr60tbEhoJH
hAdXnsJgEfsu2mnorAcwahx91lnjrVIycCgHndhmHSXvTSn+S6C0uDjfiFr/zQau
cCKYPQVII+Yy7sd3mLzf+ZursJx3mUsht+Yp3hYRu2Jg2Z1dD9q9TWmGfHhUAYQ0
VTCiRj5MQirt+najZS99mwv/urqGFvx0tCLeVMpsNUMpHx+wwl2yUXsR9VDvpcFW
QSm+NZwBWASbonY9mRSz22Iv2nJPlulYOPvjNrUI0qaIqwb07e2yJz6bTpjdb02d
VpJiI4wF6MWVnrcMAS14CkhgqKYkDXpYykI8U2yR5uZ2z7cSRHFwUT+TAAWGPPRm
M/n3oxBblvyRY1E9E2NStzIoAKM8eC+ewiGifx/+A37ZvluWkA53Fhc9x9xRmw1d
OWGhELsI1r3sjadPIkXLDz0YM19UBY/h2z9XZ5dUOGGc78NUIohQSbO9K3XeEddv
knT+m/VTB1oCT4kJ476b9PX96ru5Lb5LA+I7tCI7GVso/7T1OGrYvYQPrZThMmFw
dpTyIs9UIjLGkgUgEC2XjuXulck0rOGqZGN8goKNfKY9rYDl4sis70tkgRsn+HF8
3GShW7wCWEiSyNU2GxO0Kkf2kzFNJVW2+AzXS1XUlY7uxHnCRnogkQkPtYt7UzO5
pcFblLAJoH4c8SQDCvkxfAs80O09qs5ERXBvmpXPdIq9WjNbkrJtDWo0ecuB1fb5
h+u4tkKpt2Yyn1WC9OjOFds/bnIxSxWYdqZEBgoJi72ZtcEopAn7qBU62viANzDg
u51IRHTr2x4UKS/hE0TzxBucbV1D2NpPmv7xukpV9oeQmnNnddh73O4rX8Z0QGDR
9tCtzeZCqpldoed2z3pyyTDM5lL/OHGwIRKZbPWkekbXaNSXq8uiq+1fPt60cikF
AqgZh86uHtbXL2/08o0SK/HYbDWItNN7HmRJsZnn5yB/g7FMAFWhFKeH9NwmUEt6
tbfaLfAq6DG6V8SxbJRidoO0Wy5gZDHlCVGM2PPAsLcHoyBrFwjGSyvle4nIO+wb
XNDZwXgLCCPnahbquXCnwFPaOv6dQT4C9PzPCiqW/3hDqE8dj4eJWSfVBw+vUyG8
oUwKmjQN3w+dLdEBJG2cRO6hN7QfXpZW/NhGuQUUz9ZRKeYucLnQRluFXT3nIQ6b
MljFuBIw+CKamrb6n2Jig1I+CstIFQRaKj6I8f9ZkHByBhg2CGC8wJWTPk15TtFm
XfO1m0OjIGAW6vcdxgIFL8DEt1c4Lww/q2M/RKmbBYZRbILqWEUmUTcO5ewpwrcK
nXaSoIhwjcIHA19BGwMu5DDc8RKF4fmaK4pi3UEUgj0f7Tre+5x7MZIGOwa+bUFL
3NU9+2g+kfzF3d5Xa+KnNHjx422ie/pz+erzVXsNhJSeBk2NFt++e6cIPX7H5tcE
63GID2kpvkyTlMQ6WP4ZWYf9b/8ETqKxj7TeFxFwXmhlwjb0lkvxhYDmW3tkSuVB
xYe0qafnm1X7q2/W3cQfl5abhn3PUFg+RrR0GigV3H85nXeva+y9TXJk9tZr2sCI
54crOA9HTG3Wf0ldgA7H0aS1gZv00hqvY9NTrknBYZh6A9KSWbCHoZnl4PFc8S3w
BtcJOSGZDvOd61uZnWlqJ1YjN0Xu93BIKD8jqLZ3PzUd0wtptIll8gzCIhfJasQX
PAPjxGSzEBgFaN1RTPr4mFtYCz3fMjD7RL/hYaDsiNw6qwuZ+Kx0d/Q7bA5/kjkH
AYUV7ficYEJsZ8rmA5zf4d+CX1QW3LAIcA6c/UjBKsc5B6tZunAI++iDrB8R6uQX
TZnrUzl4Bwc/eRX1ItfK3H6j24iKc0g0z4m2JM0Zy0hRBemwb5Rk6anh+C3wul9f
TNmdgjEmRJdpzBJ2sH4EOTp0A8mli7wXX1oEfBwbdzdLwm21IsILsIdMopXb+H+/
6uUrMhxsTAWLfLdeI+mVjRKicaz4SKxKrDk+sTWmmCIY1iJQv0PwM5QovoxtHuKH
of8ymPg4POEFPk65r2HSydhUOTXeNIZkgcdEH/fJ1cBoK4RqF+/krTLh8z8N4hKK
rmEt4Kzm5f9sJPrZbjeZtVK1/DS0SRlwRF4DFhKIx1pANVNb2ZA4rg0+XTHJ3xJi
u2jv0VrRjAWmqkoOFMzv/auXvSLICCT3EPPXMwH7A/+UxhCRRvJJYhCXL9MIQWAy
3z24O5Ivn8sDV4xUx2zCxEHi1Rv3CgXgDhQzuW07LGlh49CKYOyA7Fe+Bs7QkRYT
3tpsL9wINOstpniiQV88JHA2JHdixkBJrP+v3PRL59nXA8jo+2S8fF6v/PaPY5qV
OSwIoJemt457tOrPgYQnYIb9aZzX/nya3GuZ0hh6ntC6WEme+THh1pdjrqVNpOLJ
cIXD71X0infzld3AsNb5c+ltxxAHhVrl3cnIKQdk4j3KWjIy7NwHP+mMQ5hncwdb
zODFZEdjS9yLsldlRFJSYLMCfbH+cQcK6PAKS+ZMpd9rgxrv18faowfLjbYHH2gD
Hd2WjSr0uy3QHTwWospl52Ra0/eseRiGalWVJKpMjacuS2rLrES2SwyuNIQn1kDk
gJJ4o1uTKrQIYD2LiX9KuUUkFyA0udB2j/0CDMPY6jBU7SWhAWNoqJJe5w689l3c
vkvMlafK4c8YXofPlkAnxmeqMgROJ1OlWKVVgi6zHvroYZmS0eBJgqGKTyUIdBCo
zT60EdLsbmO5mvaiga5FdyH+onpl/0xZqVMSBrUzYGv5fZcRR6jx+7GTAAym3Qlz
actjP7grgQvkHypQ+Wa1K32qI3Xe3ODn0L6koXgnMe0DSrL1ki5VzkwHNzzxixba
69BTWBadrSsN9Z4v0imlYS2Kz29jtsAOj9FRenRMEZ7OhamSA/FIlYoWPgoTrOkF
X3s8LA+C3/bpflZCEdpq7XCFzkvunMxGNnh88Y1OWWIDNS9fs3AIHbXaWFveyhHy
0yZ/DVavj4ysTmKSppicuP6jPvqcLwbINqLOyZp3+EZVK7eBWN6jPP7zI8/OY6P4
FGGFjORr9B7OfNN+rTh/zwghJKbR7m2I1Fs8ULkirlS41ek5fynJyDm/2y33/25z
9k+9MDtizCSfD+MQVAXeBBdIQ0+e4LNgyPYmZbKgS+zGojHLq+cd6MKZPdw95BnZ
TurOrLmx2GqYK/sbCt25XqNTCWNWVwWoqPS2GRLJ5WFGSL2Nq4/25ooOyspmU2B5
JdPLBpaLqPnfU6n1J8KftkEHl/HCf2kknNADmFsz0/zqMPIzoeG8o68COIlHZ8tH
El27nu06GIp/ftjm5kg00XnJc03fg6mAC51kLii64ALgT7ch+iJTdbZEf3N5HRVv
bqsm5s0MlM8VV/ui0Z/kPc5UjQ3oo1wW+qXUjwVXv+LztIq0L+oWsK8tc14+JSsz
N4fZSgzZuhviAsf8vZ9fQWSdDqKbdyIplSW+nPD2LHygI4nCXsXPJP2HNobariyv
x+86jPL/YpHpg8ybnrBE6ZUBFS482BNFLecYMIUYh1cJ9KKosOHJDi2lpVlWzbt1
iLjDodfgu9k8HYV6+leY2Wj/Yos98V1PuWEKmAlvNyCJ95LNGUTTogmDHxlpv4dx
vQ5bnOmfmiBj6CwU7oTa98zuZsJQxxA3DbBDD1/L/AbJdmWvuPwWEleHxRBjp40p
Ho0ni4PBkrRCNGHDMZs+H/FWAxFXvIP7JjyMcYggLc9uTtiXmvgqhtrze150lKsR
iIWsczCi6gxrt2lKAO/0rQt9eWxW5rzS7a27hOLK8cvn9UxdDy4SM1PiHFq3Bjvo
tfLJlNrM8ns5V5sxPoOy+o9/fDdaE//+gxDQWbr4PesdZRo2UqFU9t2MDfFr/NzN
7RTWwyGBniL9OVyqXuGVbgqfuyJ67cIWkMlLbRVVSNFUdM2iE+gtBMaxMVknLgDY
cuBtTfYnw231CFUaH3aMTVI1/yK5mSgL24TNh4JJ7fxA6KxGjPOqpd+dvE3v/QwE
8T0YzajQpBgrBRvhBY+ctsIjLjTXrVDIudjZRfCILFY0T7jwqiJk9jsj7p/B1abe
bun8wqJBaAA2MlvIRWd2oe8TfmN4tOpqupLvSaLcAtrbw2vZgROz7B0Aiil6sf9Y
kQ3+CLFFzCOyswdhI/YgKLIdZW3eVASVhfqBZkZ8LN0ukmwv0+TwgnMDMm4lq0VI
sfRRgtFGxmxLFXlm2bHlAin5itfQeB9QgO+bVPLUp1CC/5Pm+RwFLlCsVAvWcWxy
D9oUHc5ktQN3LyKF6wDqcDV/wbYUMEBRe1yvS10t/dZllFKz8nC1ZJdmBtX8N9O9
TDkTWuO6e2eDL07R5iU4A2g9k/bYb9BbR+NO4PYcLFrufKN8dK16J9NmHwYgCBdv
hUP30I82oUQ/fn+PLhadlVRR0g2YfeiSIS9fAMED29Li6yDC+10gr3d75I1qYuoH
/unYlEYWitKYylgJ9gSJywzkCVp5detwnBD+znxLWzAazH4+ZsMKBNiee4AxoqIt
+VnvHX6Zus5J5G+JydrdJEv7OVT1md1aVg/RDA8zspETyYXTH8LdB9PXrY+PCLes
yaDBOz0hz7dgsAPcuduVDGwA5/6pg5oB8qoS25x1pS8FEUnGE5ACDS762t7bya8n
22bSfZX2dxQC+lw/qEWfP/IVbpKLiruBp1g5U0iJZOlXrDEnxS0ySwh3m0s+c8V5
Jbbgn+pHibP7mHEopeUpOJ5xeGv6xLRGCYmJm6b+iOPITtgNsoW7usE558NKA4EF
qDUV943Jg26ZfgFiFAYo65avhPv+Kp6ABKwRoV0fGtYeRG+QcB87Vqkxy/+okdiF
OOvWl1k04Lrb50TGeL5ifXZcoEZVQzk5WdI6Q4tAHXO++hKBffLSUjyQzhkne+AU
efTSxBVb4RfhZzL9e/0nyk+MSQd1chcqNa4BVrbabUdYmatx1qYfC/Jg75lFFU3d
IsonMkvYVbn0m8XnCK5TTF+UbcZw8vrCx6yWkI5QvhWPJ70MbCq9WkEsobzU/c6q
SPIjR8sQHllZS/Jt0nIXA+ans0wAnV8bUpoTyzPReFa+DPm1CsVDopxx1cLr+mYX
ec32ObJgvdFrwfbUraKNJ+Oyt0IqwmYo8pUSyvQvUbuky+di840lPVTccqH7a4gP
mzoudYfXx4uhT04EyNFanfPptd+zenOEqlDHLytiSLbQ9nW7K4UAeoXysmJu/8tJ
q1yiS9lQR3InRd5u8AslrlR5WKge4DfPwa1wQiHTVhTcTTBE8RbifeK/ouff6NCE
euqIje8nYT7VzkWulcpiPgU/FrIADjmRfLf/GYIRMAQOG3bmVbnyujNvrF/FrXRn
djtVTr/fJYVKPbT8Qy7SEpiTwrSLQKAFCiUOn6csTiW/3+bvMTyoH9ZunxprZYr5
/D/nh74nwtZG73bYnnECiVgogHobcvdmZlb0YszHcFE3WP24I82NbdZNvXn73mIs
e1XqIC9bmZFv/s01BiFbubtzAoICmghKoB80Nswi0xIX+Zsgce+i5xi0VslI2jw6
jFknU5+ty7NGFtm1AQ/7YluD5Cx/j1z2THn4f9UtWXpmsJg9USer2xduU2VuK/BT
uPqXP7pI0z6keeMgUkTSuLpYalLNJPGvF6nwEfGbmbhWC0Tzfo6EWMlupKOSHMRb
MpMsdf06KLhn7B6E+BxtTRBkvaorBU0kqspjXnWvbirpIuTi0eC8fldXlVogt/6h
hWjxyjNMuaniG4xc0HPqPOGQWtNnDsIuDcgDfqFV1zgJW5ifyF9CQdHq+SRUPde5
duRbutk88JSI/yPkT9/jHxSHyiYcSSna3t8mBQZ4oZ13EXtCzCUctbu4G+dlYWac
yX3/nnvUGZ1psOrqJNA6Lkl8oR0gkzw6WaaJPia5PpxvBautfiEHGRD2bE67+NA5
8Snw9dO/IIemFQ4CMfK3eXFQTDdN8PLvsTBnHzsLztZcEIJGbpuaOMaR/unJ1aNj
0S5QseQNWETd9u+Oxl1AuJ8kQ2cDbSCMyTigHwFQbfY31ZzdZRwPELEvMkBeY7X/
ZZ2zdLL9KcnfgpvUl5wkyVEUA/Gfkvv988AKPs6sGcAPT0zDii9CbCjaHfwvml1K
CdqdnfgTcPnqXSHsaKGinuHwwzQdkiARvfWQE1DzXzIFVp4fC/FdIYstxxBIuQj+
UO9iUdB8nHLUURoMivQ9yOjPZQr+emdfAKcXUp0cpZaBrHiw7SqLA1/86PcdyMUL
s93uTyk07cLEjEGtZjmveGSqE4MEmSzv4vbWKeuJIxPHE4iHI5VBQ0NXOe6sK1VG
nj36DXPEppZJg4OIX18jxgsep+yp9h5ggxfnITy177Nw9sAGV0uqULuaR7vMSlfl
l7aLByiNACxWCEuLyldMX68RdlZob65OjsGafl72964lRrDNLxQkLMfsphna/vos
JCFFqaAc/4ZnrVFgvWEKNOOYWBkGdTgoXyhkXnDnZI6XFxKg61BZu2C1ocQItn7Y
RNynpqnzgc/1WPHoy0C5hsIyMeey/kJ403r2QMx02DhjCAKrUnNcr2GK26pCsGSZ
QyKstbPhaCjwfZIGiinh0+BKrEwxCt1XRpwqCUg4W0Oyu7maVJ2bUASqVy/VzwG6
HAK6Om3fm0p8dGTnL8+wFxAmjCMZN8cpPBlWmpwJveCSdc3KfKzSNwxcp2Xc6jV4
+U8t729uyRxWDBMGUvGCUdRWfWth2eEKQM7EhRGqQM9uTzEBIairVi/9rOsT9rpz
FRz24q1UmMdS+zOpHUUoYGrtA5Quv5+5jUQ0ibsZcsKNwVCHsZuf4dz9jiZb7nuw
Ysnh9LqTkTKRFMcKpHTx7xVEdKi2lYrSIykFCe9v8/Wwzl/Je4BuTCFIw3+cxSMN
FfkHwdWpU6by8Efvp6qGFYBJLFgkAVb6riYqsuDnm8P8RCVHW68NTxz9rE/V34pQ
Bv3lAktVB64gi7wDe9igJQR2i4oaANgcw+0TMOt4HB2cViJEe6N/wXk1bWu7M2AZ
bsEmZYnrWUoYTEHno31bgX0jING+aau97JmsPmbfJwsT51fS4WCxKWaAzSuLzAjR
W5QlY1xf65/PNypwiKHMv4oCsN1tJr037esJeoZGaZuDcAKe9ukrsBuOLXh4PdkZ
6rljE4d4EFHSd2nRBuaMbyH5vBwyhvnj2xvNhd1B3Qn+HS5ws606E26I/APDkW+r
SSFI+b0q685I///7t5eyzT5IEAgRe9bD6SBmipOnjBTuwqwp/kXP2zotcxehl8G9
YeYxerVz9UUMNHdYFumzawqUWuy7vwfXTf1mDWi67VdwxPgCCfV4eJ0HWhJBMKBe
ao2S0pts3TC73mTMwUJLQA/AnmKJZQERbH+3EYmf0yx/oc0O01ti4BX8txnsQApU
ra7Lm4f8nfigwXXcnROEF7qEnYzrhEYA06It/iWgSnhyKytcWFowk/GJoAg4k5SJ
gmd7/bGT4yeZ2QS4CPBXyL6AT7yeCMP72AAIeRRNnnyKqb4DQWhnbIO0R7gFD4yx
KjqAp1o4UAd3RpC8u6tSjK7XjOzXNpKE2jYrhNYuBe+5oB2zmmNRRp1WdEc9hD0W
WWqgUcusLpsSyCAvmeOEm+uiiijSTkAbnvQwkS5GItIp4VJy4oM3rZ5V8hScKehO
1NxB2qRwhRy3GPbNsO/chNMpMRq8DLlnBDfrKHLnC2l+dbg9opvy+1B7ytvsZyjL
sED/bhMkFYYFhCV9ZN/Ng3Ixt3epWTrkiIZ4MEgf8zLRW/2WCDkKRjOsbCaXilKG
jbIEL9rA8THlLhQq05xIffHVST7sP8aUnAr24pMvRckH70QrOEpfnXVSOFLo4uUS
LBIwX0Q9Q1waRfr/KP/+QXJ9oKXGREqBFEPR9RuYUQeJhJve45gfy3LOn2CUsCU7
YBUZGwZb2TBRyY6Ked1yamEH/24aRMBAvR4zMn8fSQ9dlqal45avtIKA1BOPAV4c
NCeV5hraKXmcYNv4WidaMD9+uDClAxphspkdA6fgihP3tOIwtm902P9Dih1yHArM
45d0ALBLyRkp4eBTYupctJHGEvvl4NWZN/pvJSOwFz8tKW6lq3/Sy/eACrUMXrMu
Egbi+jy+qASMLhmVoiTYDTRik3IG2t73198txmYvCD7JKpi/rDVsWFmpcY9XZJY4
SUCsm9tMCRFKXTNA46QU+r9K6KKseyGVEGG9pZcWDo/1NG//dpf8AD9HBFTuEhvZ
pXw+P67CK0CDs1l1HCy7b8s8+7TwrXvtu19flXtL5613Jl5OFjHMC9S02OFEC7At
FhJsYFzTE6QmC4UaNLDxfRS44jDZf4qyVlvJ+J7T/+18TscEhfsiyMcEhOHYHsaA
ZuhQoJUhtFFCD8EvNquChvlRsd2rc97JNgYNZrpNaUM7EV+t0J2sJEZ+TmWgVr/J
nQsi04TnOqbvhr36N107jOnr4X8QiePbsOYt6bx0x52wpQ07C82ZGjOeZxfSHPVl
wke7CPO55jQsdY4bclA8BBWhhI5na+ktQxh9b+9yP8+Ar4Z2oG3rnLw1BXmkj29N
rrr7XWTaTaqbsb42uJUHxsSeehqFbfhBsUQxpZMGdQSmb8dTudnBwM8+Bbp59Csq
e5l6dNTVF9RgDv8ljAwS9XmFFXyG7YG3GgfCjBJ8aKl0PPrPLe3SqnLF8DDcUBJq
auDr6y5qenWWrAEwE9bwRseVdZfqxMPdNFC5r1RusoHQbyYgYm7SxCG726LmRIT3
MFctMWFqQ/9btm8O7EYZSl3cDNdp8gyT1ECJZ9yg/msDZoqF3JQ3l3pM6Dd+KyCr
BFnn3/ecDVbDHmIQ1s7s89aOw/1PJh+x9/qYnUm0LN08xBWitXGtG8gTnuXnKIzu
vdk31mQAE/yXyzjVaX79lxJUWC6lOPiyCRZz7ArLhNHRfFf+IClSDBtUfJORiROY
3Z3MzXMGgc5CPptVUC1YLYg834deW/JVavKaeR//YeP/lZZp6qTS9Th+0pz9Bkzd
9gQdDU3wi4k/DrHiYLVIDPtrmsmm7p0k7HSvirQ0O+Iwa9DKtcJ+Pn1AyAE+IXbn
XC48QGWZk/l8yWzoghjvPvsnvJ9CoUUyAV7Re3ERPx+ySso77yn2EoqjCJqarycG
ltrQoNarWKVNEv0Szi92cXLPbYyLOIWJlDsvS7N9qkwO0kYaK3o+sUYXrKJqk+m5
tsrjv+/f2etN24W/XgQaU7z46n/ZwRUJrnhRIFiFdIvwMH2TDnH38S6zswFq5tFD
7Lh9hRfgDbBlgnhxJJ40JcTViZRrdLjccVCPp7YByerNO9YxPEs584rKamf7KEZW
8YNOpCUAl78xmLgRqwxxPkDK7rEClJdYVkZB9Uymsd948mWye4nhZ7cY6zose/3C
uKlqFKFKUOPFTVkoSZVEEkw59FLYkC3cIzGWloOGb1XL0GG0RP55BaUSaT6+ikx0
FvuJz/41up7vrLIz6qKi2yr69pj+JYIDxom8KW6lUaAcp02K6CX07GhifcIjBlle
1+nAp0IAfvjuAGioxoc9PQMuj7CEQrLdc+V2/4P0arIzTQj7pTFMLM07DvHgFeUb
qomLaGzw1JSzJmxKff4JfW7rLSmA9pCdxBvuvkX0jLm+vEHiHzcA1HWldTbg1d8D
6oa+lW2dbK6Lyi/jqQHprYd3sGohQ7PdUNymLVCJ/aPzLWndTZKjAAp5EpwkYYo2
p+AOV2loAlITMRHFBv+1Qnr8FNlLoB7m8tUd4P+DKhXSEqFm16mzgxGnd2UvHlhr
QJ/KNFHxIJGhpimGBCZwanfuQ0Cbp6S1Ue8RF06aMCQKLxKLGKRAXgQauZ6SIv2b
7IX3CgM+FJiw2UCeXLnll3mJK+M9pNxE6wGjwFr2ZQgWZQqtixXTX4RBiZdoRSOF
tBKzYqNscJSA4XjYm3fBcsxpP7LRmPivbSNJMkDzP+o4V+vTQoN3+GWwCOn1Zqxa
3ebdrBCXYhmxz1VyQuzozLA7WQn+O5qh2UGhcJ6eMfFUDdpJOUXjVjzwkv2XDMh3
RZtyTnGgZyq612A9AyZT2o2ZkmXOwZ66DmBNn/QkRstu9y4F2fpm3PeYe+920lrt
GEdD/uyXcObeFWnQcdhj7MsbGfwQwqArksoqfNJnMptHTnKvNwtN47kbkHNFjNbQ
LAUqqpWlSKXRAj0A6mWT4mz2Bjnlz7Dfmo8lCUQqpnaY9EUd+u/WTGn5aV5aRkgG
lsQ9q2CbYfztYpE41W+anvQriia13Z6OGqwTKJPZwESNre3IDtx9Qxb10OfUXz1y
IMoBtTcYKa/x6Ku7d3vzGkFZtFbA1TBH17qPHC8oVMbM6yu/1AsSTJf2lF77q6v6
9mSJYPh9o/ugNeNJR44Eqzciiyy41IzVEwJi7o0hMvKPaVCIu233zNcxktSR4ERc
uLIpIL6iCtuyktDoahG1mjam7W/AbaNI3kLjLsGjtQ39Lpnw/2yoC3llGv7ZGRzB
kvSEclfbs7/uNKsq7v/mGbpDPwzZ81VO9qoDQQC1P/aw/DdPNu41Bu+z0+Ph3iUS
qLd0tivUGhCb/pnIn3D3YJTuUqRIU9OOcAVpVde+IBWL0tAJDqdYKCwZEvj669mC
dBudJQbZzW0q1BnLLxD62rVJ/F5auPdbUVEuKpfM0vRyUaqiDdvP5boGVxLVYOYM
/unAhpTjRbjPYAcbh/jwe4hbDice++Tl5gLVeHYqowHurD5vO0SA5GUODKpciboU
cdBJnUkGW55o+gguv1zajjhJGpJsZjkVEbweS34FcoMB6L+S1LmY8gx+2ukf+GpX
m04FMkFJPrKCmtSMzJ8BE9CTIZZ/Ua7ou96U4XMA69SChJu3nrHYa+5liny0K5aw
nd5oKqGHXK3DoCOdF1OwlUvXupto8IlBKYPXhWjGro8s1AdCKbKD2oXhRPlHqzU4
2PUBqlSIZUyAFfcIyC147TiyOqTZAf0sEyjGJxAf51+d7ABPrfpjFWk+5DMaGo+0
UMnhX0l6of9KIIls738iSIaJtHa6SjM3A6Qc6mXH3U7ZZf/XYB+YCkROcXCG4XO3
eUnUPHGoFqkW6+LDkse83i8WbApGp6/0Y/+BTHySNVCm+5toEJXl2FcyMSxC+CwR
iolFRnJCPJaeI4aLdJSiMNblPmW37SdLhWt8EmR4enRjHB0YZg1xt3wVzAs4WEB6
jtklShQAIiMnt5tzJycklAl5wcClvPBTvHyxgSnaK8OSliHAgtthBXaovMHaC7SH
TbWdiQQ9vJPSPnxpd73BWKWlZaRPUi6PAbpbyuk3RGV051qG2bSd8uT7j94Nsu1f
E8YRZT0PX/Pgg7g0eLmT/8d/pDbdttv6WBWF+bFaoX0XZgx0/VEyNj/vCvKhgI/X
vSceWXFVz3MqotP38w7LEuGQ7d+MsF5qvNJmGsn+lFVysxUx8VsfVNI37RTi7T7m
IKDGwp0EBLcBAA5hb3TA3JmeYmOftDTxsYMKRqj4k28lGEVgQMcpMVTMDuK+pKti
Z3WfGItY6Ys4jtvCbEIbFACzHN6Km7V3PVatN45T/mFHpYBUq4sviYZoGdCK43pr
OKFFl3wBsNHzc4RX6qTgiK6o3lVhSWQK26wMIB5LnXc82lOanIpCqTOdInoCWo/L
jPqv4mjnECcNYIjrF+Hwo13Xxn5xQQS8GmYcGXRGpBIHeO/aG/giTkEgORZGu3pd
eCewCjzQP5TyO7IzBJOy1QSOVPYkn/xZHlgvwfwNZDlEeBD5Flf9AWqlbiSRw0I0
uOauLauKdfjVomoniOi1BI1SY0ay7gKBp4npM17Zd6ohqJ89q5WwdMrmLm2ShdX1
3g94WIEiIXO1C2WEbXV21Aq91g2MKmgF31vCi23HuaLN7ECCrb8XdJDxlDGsduWt
kw9p1rrtB9sgh2Wrzjh+v3gLFXFHrpXAT6d2bQ5wKnLkHjlbWlnXQwrmK56XghYQ
+c/KDFivOwVzAm352HtK9AACw/tdrkZoqmM1Y55WV2Dxe38HinRGQ3irENxIHuu/
KBITJCqYkkqwwMNsfzluXMnQInF/PMotyRZm9mn82RtdLlvtQncGMqZS21IJGA++
YmtxVW6OYp6JCXz8PBQIkFfur6NIFlILgMls4EFrgUoNo20EVRluaf3O8isj4nPr
0uj1xb7G0WLFh86B6K6ZijEwTHKkqaa080ltxJQNdGIWJY96zVkavLl97W8NCEg/
mzTOQ6d8u4UjKr+giRWOEufy0sy+hTzse6H/8zaPuY04ozEYSdwqc9RrWfiOVS4j
Fns9jhkoTTwn6LfVNLjBq0WTF0r24TZu9m1BllSDo350wYKKDfbweAKxu60dlGPo
e0lkhEsULSPQl64mxtc8IUYhgh9qBblfd4umcw4B0ytX0M2aZzq8rc0QtOv8ADqN
hBBdXI3z1RgYFHRo+MoQalnxltBkv4Z8FjpIeIpfzAiCjBzvYTTuuYmbGHwkI3WQ
iulVqmoFRHnMV1s1Q5/WWNpouWimi/Ut4lWM0mdvnn5ajtR5xQRo47Agh0b0855O
b8qnvGj9BVN9UeUMeDW+4XtaK4QYAVEdLnUP+1ARkiPe2/fh6SeHHelWvH19uIY6
7Jiu+w6lp3p9HKvFMrRJNPA+BAIzudZd6wJgfHe5yRwkkTmoH4HkzloMAvAhW7uv
eJpUfi5kvYEYTjRHsqE00i9HZQyC6U2euXklEKBFDwZbaI43yMCzIH/QeGjQXc7B
sOe1imTfMiPZy3QoZx7fvdcyaQnfu3sxNEbKeL9Wc5cKU8mHJPlZ5VafTtCpFU/r
CGQ2SRggNZfPgbR95dDgk1mvhnZw60zHJTVi2g38pakPvNsQ2cp+V+dk2Xkp02im
muiiJQ2m99jE80PGsxKqAppnAYpqtOt4Ofmhv8fl1cQHCCP8yjNMErlcNzPWIlzD
bGUOJZiqR4EaPWgWEeZioswpuAOOy/vSkWG8IaZRQpuFPfehfchWFLAQFOMnJWY2
5ARGDF00/OGetTk9Vv7BEzlOneA059IfytadI4+UZ3nYb67MGx8iBhQPZCMRB+18
E9D+cYlRThhqxDZjM1Sj+yKxrj5QuMew7xcaXvczfipVZc2CkdeOWx2m7akL7AHa
X1A7ImY9EiVziy7jDe+uGbvC8yDuSmITWOVgzX3F6HUu1oU3L6x6FN1FGSQKYPna
Efwk5fqSVgAUN82eX9XPcJ+9yyTOToRxA85u4etqhJOM+Os+QPDEmCP7krdsmgw/
RBpD10XEtp/W55KrdLm+c5F2hONcgBMMjwcYqKtaTbsNdgTTx8NaC+WWusxnOMco
+0YNkUR3GCImk3621PXVaLid000ruIR4gqVuPkiNKHFfY3vM/ASmMSHjS8SELw3e
FHH0xJBHgo1axyK+dCSxt0mrUfz0rLBoYxcTQ042hdGHiX5f1lWb78P46fXXAoSv
WUpjDpRazw9eXw+wpN4EwV2NsKVofW1Q53Kf3EjIhieQjvgyl69cvY4jGoR0Mx+m
M6U26vVY6hbolE/dXlLxCzDOj9YFEXLelrNIHbHn8l01CIPsRuI8tmEH5KYOP73u
qMNkGZ5736wXdoCxr3AX/GnaCf/TZ8pyzB0PgNxz4wE18/SEkxUNEVAjJY/fklhO
qQAjIyo8CDM2/52pyEcSjAfLVTvR2uvkLpuIosik5xdh1Hz8FKWNGUDeJKNwqlKG
h6RtCAa21JDRMsA8Lpe97wnpvjT6/oneukiGcT1akl8+O9VxyyhWfYD68yHgl0kN
QmjeMf+/Ys02LiqtGjl2/Kv0goRiRODVOFM1l4ax9Ew2AoXs91eDEXeHEEqO9IKk
AJLeIUepSd6fsGOYwXfKrBPJffCFmvQ/gsI9b+YNxL2Pcb3l+TrR3j4AZ5P/trW5
W/qJuyXNIzEXu0LuwEZyA2dDMhvNreDuA42AVEnOf/DDbPvltiY6LPC684xtlmpF
6UerZa0wQqzMg0wlgI4TGnaN0wk7h7Uoff9SRYi5ZZWfB1PNOefMoW4MN1k3oDNA
d8+70tTmgCIdKrNJ4C1bj4GGM7lJv39s+RCITlp7WScRuXMQS27ieOcrbzUipYpT
crwRzfhWOfSff0q6dyowebLJnP0Uc5edMpB6EfDWqA3QIeIye/QYYjX2G3j0uVBt
7oIpFqQ3SPFQGR1leiDbnfKfCr6s1RbO4Nh8ArV0a5qlILoyo5wq9uyIafxd29T8
M0fvEuJ3a841GU3vLqadD/TMqGdx+PsJW8tre31RmezG8n/p1krXk14Gdtiqk4gU
WBwaEeFdXCgF5LogvWLcDxMEks1lpEvMSigsfE3+GVSdWEM9VAGuL2UPs1mGSF5R
PwTFihmz4k5leILSzesL99wpeTIlUAbvmGDVJg5P11u6EcwMpBQDWV0J6lcstkkA
NmdUxDZov/f8xkkHojoSz1PeS0dtwwteDyTOQrF//7eqrodorlZtgyqXbxDulRpw
WCeyextCXCuao/3jpF92nSYLegxeS1sa04BHXbMN6+o0zmz6JgpzN9Hz93ULL2Rp
36feBvIb7RLUfbTwHusOtmQJQB07vvwO7wXN7VfN/qe0vL6/JL7VYRcJoAs+NtPA
dhCRgVlkEKyTsAdYkTKcUG31SZvaD40qLoKVshN6ICgsc6Ye7t5yq+xdWZs5Pg6W
7jYQMzhob+lnkjAo/m0tUiG9Jdn4yNgY3gw/ib30D7G/dgwSo+aLqK3plj+ypA0g
zorsVinZdAvAP5VBHGJUakf5icE6PKOoax+PPvyyxQXKny5rq0SoOPPbrpUNBlR7
bCPcYYy/kKzNQKWTvrMsJ6WIIGZ5CRJyfcUfVdRU2TFdaJKZ4ft3CJAfxl3uRAlK
POxp9zwkQzif7dWVCyD5m8xeuZeg9Hln1y9uitzI+ToHe9N7cTb2SgTN5eMBhL/w
JLnZUvwiQDTorpmNbwtWaRCtCtj2Bi6I1c50kcCfowK6g1a51IXTmoZKfPK3eXFw
suCf6BXFBiNoh4AlfXnfKLR+Tkot9XxTWbZyiiWvFOWTkJdahJHLoCxSE+Zq2WYQ
ze/8PZANsZSmxs/y3/9HWolmhcI9FLvzosczT5oyQ9H3vhPL+5DCfWLj8edVsm+G
L0j4PcAKREVu2krgoc0JXXNhBhFct3Kl1SxC/X21j20Yi8x+NWI3bPn47V1CJ6bE
tGNxnVu9t5LeMPmBTq58h0nnbdLhqLmdzVs8jbb/TtM3KQuw8vbK2ykvkwalUkoh
PMLJ5n5JZx08i++Obt9qgr55/MRieIJ1frOnFRbMErr0lZ5d411z3oyh2kVgTak1
wpwoHZvFrK8Eou+WOZtpYZfzZ6vHpoIpd+lYTR/ez00oQM2kEgsQvF6+HBIDFOAo
NKAFvgRT44mfLBFO1ZX4u1McXrQFswv0wtibpH18tmBOED/Frmhlz+K4o5IJQoP+
Dje503jBG8aM0y0UEGOpAT0BVx8Df4aY+hZ18MPO9eAh4Dw6Aj1RVgPEk55XbNJ3
4Z70S/BIJSHfydPy9msEUVmapX3XkD2jJft+6CSpclaNkAihr18wCNg2b/rvPsSs
yJJX6dNBGCf5dskhVCQ3sAF+6iecxYa/yJ6T7umJ0kPufl1YFdFmPTmtTXevFUkx
1ecgLIX+FkUU7r8FAEQlPxQGoeO3Ov3hbMKYmBHdc4SRi3yqJWnCQzdMrIXRWdva
Fv65rP6l2iZcqx/Bnhxh8tX43p1BQ0zDBacLRryGUbgZ7fOiqbY0Q4/2lO5BuqDp
thPz5A5qSpSWPyUPRtXoMhiah1P1V0XWBykaKeqxNnX/oiiaQMgPldlzxY8SJWGo
k/ZGCUPdBI8Y/P7z4io4/Ei69wAi03xeX8YweKPb75tucD8e9QQxLGURFYbyqLnX
8tu7Y+x1QOZ+YPRmTBxntm/mEdHiY9SHWtDCISMxVWGQo8kzunwGak8HIAghZj1O
0wFneQcFMWYG3jWLZb2RLq/NejYQ92yN4F9W8nkJEsW411+BfDJKn+u0ifptPRfC
W5hFco2ymjcSZBW/mdXv7jHNErmd4ucqaoc+G6Rjrn0YjZy9OSjeNI1/1OWdMQIv
VMa/n4LoUI36gAzq48/cVYWCrLC37D2aywY61GTawjRcju4PODG8GVkJMR0gGhKL
mssYkN0PYiCy7If/OIHE8iHaZXihv0UGtzgmrs8OgKfIXKjNI81x1FTpzA8rr5PH
E1l449WZQrRS9FgPywn+HhwD8iM/6l//ItgMNPIK3GRjUANFoLTZzSwstQxViErf
KMqUCDCNpYiutyQDe5XAfttQ9zR9ep4JMTn4c+3+9Hp+DHhRvwa6AVAYutsN28g9
CwH7xbcTdxKZl1mfJoAO8zg3Z5dt0x9ivnRG8WUsDSCFC8Mik+HjJmCeru0JdvFR
+0sghowVuZ0T1aoGuCvodf+wEw2Z/vRgc8xmjl3rxZr5sUn4dtLfl2OlwEdGRnRm
bBm9LLSMB8GvBnIIBIsKjv6fsEV+xlHnDxirmL8+oKHVfaJDRFypcIUxp1EQjb8q
FpNVA4dH4+1Dj3lVm85l29fOBPkjsUn/9cEy4kdEaRpsUSKmS3mWAUNMJSRNQNet
fpxp1StFkJmVSqk3uIlZx+xsSJSTcGBvUNOufy1olLD/iVASvTeCIWeyzFoF0j0g
U0x7nSMbam6JMV4AqsFeh7jbVUm76uY/RLv6AU4RkilZWbQmc61fl4eAqHsPlFmb
srKt6qSSZvMEHxNYzMKFnl+R3yuiwdBR2WIreLnAz0tSDpXz4966NA3hu57Obk4H
09odg79o67ycJ2LMDSYheD6YnzJGyX+y/xXG54F8rSQF9BBtySTan+G8aZvfzDPB
nQBc9JwcjnkVp651HsELGeDISoVP7l4k6u4fJ++IywqfWsqguAywZ9rXAG3U0D84
IpA6bGmddUnkyp0ThDBVuuU0CwaaUfhZCnGyPjYwXw1SFn4BwOF0xf08lIei8/uZ
iLFFiY0/zG4uqm7GXIlE/xYLRvcB3A2IrQ0h6ZGR0Ae8ZQDgQs6fjV8kyB2s09sH
V6QjM42EOiNa9FPehMKFCjTrtR+MvR3PvcA2YC8Ou0fzLEwKKOqB8rBbqoB/wgv9
IeRkYY0PITCW/AvcUGFsD1Yot1WHQzrWY5L59/HeJNhaXgNtzKZseKkl+x7IIU7A
mm7j+9+kPwYOmf+IsismE+77q9tLUtTpCnxNVT898PMNMDkO+sNfnAXYZ/1szH26
qHVxGQzTEidOHjapesxygbpKvOt5EGDrK1IzmhFeji4Q/bs+gc3pd9fB39LJtI/m
WX+pUFzKM6bP5jZJRsv4Msjgz4pzNXdHoTcw94wIJy8W04AccR+oBHP3sZIlrZ+p
ZZyXyP/udTfZUTGwM/gxHew1CUlBKTVwxGAUjl9n/Swzt2hm3PoXF/Nc3HUQaZ5N
ccutPquZ3WXqvp6a7jkx+a+/xYnka7D7QuqspMDduypTtJe5Kem7SreEkRDthw1T
HjuSrFKCSSyeH13bR9K/hLDmhms9MIlaQzXy7qYjGkXrbQfjMpQMpvpELZ4cLezo
GgfgJpRLf9JFLdE19uftHX7rY1vnTD7uYahQv4XP8cxE5gCLhbIixydFhXMiLnON
fOwW3ZxeUajP0edH913ynXLyub++ug70QfvquscuE6DvsQgHk/mT7BMrPdBQVLqd
FtGUVePQ7Jey6lOnwabnOSSdyYJMwvFHUa5kOzlWuWF3FOJ8qoieoviTvsMAGZ3E
EZZuQPgmNCz4j5AVBHbSBFgv8qsYhacXlf3w2Ath/dF90GlJTQI8pXtwJAQ+lQBr
rVuywECnQvp2+iWjDCKCN7mX3PJl54S7BbR2M3mlZqtiHR4F0u2txY4yZ4LQ2oBF
8BpTdtRZaUPw6vQLuovnb0+dK9RTKU0M7Q0uRkDo7hpW+1L1/TsqdCv7XqtNBGXY
aE97DQZVUsvIIneJUeieyhZTpEiGyS4A1qdrgGmC83iOkrJiKE20bAO+8nJBOgbP
Q/BpChK2jV/n5tQNvBKpLOZbvy08wgEiYQDTd7bc3goo6k3DleseBtRQnH8NTMdM
Z4Yak7I82+/dTU2let3onwKlUxQG5GXUYKNHTVO/+4RJm+Xd9JSjEbZq6mbcdwpE
r+UfGTZwRURleN4nGicXV8WItbE3jX48BWSSEqR87qGd1IVO+0uzKTcC8cFC16Js
Pcfo7G8J2eRHPaTvOZVbI8kguedNJ6JC2rwkBe+lcTWocRvBm9C16V6TQBm3LUhJ
iZazxr6Tt0sRM7M+OAGe0tYwWAQBStDYZWpnVqOx9sfTMHndYmQFYRlVhZToHFi7
H2HBgm9CRfooWaczi/YDbqkYHzZFfd6U+tbLv9KyXJUhyk06MYtsMokoWFwK2YPT
qPvSO7OhKRGtD3/MKfwUutCJkayPdamH37H4sMnOQrwG4wZyN/v7gpVKq31j/l2U
gYMwaiVjiVA3HqJ6tLK5cEQOlFqmJHvqUv3xWNYrnbwVeaR2F89HqM5RXyVRpI5q
+Hq7cxWvEksuKe6NSGNZDnaowQ9pVAlqHWXvxnqspZ0rEJmaFO1L9JvU/G34vwU0
xqrq4VDHI5ASjhZKSk58EFzZ6wTlZ8ICmONE/qBX4P8Uai1tFlZ+bibU5NSBva+T
hvwWbtQ6SWpDS3jRHxLTxqod5t9W9jE7UetvhZLdEvBiwahbdBJwNKqq1FysmoTU
HTtKwVZAG7DIJKn3STswltdWbCsKdKsaWHNLBZbqOL5A2YAX0PEgFZyQIAIK0bY3
OSlaOw08ShZt9/XZBWV3sbAeDqhhTJjBfJxCW0DZuwD04UTAQspM1WfI2LXQ+FMc
g65dNEvA0asHYNlQIU6Gtc7gCMOT0OL0xczucz8/ZewlA32TU+3hN8US2H9SlNeH
dzqssyllxxBuNJkVX15sKeKsWnyuqkGsB663FnPdAmtDBBIg0C23viRHxLjFvJSx
IfftOT0vxe/y/GHFYY8ASZkiFsmxd0kDc+BLaAdg1vMg8g0gKJVpb4CiBw6r8KFa
lanC2z+jE6NxXVj57SP4OqYraCEORnAu/FNyhQeUFxxWOiAWIPoJQG/7wtvjVGzS
Rp8bcB3rH+fFNm7UqN6ELgIQW6m7Z8LFEeDuKP/ND+O1o538IaiZZmDlRuIz2g0Z
x8dz7T35bNflTVGfVWH22ACMjfc0upX3mA03GlixdnhP6QbX7D7MT9OJyhMm6Cur
VKHBT0yTDnLjP0FMZ8ChWwFtfPwob2BDTG8v19zORcmSJbiNtdDH42N06UgI54Vq
C2eySoAQv0ObYbzPD6PgfOPKojY+EyFGiM/oU06hawduBfN7XHbf5zEwPnC3YYLv
Q4E2NUgqmrZanJF0Y38WsvuG9HpazSl5LluvYIbfeRg0XDykBC4mHHuZjznDV53i
nciR3tPhHsmpGbSHj1pQZcnbZ7QBTTSpaPUba6GC5XFRzPhnQAts61wB7g2X3eKO
xTx1onWGKxQdB+fxqv6+Tj3Lqljn2rfyBclG66ageAxsDohA22KyjAHb4faXu0k9
PXKKFODvFH/4GFZXJ5GUSPYOGuldtVmmJ99U92zLmesw6J+RGiqCxdk4iXFoWJci
J3vA/xGrL05Atz5AjofGk+EkfgcJm2EU7nsIdo3XRcY+9hqF1APf6i5nwq63Wn38
ihZ9tFDsDlSa1kaqhDilxzGUbKzhzAA6Wm0fU+wmj0Qj+gELs0Eb13wo24fnUDbH
kqT0qOZQdEF6LJQtLAO0KhIV+GHVARdDo/kFO3edPir3weAL5oPi4BHxnWdRPJKB
3eC4aDyo3Jq8NK2BOYMLnPAQRY7i5omwa/9nQuVTuk1ooIXX4Fb+PemT+zaWNi4E
S1S6mJXNBtLPahnrx1DDnVzsN60z1xU9ZNszaeBVZ9Wlu8nLxVoAGTqWdlJuHIgL
NiKyExdmwg6DJloFHZarZ43wLU1s81Q5e4A02M2DSMasvXfEA+8i063uKrvhb9IX
dq/MwYnpUHavCMS3fxGqCtdhL8mjf4UaS7rYXytrC7jH7PnD1YhordWqQGVTsvYF
0W04fc+U5WGXGGirOBPzfy6mukFyz4YOh11CvpyQDyFoNXAIk1RtcUBiy4ZHfTt2
gSIdoeEA5gtmfxKFSEk+uPlwe2o8nYyAXJ8/uy4g7bZtQue5jY5o6yNPPUh9OMCo
0nKXFzNyiMQ3XnvdIBFqZr+QHKxlm7sP5lyLh8Le8BH/9Gv7PAokJO9gc9F0YSMJ
MLNP/InHVNCJriopTKtB54kUaV8fp/KaIIXYRMks2JPB1nPJBLGqlBVq7nwBl5RE
K8u/NVz2N56QRccYVL7illaM/6KBHAGABAd3pE5dkRYqClWkdlkyWljj3AaQ1xyZ
/6ly1yfvToMrR+3iJrhURh/Ju28ZnkDkwjdxjWweuXb0g32vVBI8VVbEmr97Hsqi
XVsvcnPd4ARYArJB2S8wITunGdMCNRNGHj7aqOv8m2Q6ExHedlXZlp6qryP8lESk
KBdzFqiVhkVeIeGMMxZk2Nm6u6c/7uKH+Ro0qyU8G8T+QFuhWF51/VOhk1iS6DRP
gT9JNmxvMatkvkD3b4nOxHWCg3RPRVb8LjvDyT+o9EXBNM3uxsdsP1oDsbRY946R
/Am42t4l8VDOm2yQdKMiu0t50dq71KWIbrNZwHCGNhRFr1ZZGDFw2BYQGUT1tkpk
3foYOrk8ybokg8XjgH5Om6OBcu5H2rot3QhlTaB4mRptpVQ83EXbmnjYxGhJhk01
RaJIIt9WUp7Jss98QDoMQBhtrTGGg801/gvsJuEiEwBiB2R2US8bEH8ySnIGXghN
o5X34WR/MV+viwNG0x5JID2Rz6HiGItMCX3apysEYzZ6O0ZKlABwRIVt15hrOTxX
hq4yVDshDqbEBLyZ6Q6sRmMoejLlS7cXaMSVFyxxdZ9iG6Ulh5zqeZ0U7V5OcEgl
5TxAmO9fGL2C/BJkq8Fn7V4plXadUeFqLP2m+82F4BjU9Ivhq89w7U2a95doD9eS
QxsXepBF2fPojDL57PekXoOweVy/sYz4Hs0n4Wqf5Cs1y/impozF/E/tsACoov4z
jwsHSfPRbswz/0tOBcmOY9VBuPwKbytEE5Bvc31e8v6rBPaEolgQUPoeflkWVmci
x7MiSz+hp7AN/Qk7B2Ds9doE4nlzIqga5iUi5hD9lwgGwAivkyedA4FlYw9jZ6Ua
uwfVkhptBG9lPVXMJyd+06RwIZ+cGg3Dga5q8CIGAkKpZqd5VkNB8Qei4w6SBHK3
A3MhhvDl3GWm6dyC+owBHKDY4SvuZd4AeD9V+jmarvD7ycG0QSL3/nkx6VNefWnM
BvCrVsC2WX9eMkBAl7nyduiVKLZP1hoz0exagayqkVTQFnyxHf1nMrkPLbIsee37
+An0W7Dh27mNjaVbuzoUaSV8OcxtTjBDxoh+fUgqLz7MQ94xz2zjYVFqWh36OLXc
MJ5Rog3pIZ4MAbGQVvU5Yj3RaFVfSVp/sRNqMuUa7++0yATmo8dV1TcruI9pkEDq
IVV2PuJj07ls9ho1QcGHYsbwH4L8Y1nAvJqOjQMn+lnYhbXspsSUFEJK0JFnVdq3
9hclY778O5/81Ns4qhGJNfsTnBkiTvBOm3mVvwFV5vJezoNtY6S3R9vcgXZi2/4i
Ip5x4YW9sONZSdAJfye0PFHH42M8D1Pn8Dlx0xVsc/AA8owBNyy8hd5prys7ODSS
L8m6yrLK/f5SqefReKz8ik2bDAILWy9GK7O9QnEjhGgqURs+J7TK/bVzuOkGEhut
/Cf8XEuXZVO0JdzD1Nl7+XqzahNRXMbFcFO4+F3EPWUgD5kmDYoIOgk7TacpTAn7
n44zzEdPow4DFCK8qCTomL1OOrGHL4U7w0TlTyHKjug6RztZxj/KTsfEflEoy9Ni
dS6fX9Ws+dWLvKXuBdxvwE8alXNo2GGKnEOf/4LRhacNiC4GoeYw3TAsCOJCiz65
JK21A8QMyjsfIe8mSvLsXdSwYlWKftOkBfKS9poJ0up2KrzQ1llDR+GcRzlx++Ew
hLEGC/f6QEP4fz2HygK35VgjRkVbboVRpILGX1es9oAzsCGXMPpsfeF5TRys4HYg
5sej5sDCP1/nvQPoyeGv75MRtZvEHUuEWu++DbxXkQ19m+yl0dezCA2szcWlGJmB
6mHmAZ9EubX7Vwn3NtDhXrSXRIJq2/rB1eUHsvYpyt5T950z55bmTUb9iSkJrPXB
Bd6Ni2u8vTNIfjaot5h52MJR++NVmIDaHuFEW1OUws5x8GgIC+C7EmJPLoHsM9fP
s+BW/lImR+6Epg6B6WvjCSNA2U2XyADQQYbOBmqq7rtom0vqM0JOSD3Rd/g5rCPH
jk8s3uZt3JCfsHBt2moi9clZyOSBiA0ecwRVp3fFJEmhM977jbU5oTG0BmUk058H
wgVgyqguwBmU/b9u9v9L/7iidxNnfvCg59SEQg3kMCbBKwpsVU+StF62NxfDMPdJ
1zr0jfxNv++ekXohMVueUy9ryagv0odI8jBpDRK1gffRj9Ex8nBbms6N0OOJshrN
a3J+7pWTsSOrGih4n1kJI32YWJx3tlZMVk/DVlC/RH9HvTmovDHmJuUJutFsqjEz
HzWDTjuFdqS7siNmqNnU0FC1FEN+0sxOUNpyvy5UCxTT2ODhV9sGzHi8p7j4Ds6l
x0zV0+r80ypKT37pNjLlAA+46u8FyRyZjUFy1Y+pgrZon5Us358iSeOIJR+x4bO7
c1SnENVj+KAJN8Jp7aEqB667JIExylRJHz38rcELcvqDYOYt7BhaZ+Et7ec8EvLE
EwqYemlNF+tIo2CdgTQFYWbJ3GFmPSFz5m3lFu1BEq+xUQA10AZ8FEAPy/Ag4XGH
yhcOqFRn3jTZ5IpVz7OFzIV74yjS9rrDnIZG/Kj7N3XC/I7sZR/FeTlmGi9JsQzt
x20Hq+ecQHpoLe/y1XbX3bvkgqX31oZ0qn9k3CFWxznbl/3gcfxEtxilPhn28s+l
Mu+d+9vHQ+H/LGpSBtUEy7sTn2HaAUlOebtlL9273S/dUbkSEXYkhYr61Ov4qfcU
xBNJWRJu3ci+NuZJ1p24lulI/dogdczZhaA/zlc/uljmlHAv3C+Gj12E9NBZBbcu
KMH+kJ58a4WtCcutNeV0SJD8WCNrxIrQ6BBlma0po24287992F3doG80kpssva6C
1wNKppBybL5IdFz4TxHi3ZSQCmLxDuDmEZziFqN31e/bm932qeQWlz8AKOb+23Lo
oVg10TIElqKhhONycAolDV9/onCRpXeII9hdYBcfr/dwj6MkBJcLHT4y3PPeBDhG
FKxmR85SX8sEpYDnVDMe3mPBvMjhcbRrhd/kYSiThnzIJBp/gpj0FL9bALS9jUd/
918ozt59dDFuB7W8fjVVzoHbQJAm0f81XuvUeGKjQX3Dco2l5AYvtFpytjY0gY6G
wshYI0zfRplVB3FqCj8VyKZEUC4tqg+bPUAL2bxSvH8+x7TxmLzZUB8e99uYF9Xe
9VrnQywSj6jUomlSQ0xJZKlPcClDiQVWJNx0Xw0HUmC+sa75xU6ZrtGujz6Xctpw
fZUyiI87RyXo6iiS6WY50rOfR4ijh+8s1x2RqTszgdEOZJ/pw6VEq7oanejpvBHp
vzUOZjXwKyXUJBCcsKGXDf2QUVsMlAxP84otkbkH74jwVK6tTlMUTo744aD7WHCa
3UcsH6+MrtiMjRG1kf4EFwrhCSf+8L3JIbINo9hBrZXHU10Mw355PRrpEOD4xlm8
PRwQ9fUF1q1jW+tAk8nBmF840KcVEGBofQHo4/PefhU7HHyWFo/5zv3JDoPCrNa1
4LpL9DMjf9Tu0fzceBvYxxm/rI0mVvc4YnRCaiPVcZ8BUGGugQ8NQtPKSrT40rhk
gfYc/5oq1Ek407nXJgQ1BicN17JWrgXORooeza8lJ5Agw3j5wozlZFT2QgP714h0
1M9xzSChK2CJle79IUHBtZU51MT6nMpNgq9J7pEUky0gOVjQQL63xiBsG3bQ+syj
IEGcTmfnQv/Z6ipwOwID9VoLRfigZTrbsaie9dH0Ci1YK+03LwUvuXqIVX2Kx5M2
ml2419ZbSssIFQIEg59+IWFpgK8qzs1YAoNK3Ajg36VsTZkPv0R0xUw7zoUBo3UL
UCPZks+m/aJvNqg38hL73NiqykmyDehqqhch234OQOluUC4vFeP6oEfRGPDD/jEb
QevtrBZUlLlYbHGktnzN/Qz/VSybfwVkUhUsNvPc55qqiUEem7iLpT/vBDk9ny8o
P9H/pBre7vNPhGHJt/dMuJIwGuexucOqg2nR18sCPiYNlkB78B3l2uqHVUmMhKRD
rrcug3tJphGfXSL4TvesRN9ZbKBpyOiOHlKMetQ0Y1H1TD5aIACd77ZUgzMuhY4V
4VOOx4r5owt61Ku4LLO5/5Q6X8vdXozp+LdVteFE2NOcVDT+tzLYFIZSNcIBa3H/
avFWrgDn5mWjO+X6OeAw1PSmycNfaLz1O/lopjTjLVhJMqGLDRvIhqzKPz04fG/L
0vaxV8L9g9nQEMdttPfu6GhX4zUGuv7leyO+5YNjiOf+IeHRuyOC+7CbZaqsUmjN
Cwtbm9DGO+4oF9oB83C+wjdB4JygJz84bCe1DrLAhFoblslIS7xmbPJHAvsLIJmt
7QeVjlt3PM+NONV9hC16R1eQ0KAXu7btpI8xdtgb9M+qTrruH5MKBxNsBctYU68Q
yDdCoLSzqYi27iZ9fExIi1obRQn2w6lrAhgBob+lWF8A5uAzO+muU045cquIp29p
19F1WUQ3+T/fJdvUMLWFzmGZx0fu8azSIVvhhnnKTx0MM2A4Afav7zUobJYXr7Ne
Vo0u7b3fwhYnvG2BneiMo9yxFpnW8wEmj7JhaVgUsAS6qK0ltOucNFgmIwaKttdu
MABpluMY9v3XI6KLlETPpXF16Mc25otDSwWKZS61dUVT9HThhrupY4TpeoxugePA
c0rUyWaS3iYdjoKxyWZTBOFhKgDq+v8sioDu/mVxXgwKwAt2VCtNxy0if3BT9bZC
YXrzUqvWH2bJWbAHOqyg7tuqP+3cxzP5u/WvXbwLsqJUkxBuihyQDVMPueEf5AFd
04G+oUm8zE4Tg9wq27IjRs+gJYuDiQAybauU3vmhqxI5vd9iGbdpic7J1d/RqCIS
NVYYLrN2LDLU+DmScHyyhBREoMOZVYWB9seiJRf1e0jl5xpD4qAO7KiwMTOfm89J
LyxXBoDqU5TTTo2TcmfT/lJEh+Fqe8X5fri1TLpaAnl/EhHRcUy7yOb2IE64omwP
bpfKZyqTbBrn5FoQvI043IoZniEqP9O6a/tJ/Q02bBUx5RkisfBaXf8zstCidEFv
+I4CIJ9Njl1VaAh6Xe4910QGwHobtdtWB++BvkK/IM4KFLGuPEy4pEj9eXJ1LHN2
oQ1yqxjNVDl0BjfOkFhM1kVMw3bTba4Krk5zf8eJnGftlNrdq89juEGu3iPt2QCT
lMb959kFMZ7hLeQZZFd0NLqZ+KA44ajrF/cqVjYpvc4+wTqNZ+E7tjPDidKg8SDC
OEj5WKCqSy9tfl8oG6tBbM8qDJxQuNHR//G5a9iowoVrrEUGCSNZoyzd5YjfNHgL
X/EurYWRoS0hCrpXyyAg4txSeDzLlQBy7delcuvxoZJg98Vt4Z7VEwVUy4+Mpgrx
W7z4GAls4E1bCr4ZmrgNazi2ZpP5Wj0onybjvmunt1iTW7vPa5g+FoUx0N6l1+uA
NH14exhdJM5K8m4UBHxViTBMOSSdfmZvlpQeqtVvU/f1IeQbVukDCGLpk7uRJGTz
BPWTlYBCsW7KDmOe5+ZuPJBWGfkN2LQLyQmsBAsHuQiaEMNlt+JBb/Hvdmv5WgKw
HP2O+gKxdospwTguJE/EvywELgRjpMFZHcAzmhGZu+vFDVjF1jgQ4qvLqDbFVrVF
ivvP3VdglxC9dvygaj+JJeGAePRy8XmpXaWtPML5/VAHmroCPl0RRI5o8JeZ86ap
tvbGE18TnZp1r4cuHyH6QY1ZmWehXLrWQnRt/9nL2e7pisoXEYYcCwIiQGghMCrk
fazy3UFA4zFPwST5twHKSH37G8l9pXI5oYujzR1Hi2/fbQCywqfCchZwqxtlUO3V
I5k+wtC0jvH30h/CIdutwdvBxq6IQ+vTWBWgQKLPcht32vPomnz1cRPD/EFG3Msx
bTNtPW3Zel2rxz00YhrsYJhG7IAWUtCPOebqDevlIA8dzusfmLcxMf9/loAeakZ2
XYIxCBptXi7/1p8s/UNgqxjQASzP/keZR6hUiGWRMG5DW/gaicdVOAshUsR5Qz+H
8n7VuMoi+/lII+iNnZG0tMDLZDOSfbIOqV8uVQdsJ7fNxY3qLyeQCPZlUS/LMhpE
4ceQbkh6b3zKjAh8H0ovawSlZz6v1JYPap4QaSgzhbdh00DmYk+3phRzDqVt5/Vp
R4V1UM+fCOmH//03BSz7A8ZmWIzqsBrKzEPvXSqe/FfB2xc4lof0WABqbiHvIblw
MEXH6qP9dXLk2eZ1M73f/sZ4w5S6oIPM0vvojBC5bwMrVe2pCHcMmYKr2P+xUpoj
4WEDMfnErP0m3EmrPKEzTgUa6gjgq75/9NYc9VF9ONSTUbAeWOdZKJikXz+d+HpE
BSnytLgUfnqJbtoul5rF/QfOslJPhar/qiIIhNc+EJoCgZ3kX4ImYfc6F1Lm9168
WrNnEF3ZGCg4ccanUbchDSGPl4821oPsW2pcOuUvaMC5jdc2/6m98yaOczFPoyeC
5vn3ayh87BYe/FAicDu+YUFhjVdSZwFaGGi5zSrSbPX4WmoCECAQcFQyaSElM1BP
9zf03dWUTw9Wxf86Z17pUnLipG4UwsuoWwXGGcFOyTQRqDOr0VzlglBWfpBu/gpa
zLgjYTEyKHupgqyUp7VQNKLFnzhEZ1g0oEKEVJkPhZQJZ4/Uw4QYgSuJOcs0UToK
o73CgnJr4SXtuANNvg1yXLKoizs+OyQl1vD4/jNLz+zrrdaxTf0KooZyk8uPTJEU
P3G/3IghEzSBSoqKHsZFcJn4euwgHaPiCE7mtANOAjxoVrct7njdLBQ7UNGHRM73
RksZa2SUJe5ZQwU6FSalNnSNTMLCKQVn+Lx2Py54X/IXK7BYYX+vAnN1cvkVmDwO
Ag2Y+P4Waa+pHApc8t2nxb1YoCIj+cvkwWvOLiApi6ja5DaRmqEqj4yYP+o7SRB7
+p+cqcsCSyf7RslWC+IP4paYsWHtzNuStmmmn/fpTUgw/ZdpQs/B3b5yOJVxkb4Y
KWELyU3Qio5VUUbj1j7kwJdLE5Cc+PUABsq9Yo6g710ve8MeSkGVquQVgm5g+AAa
WV0X/EB+G5dGPkCHjB6F99GkQCTLHikSHXQnAXN3+cwpJTZ+7GUgRzeazNTUIfTM
0WcmaouhEsqdyTDxmrCObCBHG3wxkW3IV8XeuhhiVavAo9ZHmw4X9ine+dqJ/qaI
JyOaAYO03dfpEYVwF37zHObz3uAqNctxvGn6AONqtl8PhxVsR07pAWviKCdd0SAH
YbqS7HhA73AVCKcnmVa3j8bMOqgKpp+o9GFb52jDc8LSSt7os4PR9mWWUnvKtyXe
3csfpdVsuB657SQXNJeYHB3fEqiIP/1e+DWnpdchyYmn2iERWqj8+X4e/uqla0Js
pgb++ZY8ZBg1YJCsSavw9sa0kBaUc3YpuMFfCf+hYDXSguhsVCgDwNoLtWRoKKpP
Tr042O/00OmJL91vVL0yq+wXuNnTw/ofylrYw21WsI7O3tLspfGZ/lKzODZxoP0s
yR5DQLJrQCktYeNZKJ9y5z9OloNEzmttiULA76Z1dRkJl1dA9isM+EiXm5hvcwnP
YI+v6p68bu8V50IFkI9qU2nn9xV+qnBHzCwVhXpFNloBJwmeOdte8TFGmdBf1w90
tw78FZxM2ooYCvQNGbae03+tre1GxeakHXWZ7eoIoDNLsocyJztYFKCJoq5nZ5Q+
sa5QvKEk17c+LOQVeBFF0EyNlx83Tk/XaV8kKET81CwJEibedsZ7bg3K5wMu+Ubv
nP/U0mWPXuXONGZj05A4WYGWqWAs9P8jPklQuKFv9cIgeDjTRcJFPRGqwqAsnA3K
UBnJwCf71RQudBK6UYbg3Qn3+6rwmhcECFJMPbhgMh36LD1GtbPLtCmlqvo2UqLo
6diX50rsgABnd3wNwrJJl2OTHfoalLGr5luWHRkq4ph/ec6zoeCzXjsWoGFma0Jw
RDon+/6Oq+0bLGCMr8YCf2qxA9P5OopIuZYMWUU8AsOxeHzUUEhsxjckTg4Rx4p2
tJCLhT2YVkoVP91cldtM8QHr5eu7IRYFJk0RBXMgayEx3cfFGuIs5VYdLle9KVhS
66A8LGiXz4cs0lzq1ABG5F5k8pVuZePOsokr87o3J8xEwcs7/IgysZKXrwNjiICK
cXTpZnF9rv/HSjd1WwGvT29UbfjFpW/gexUESOyGhFRYCsblGpdY5mddxrzvot6v
JSyhSjdib2xDyM1fshhhcpFpoa3KDWJlt8rrI8DDVAKEaavVU6yvK3jHlu4AHIcg
QvIqMqtO5I1TtwtMOqGqpc4ftned4qPveFVfvKNYUBrWUjWUF9GnCG5ZivoheTMQ
MVCXSmCMi79eeRZG2VzaFjVkV392h/U+o9aIRPMFJy4WgKd0Jo5eMAV+UiqXTX8x
hhGDy1+A1PpFL1Br1tmdFJYPrprj3oztf1ittdVF6aPOgY1AUE9tCkHrOsaIsRAM
Da294GS3E6c60n9YAhX6ugeUhcCSR0eyV6lJyCi7ELVtrmNF1YsaTEKuteVJtvGs
bAY+zAIAe8N21e3nU/XLJq5ee5arY5Oc2mmLuPttqNRg0n5gOaAVhOMHfuYU7Q5n
ACc7vi5SCY9SjGzglOexiq3KoNCtbYwCqHTnF7Bcn5T86Groln6zAPa6YAgdHYvn
VaCbvg9n1l5cbG8+e92R9he6QQ11MMJU0B41/X0rZOsoHE+sojR7Sf8JlApE230n
Mfw0c/E7m0bUjBBak6TAk4367uIrbgaw5xK30umEo/sbJsagWTsC8dmzRq+MaS82
tiU1J+O22w/AfCCVHEdSWmqLexzsTMU75IWWB2ueuo6MLiEpY55/roQOpqLx2nHa
95OZCT6Zw/apAh4Zy8UOSN35lzYGKtbChLgZw6tO+UGEVPgc19invUfTsfELsTwZ
KR/gghnqKeORdbOfAOm52aGXmKUNvTkgMIE3Fzmgx9u87SjJA445djDcB5fafiVy
35TZW2bH6AN+SIhBJj7eDLA/RarjMP0soXqR1mQN8cyX527NH5Y4wl742ljM9dB3
1n6T7PYgx1CUbHUInaN8oLPnfZquKh+kK+4Hl51p8iNYusPq0WW65GePMsJVp30M
cnwP1iyoDhq7/Qh8fUFc8EVYry/SlJemLyT75fSq/OZObJznWUwsAsUr3cFBNakZ
oF8tUW7VRiWLURmrTJjEyWx4VQbqNkCXbJljsXr/GvlNk0LFwD1ERNA+9lxE0r2t
qmD4xmiHETIfxM5vYfzaHeskJk3wCdNhXEriO9+pGg3yttmIQ6UDTJtINkubeffX
e94iYxZuvbs8CNRJrZyb0Uw+qoWWG442yL6/1KTGU7jxh8Y7yxRupL9LGK7zXvRd
5oWA/4geS9RbQlxOoMw8vYQizxTTnTCZe86cPVHR4xs2IZrcd3kzkxMNsyMfvli1
/1x9kRFjnZsPh8X9eaeNccXVId0na6HHkqHUI2LJ2SPeEyZUhSg/PMa1sThE6Rn2
6YBZtRPG2HJDE97Bqg8A3kjkl/kVoCfYPxTeoKLooAlmY1tFU6senrqj0vTk0kqj
sU3Kvy1xAEI6Tnc56/i0Eoe5gz3rDeD2nQnATiWXlvCrsQxY3nC/B8HzlVV9XRQn
oK9sWET/FSCYHmNj8Ogsw8FHbWtFxBaKTI6GppKljHyEqWVRNm3g1cR9JNQqESOL
jTCuw9BGav4a83ZLEdq9dYeCBio/d9vGrZxSMgkOi5lb8yVcukPA92HWwlvH5+hf
rfuK4RMk0StiM/OKvJcIleX0Qk0s9cb5KwmK3sSLS0hC/XyS1oXODVfzE4rQHIEa
qR7kIiYaFXXsOjucUL8r0Ar0sdsLJbQ8InA2HI7k1LAQfe5yIEN6E615pqQFJTgG
iCP/yUQZBAsjgKAduf5sL/h48O76W6CanLeZNv4VnTm9gbYw2sm414QSgHT6KdRk
QxY28Pin6akVVIaGwC1F1bBNgNQh02OCzuOHdmAk0sHjPW87gt8B+jSkfbSbBqOl
9cGta9gccUBnfMNEMe2a2FxpCjQjGJaWEoZ0WPPOpshy1aP/RsqGnZV5ovhaC89P
Nn2eW36BKimIRjabAjlqIRUEzEj/c+xf8Cv/yuEuD3tWac8Jsy/vhOCJVvkU8106
bY+8+XcsknzhbPo/YViNWhCyq+YuW/hzrE7uyL2SVnbj9b+F2U03o9d8UVjD743t
gRxb3mri8yilB/VeNhgNTW/gI58unVTTuOF1IJGsHYCHBanImbKSHC87arj6jUZu
r7q9GtW3Qq5+/dX0brSTOM3DLxQb5ZZ9HNy/kU5LN9FrmBHnpan9hTMtrpWwbXD+
aeRQTRda2yj6l1R/RVHZXje7CbRZACAS+p/qKyzJISg8tnWulPSEI6uY7BOFlQCz
+z1IoDX3A2uZYSfxCKgUluMdjYPz+Lt+yTc16KuFfccFLrzrAyCqfSh8EOWsDvdG
J1x9Xe128M+cMio9i0kLjkrBbw4q+W3l2WYMOTLpwVfz9iAFTXKsDUun+JEDbrjL
Os8yW9x+pG7m41jA8tmVbAvR6jya53X0TagV4JMnN7u5R2OCpd7JqUdmZjpx6emF
h5WjM15Hj5m4kNpecyXS1UZEeZ0WeAHtxjn0sDIWA1Xd4zvjnZGVNJdo+1PvR36o
j41a7xoW58UWkL3ovIQ76oOo6rLZpFeGcwUhl9i+mp7K99qjrEAx5KIeyfH1FbB0
ybFRaak2uS8+BlykM/6hrDgc6gJcmz5nzzVY13ID0Tjo/869DaS1EOl9EGitaSon
OvXp+PqRJahxqtBl9pX+aKr4QkkxqKMgR8RXgQm9YOLmNIUUs/feS9zpJE1/hlSL
JTi8REWfRvIOW3aDn7dh0EAjuM4Co8/n88w1yN2DPTAilBjqmVBnHZ4rt3QKTfjA
j35S+8lIyj/3QrQ3MF+KrdKeePwQfvsmiIpyzxMN6IGgwiOZaL9gdFFz5fOcUxN2
zWUAFCwB77NLXccxllfGCGe14N6QgunDYEWMRXZoQ8l9bbF8zqzAQtckMUbfo2W/
3OTJpr/9AeMfYZJvvtN/y5SudqlUJRXtvjcnHM10bTkqgw2+C2YqEp3YVljiVyc3
uX1j7pDQhYU/I1M9KbvpE5u2KqcZ8pPUJZ3NUTQA2iro4jUW+O+8LHzdTNYF+7zY
92Su7c0GZdzeWlFmMKpcOZQLrpFZ1iSxODPlAYePAwqqLcCoR932ioqmbX8RI4s6
eVNZkpMjVGgUHYHha40QHEt4EMvvFv8nlEr7aoWhbmoFRF5l4ZwFzwf9Cy76Am61
+4Wd0aZBSI72pCy9AfVDPx3KDW9PmsSCJ0FehxGXegmtnyxxgMSVKnLNhDzEgPs+
2lfi1nk3LQ31QwCYQ4OGd08KSKHN2lP1hIj2DgqVNZ2SwMJfuLH/rcoh7tdQAK4W
ruZItxzrCyxqjTHuDXaM1zSMfUF6rHcxheX7sRgcHpYoeFJ1CrJ3yWWTTFq61YSg
qIFbZCDtVwivgD6qIGHVml9CHSPE/58l2wsN4ROeUZof9vxHwykkcBgkU5RXSO21
PjPBrnJgbldU9DYj+DKrYKj95o68mOjuWo6AvjjFc91F0IjahCjFtMOJL98z+hEh
ALruCwHZrZ8lw6YY7cHe+B2BCWAoe0oNE6pgvmE9ff0MkE/bgP9tnGZyt2ROqsH1
6hBdgJY8Z8YDxhqOUXq0g1I+bOgayzmAFzMXLs1BU7QUmKjUB1K3Cg1ORbj0+MV8
B0CJcWCBXvSlEA3R5hJik5aKD0hc5TFOEAIUU62PxdH6QfB+rsY2fxa7jIrLWsVL
yvbM4vLW/0t+A7F47RSlXkkySLH0Qu17ZCQkJxvKS9diGWUe5kfNFvrWKMXErOpI
Kvpb6fRCBbAPoPtrw73bLsU/aM7xZJdBAVOCLQa5Jls1ZB1Qii/oRbP2bf4io9ID
xn4Z2u8VGrNYvKi4C0IlXijoHHvoxSJpnmgnlVgSWk2E8xJLee7rg4J8SUmXLAvt
CYRTzNt7vxFxI1KbUlmgY3Z5lXpoaxBXoelS7ukReGhUyFhodT6yct+sAyPr2DNN
UvXiqHpGf9x/gOTggkesh+xXEKDISrEaLy8KVlzez5cfEO+i0c74zW+muaEeV+ss
wHSPnLG9tfOINyPckBN8vEe37BTfl1o/dVExux9liWd09/BitleMEo6n7hFKBjMe
Hz2aXsRjj05lHw0ZRObXJZz24ktRUkGkdygjHDrYL1laqVASMkpFtrvKoSPEqjEg
ObinHofgKMFKVerLuDS5f1h9/QxiEM/o69wJOjNB+yjNA5Dn8B9DjGNSea2pU9jy
leG/oLULJNtrsbT4NeeN01oKQqVoj8pE3Ee1zUPjmhign5Q4HIqaIhaMTWFH7TxO
0F0L6gJs0p8Hp6vfstq14N010mDW+i0HauBDK+oaT/OrIBY0Bhtn4VHSi+L540mQ
6GtFysha2G2wsHX5MRoeaaFyGAvfg0/rAXzaK6s9VlZQP+nLzTXkbz8og2V7LRwv
jqMS/i4O3pvELJbkxmDhkKosOOZ1T8GL31tq0oulD3dWL9UIk9T4wBgzucIl0C0Y
fYPqn3wzSc0QcgyYoZvvwnkj+S0fI89OphfuBVxyPtrlaH+M2GO99Bvf7osxbZAZ
HC7RbgJo2ZKpdPLJpl8yx2e9y7qmQHQ4xvBlfMpdkvJoWPXnkpK4q6J4BfkN01xf
Io1SXcN/wA5kT+xZnyLNPsGPGiGl/pQ/0SEpLDWDD/h0PRSSA2RBRRBPPQNNTuPs
21DhO0G58cE1HQOb7Xm3bTVbbNf2gr2yu/V/xue0nq21tZ55F37qR3MyI55jM6/H
kCc1B9BTYdy9j0qAtOydenLo+2X9Kv+dODLvyk8N9xLIyi2WU7HCbI9THgUKZDCi
UCpE/qWyJy5WIOsNuQEM/5R9FYSBWAF7C9MNUAScbwq0bILKUFLxIBdHDGm3V0HY
7IRq/tgXI1lybqkUaCFyTUyXpF8yp9s2iePzF1L3NZTZA7uNaMa8lXG6sLXExVxC
KuDk3ejkTBoQeQvysb3u1HASsyz0qUsCMW6MzdJkauI4OzT1aXzMHIOnR0RaWoZJ
veT3Rabtb0xdbZZwVU+8wFPdhEBE0Zzvf2+C6C+8ctXfS2VLQx4lV8ZiEBZ7FZq+
B4zxUXKcCkBX9itBN2CdAyIhJbzH2yfdwISjEvLTaa46V8DSAaNuc6/wkxnx0CyZ
tn/wMakTmcnD7Lmu4N1mSNl6yPJ6JClAikkr2m/dF038c4WQRSXb6XM+s+ot6qAj
5wTZjN/iT3LaL46uGvIXd3xLXESjgHdUlLKBM6UOC6jHO2U67dM2zy0tPQs2VJNB
iNLh35zX1OfxY5jx7hXZtkK4iKhXHWyDt6gQ6bfkBZRZW3qK1pTLyPLLvhWJ+U/M
RfCkSCgvGTvov8iq8Ccdk/ZhHP0sog1btUBWuO3KUhZg/geokybbfqdbbROHpb9p
UHrOlj4EUQqnhNjKHYD56sKYvxf9NkOGqoacrUVaZeVj/x7yd8B3+133BCEmo8XC
s8wR5mko8vD9IekaMqEfasGofBlXIasLbYBdXrPUh6utiwgrgWyrC8mgHSLsiXfa
3xMvvS/mxu6x6i5Ma3wQdtdeJ4pSt6iEFi+4BSscT4FsM+8TyfiE8USYoaN1Ib2i
q8pVaqAYl1F7+8dvd0etuKgoQ0AeQuraG3iAkelD4yt3FS02itosH3fMdMf7N4uN
VHufJCJd3JbV9uS60q6xYdufNsP/t2i3tAlQFOjNlI6H7wqKeP9kGT9K9qti8g1U
O23fYAHE+igEMoboz+qhOFT4oR5RQjiXS0tN6aAY9NEqbOyC8D5zfixPz61tpNFG
C34BCgowdrbFynWHwN6AA3y4jT3ijk0GUZAluJnE26gllsFEYkW2b4VA7MyN2ozj
90eBkopJpQd2WhXVdvDBeNoZbE/Z6safbwgZ1APxscLw7nhWbKnFSdwceTO7kmZ7
RJWnZrp8QwAocQmIPSaUhfMqSG+Od9Kl6NjTDmydPCeKYYVHd5WlLspPhnDz+XdU
MzSnm3yXHQjEU5hTdLSQ+YPGDzVQwUd8607ejx2iMIUZt1snhJN3oC4tFmuXtGVP
USptzDjkM/8ingS52BvUNjy82bi2TfvVTfQ8Z0LTC5Iwa2OhZdcrIE4UWi4VDeFN
xYKASEEp8310o1sMuJQ31v0WGxwlWFEIPOtdwHM+T4iq06KwlaLf2FGhOgHQ2mvg
6bUy/wHWsmbAnwqxV51QMyOqzC+VCZI66xvaRotVd1FMjKYQApxDA0HB8v7hDs46
H1OYB0HfM0h7T/B5Z9yQCF5epAYKifRkwhvdXfZ1510cX299HqLtPzZebitfiFFf
OB+PF9bMsQRXv7PRLPoMtycwDZfE1BHfsBmInkgqi3lJFDXVYgt0aQyXxKTtBWzb
ekcz00yT+ZZpYgoZj5dY3efLrRbRn706y+1jyPs86LbRb8LGTa7UMbd5LrnzcI7N
+jIvoEcuNIgpfGrjMprtOBVDSXiHLp/MOnJpC2YMUx2cW1RGmoDLe/uacoWqmtO8
LFeDIUIXPOGc2oIya0S92sDQRNA4yvHjXGW/qWjpBqpUM+mZ+KJKhNGAWvSl1oqz
TrWFh/4NUeuOJMBiw8ul5avlPsBbr12pc63RRRRT60AKGbp3c49CeocAzxRXhtX7
2CNnWguhSvpU/nmxlKO7oWWl06cfU4oSdKvaJ+9kngdr4/c1/GFrbNAE4KgTTxfS
J404ZvjutY/CrcospGs5YGVcAGk4i9L5jLzVM1D0xBDY1ZSlp1O+ZoIuPeAQsftq
J22FN7IfFa3Gaq5ASdNAF4tLcaYl43H/sb8YtEhoYDe3Fy16DEZGCqvigfWxuhBk
xKLojQwVJeX0FGSTZL8RT6j8N8e9cDUyWsbwP+8JrRvHYDX+u1xT3cJtnGFYPll7
hug2Mtd/nTzs172BAUBYIPdFdMHat9Yb+IbyuNqMJgzBF2rsmd4SftU+xaYqDe/+
0lnGM3Tgr3rQETf2mU8WmZGGdWZAdQ4vC3+z7yPNZI66a+I+363HWxzWfh3GQuMd
2jCmWoypmLqPBpBgpVioW1dCy3Q7y85vL0NRjGDgIrS3rVOOWCkjFE5yQkXctYqm
t0B/dR611A68qja7G/eC6MX4EywcK9vlKnHLgQEXcMe15CUUwLPpcOuGQPKKbmF8
fvCIzOuz0rvND5OidQ1wxps+WD0mc4GuEcuycxAKjCzmtra/6WvnxHko5WDGHQZL
ehY3eNurl5qXuFufyzstzehd2ZkUee8bI10O7P1YLLisOTj6X5ZgtXaNRb0NQevU
C+y5sLpB+lPCF3NIleHoN+lx8wTYjTCHhIOtZmg//fuXgt2SYZ6tYwKq/M34UXo5
TF6iF+eglkMZtMFvZHAKJsR4NvtpFSZYfTAWDIrAlguR0kB2XvAhayAmQek1Vdd3
HKm364fzhcdlFIEMNjrXF+0PExMPrmNXRh1Ad8B/woA1HVelB3EkI884pP72/QmO
LhQh/jscOs3Bcy4EOX0AXLakJDlBQxk6POyTla6829ixmNDNnskEwV8vm0kiu5ds
UtkI9M5C7YZpqBh9iSjNrGc37MRo11kj5FDdT11PjSVnUPyQH/RUyJ8uLx0g1ygd
SnSvT5fhYUv/wJEnT8LHcX2e1SnJ68FRfM+480JfybQklBSc4NDwqKmz4vPs93Ey
RyQ1uu3GPbFpCJF+QnlF0gY2ZX1nhTQ8KREcaZczAYlkPOez3fPYt59PJbwxruvk
V9nM+qiNAeKvReSbG/7Go0yLoRYDcetDaqsuW7EZG0/Aaq8t0hGbtBQnd8OepYHw
NVglLJ0lDP3uJuycOLv4mhyFf1PK+jeEexTytn/CGeVjv7y+ha65xOLJmvR2mcK4
AUdiI8RYXUO/n3VzkAhzYfZjBBA11L4t50hXYsOmL0iOUgy0cLAReoCJ3M4Qztva
CSkrRKtMI1sFFV3GSAhTeFKrOCj/nqHaGKgyI0ftlGDGR8LLfk61D6KKa/b4xdib
oLiKU3AFYL2nvdImSzZmWBLQc8MQfjWgCb9LsnUobW3UoNMd5kWgrQq3LUxUBlp+
pWh0Id54smlwbRBjk74AKkjT+56ETbljbcFtLETzNNqF6ZbFGMnVshmYADbqIkcL
GSZ41yJ7vELO/pHOgDG8vHs5hZGe1AsA5TFIaRtmrdaYCiki5/OnTDORB4CL/of8
K7ebHvJIGazA183caEglG8sU9Van1kuAYphnWitPr45Ku+fbgb3FP2w0E+ZRn+Im
O6Fk2iPkowBFDYeOM4XDsbQfraPfv+TH0nuIHANsAnZki770og9ATa+xaf15Eupe
Ri4++l1TJN89G2VmXufe05kvj1n6YjgRQ7/WKz+jUv1hqk2dIfLx+d0ZSLv/j0rA
6V3zpZ47Wf7RANCeMK+hmf3HJ5YkcWDg/7J5TpJvFGpFVcsD2nrML5kMVeCQFGq7
JB5cb6KjUZ5TdNiMf/QL62byL9eaX5zjS5Qk2vUZF2BOV/gOUgnefxG6xcNjaofS
Sb1YWGIlUwq5jzN4l7LclGK2lDzZS0hW45qElSRJVZ0ZQbaJ5KxxSRygOzscf9hr
TgzVBCEPiqDFZ64t35V0KL++FWSe5y2uljFJDAQXD4E08Q+vgMoeLpZLhetmIRJJ
ESfSwtiI7kQLE8YF0s2TEBJjdDPemuRUtyBb6JXdM1Sr76ip7XjSQRyxVrL1AYi5
OT4ABibqW88jajEUtgbgyn0PUIV6T+LdAJjisxrojwlgQpIUevu++NizlHcnlSqr
kH9rpX2SbZ5I0kRwkL0Nn864sKmR7Hhc0N6i5gdIxeXq3axQdwJKxaDR07ZPG683
JpGa9a/aYtZLdZWjdIOx3Z/wGEEncfxHXjtRQRsTUPFDLHkyfe88XetHqYTJUudm
SmNXwPgca9AGU15vj5L2RLnvwNDczhb3UMXCX/aXAgKORketGUVWTnVO/+A9SJEE
PX0qpv1wad0mGttXYr621oLcb5qkReFPhlWeumPXWgXddmacjZlQly0myjXLPo6l
bNApUEd8rdZWkGyMLrdMfDKLKm8XEVHzTJQ6L5yJMPflmxTy2yk2syVLUAoA8Oly
f701hXgBu7RGFsovpwwK4/U6Ah0+5JR9zwq24UwUSj6LsWqHO34Lq1qAkZkntC/k
gz5IWHfjhj0HZyW/Fkt9hNF3/D8OFIbq1gQvxPZl7KjGpCP+sYLfYANPYZe7EOB1
T8hizaSuwbSi7QbmlI76XFrUYlOccIZWTbPs+0cWs3FBgILwXt7hL7Nr9lPMsB8J
ejQ6TdZ7Y2D1/ExjvCBcYs29FzX8D4ugIU4fGWqmwWpoI+41zVNMsZFu4dckxt2n
uQP0anxbNDEOTq7/ydnsJi1e47Ra6x8torqLD10ND3uRRlLmP9AqQKOSBGoTThOr
3N/5/pcNXqlG3TNq3intFmRYKkbeTAlwDO/KbbZgydgxHAs4sKoAOYs9iTwYMpSX
8Jqj3ymvkLy1VddgRfmA6WNNF8zqduZU1nbn9JAxgRKvcoSBkNlLiymONiU1/5kg
EW7gmtyFuIikadujynoU2E63DgSqaurgsTkxDjTIJITCML/6RUCVXwkqqspCXDj7
KBlNvIz+6WGuCXJzVfzHZqfFJeZzMNtxDI+OM1OpPiA5x8dvrQeFi4O9zAym9DFA
j/etUZJeZvqq2hUFkZYR7LMcr1LmHBEVKLT+AILqpC/W+k8U5IjXHNKb+ug24USW
OrWI1gCs8/ta1o1Y+hilZ8JaDVX3Sg7uL8V2AagCij+f0HFiihjtqggdQCl0Dicr
CFpS/9JXxlchwg9aULa/17/r7qv2R/YIDuPD3nBTzubkX6QvpSEApjou9bEdvkZ4
nlUjHoJwfh3LSR699q+s5TCGPvTTkCFd0m46ztNnlJWV3AEgNPiNAubq7JDUU0ia
J4WwjTNwBGUcUUV+vqsE3DYAoR5nKuCk524+cRjVRf0BttoJlZbImUEUq9gGs39y
x1zAoB/pGnDiN7OhIasPUqfsb4ozrDNIYJzUaNsnyGyrZoweeT1FiGlP/P0mDMgH
IvARYQQRpXsZ2tpb6DHHcN86c/jS+P+icB7dNiXz+D4WlfDdAA7k7viIE21HYvOH
mnModnv/pzozHacgbMlwTdE7oBDgqC7Xr4rHtFh5GoiuB0DmH/8v8/QGoYRE7VVG
/d+Nj/2HjTErWXBms44ylqvbK5T7k4VSlv/Oc99XtW+YEIMYcgzngqGELtX2+u+9
nRpVQc2dgNMSnrzOBlOh4Z39M2gHO6DuWuHk5KOqItteWsMhAkGCUQb3RajhVMaG
blFRJE8M/6oRDwu6BJhlKr9mffR30Lec+QAAKETVun4rpHhN5RwzVmzDepSHVndv
ZxkpRf3mrbaDo+JGZiaKm9xx9DPmSpd7vuJKSnf1AV6h9MJJI1w4NU7qrD18jZN4
s2MnfB5Mm8f2/U/n6rLTvXM5a+Xkj268Kgn3veaIZSZrMiGu2Wu1VqFmqLmdxs9I
E6I5e3Oj+RNsIYe42eN1MM5BNaAUWRjzc1XsWq53SwIJO7RCeac1cKb8UZQediYU
8rwOX+8GYoqJDr/l+ouoXoIWzJsksl4bLzLB4nVXdLHH2ZCjyqgXdC3N37l6eOvX
Zc9FOljPwcoKnzAV9hZslTRrZMqxU0Ask9e4iqvVDzB15ZbwgXWBmbYNWmwmypoV
vsvI3dtDyOz9f4iY2NRwQE41N04omb3d1TMG+RqGdqwGKmlPaJ1KTa6VPM5QIwnE
BqMvUKm5hYfqB0CIxlGLvqcOqLXFSmILTbPEZ+pJ4UTUTW1qTgVUIH7RzKK1Sqt2
VPpsL50xR3SLeL1zyOOg546BECGM+4Cq14t1ym3gAl7pqKLS7mShqG2s1YkRWu63
UPelMNgeCNOF8EXJ27zdJt/t0sUb/9A5ZmzdwhUCBiqhRba6IcmeJFousm5GUIXa
5t5/v3z03/tpC2tZ4sjwXSmgdjyAiR2yvDcOrnlNWymkSpbnUSfnKw1hptqCRsI7
8R2NgycY2z8uzooQn3/ulxkqsOFh19eJR5zdsGlGW3l1bkYvcSIbUCgXz5NY6xxq
6ONomFPx7IDj1qTskO/7z6rViXAFo4Heyfs4k7juP92UeX08fYTRn1VQjr4Uw/h8
n57kBcPNasjEMJmH2L3n2z4cy6bf8HrOhIamsyLSb7zFVGQy8lbK0YJeVeCvpxvC
ULlb20lqdjz1oRQVsvzGSnB+TLqpTbW11E61/KTTO84xMG6VMmVEUlCJOTMJ6B+y
esNViMFvmnsQScRcXcebbB3JtIF3fkJA+w2suLgHvUnh7G9w1hGJ4I1A8jR4Eumt
1Jxj8xblzgERn7F1r3sb0M43HpoBFSikL4ATP1b5gmufd31X7Xwj3TdgVPKSP9BK
pVj8mSfUApG5KKxMUP1V6ayhb0eI/bgHVOmSV3BE3+4C6/cxTzvJHYZ7SvEj/Alc
NVfB1jQc1dql+Jis52bwVSOnVwL4tZOiKH5x35BihyRLD/i+5RQeJf+/lbAnVtDH
t2GVLneGzlXV2D21R7dNRTryM68wIcOK+o/xmNkdqHKrM0eQQ6AaLrF414I9Enb8
e+FzdeGjStYtvNqewOahNQy3LpFuYLG/QgKRrWqObrlA9QkECPrZKNSLg1CWd19K
TcTk/RS7JQQruu5LLZv+ke6+bQbyEyeOIOyadIwFz1mNb9lYg9o6RyGVlkLEYkUY
homl11jK/qp3HNGHGtTB2dYPEl/vy6KAZJV8xnQhERM+AdXcAhtRkVSIDD2QB3nt
jfLSX5tdKfSbJ1NskIF//DGEK9pSm2TLx33wjKCCl4LI+hXdHML3845/WmHlP4wE
dX5/MMKKnitELS/yuth/o/km3nC+5Af9W3rfeHiM588gontZWy/9ScUS04RhpbAx
x98vBLQyDW0CA4hsibAJvWz7uWb20Piy+yoNNsYK7VZ1X03hq+aPYNdIbBv+3c2B
DzjUYNwY9+1NgRjGhbPfrxv2v+O5M5pYY9+/qe8NkBYHjzFjJc+3D5jtPTjlp4Tp
vo/IMItDHOZLhA2giIUiaiOEWGEdHmOVXB3Rp0J3yZfDelvAdo8NN8sIbdLDGdrV
oKPSWRAB6Caay+Elgrg5503dP0wYfqFTXmK+9D715/t10PaDgXL0TBqCASEiFEMP
7GEIANd+S8sSQu4aZ230OaWdGOPzRk+cXxqdwXxh/gG67V8wpbJhGKb+V07Cbzzb
B+CVtr+9m2bk9MTS/d90XVKBsfb1e1pfVTi8SCdahv4yfR3BTUk459jHU5t+UkD+
hoY3qIwpJjYGI/p1zmiZ8oTfpqPSMcJ+cc3ZjAnvqUmS/DdIjZgPrHgJFNxoi0RC
LxYP3/BxioYKHynQSnWp1j5rnuhLppae42QId77Q9gO+0/w6XOyCPIF1JkeJ+SuG
hePQvPpRCJOVC6scs9KROKHJBhdxFIJ4YAy+MPgDN7CpUh0zxEaXqAluNfsGMmiT
YlMXhqpryhSKrwLTtv0ymzS/1k63o2hbSFHJ84KYWZi4FglZWtXfIWivkyVX/Iq3
QjCUFE7VAh2DrPpjHuoMRlM4YH6wtwvo4yW9kmoJmXgJ9pLU2UshGFkbmkLeqydO
qEzVoXorJOuGOipx6wePgOTpVcw/zJqd46nTbFPOkM+PNGpKN3UPDM7SIqlSh2Ls
ejXmvKQ9LgSbZT7qD5C3TuJ9+DcDmfykOB0j3C8mfts6diV0YjkbJsMXxlPXjjTZ
KD/nSh6BWnDE9F67TT+UyBHty6OR6bOmMOLX1q4VQrjwbSc5yMbo9z++WPPMOqK7
pXZBT2DhlGDDsaZvTksV+XRQOuk+JFjXi1tZQIODV1xoKg3vYYEmAICWA2Zk1ger
bsLGl7pjy2/6CtifzSx2a1nZZPUgv6EQ2aVti6TLrEyTeXPblorYS1XXsAC3uBEP
IYqbwnXv4kUnhIc+g8z9wfwGSpj/yMeawy7m+1FjF6bGVowcbLzvKt7eARP6Afsw
PgdAHrWBbclgK3etCsJ3t4fGWdIuYOnMZgl3mpyJB6QAJjiIi8H0QrYX4qvGLER8
vPRPQTDuV07mDNPzmw9vwYZ5gZa2yBLbK0qp0uFB7m4AxV7GmMmK/HkzsRkLXXPx
d8PbMk6LGcq6hLKwoembmQFWs8R+ac4A6TgziDjrYnxS5PoeZlyZVfDildnyIJtG
jEPSDQc96maH4v2DPjm/DjDKrDeOsn/hOWzVIs38YiUwC4WfwK6bBTfMmue/MUOI
KfhSXwJQ52vXCnzBSQtdskHcg/sS5a0TVwxN0DoE3h5d7ubAJbM0YiRhXAhGdSAx
RJN96n919lkchYn2tviIR5c3EPnsPbijUXCJorQs0H7tlsJ8Yt8AtL7zpI3OBd8B
IoS1dvnzI1rkepPdTEzxPCZdL2u4krx2CPtdJvBWBFcyt9Ibpq6srQJIdclmfl3u
h0auqEW+PhLEuQTezQd5D0lWLh41aO7q4j88GMXAUiqVsMckSU7AYzdKA1wvkKdR
ga/80vLYc8ioA2t0FYfesNxHt6GMw/LrQfBRK240A5iZ5jmlg186pxpCMTrQvXcq
IejfXFXG7CLjXcZMZTgvaSB73KEQHUmvAy54Xxyty8ONpnYNKkgggE1bxf2PoeF5
mzWzkP/h5HtU/2Xf/ccWq9COAFjeoHE0xr9KNwlz4BIvjKiBgCe19fYK8lTPbae+
kTsh01bYGgVRspyRwWyrYpuyPFf9wAc8Cboefehzkv2vDgtHRT4azMJXUxgBL30j
AUF5hUj1ixEic/JhsM3kr3EyPsF1GibNaPAiESC+fQklySTGGqhQ7y6a7OpcTS+O
XXEd524ECSZdeYvMo3JhvTGoaAwJzgqaOoCQfijX9j250qh19ksH1jLYHXxkJORX
pMkczRYzoF0Q+3oDByTojhxiKsGgvPRynFYiNnJFraNxnYWzhSBpjVasbzQuCGJ4
+xnkjTpBOFjRb+21PmuZJ+lkygDDWixu5A+uoxSrR5DINDcPpYhzXPVDfJ6VSP+2
BsdOWQqLyU5RRurNxptPVKGHn1RiTSlVYFbeoyoO4rteCKyryCOalYUyXnZ8N3OS
hHHlOe2MV0wvmUb1Goe1/ouMGleBoXSAdzY/x/1NNl8wK478YGXeONZ4kVfr4rnv
9hR+U7yxCiPDW+nL2+rV9jXPFNZpAQUC/m9Bie/Nm0xy20UsNBHryP0MPB0zIhRV
C4C8i3HGidsrGOVlNELZYBAlta+TrNKjQKrYMjH2MQNQVNUNpQx2gDnCbcWwbIgH
5l1iOMkM0Nsjj7x7/INBweEM9N3VQZ7DLtEl4rOVwcwMLyn/v9Dx24friPDW+JP4
WluhMIZNbLmBpJoBJQZeOJPB3srNPwz25orAnQ3OY5uPKH4yDhJ2lKPEKjfzkwH+
jXE97H2BNRx+wcxBgp8OLwwO848hjLwrB1EmcywVzSTZF/6miI21X+5Ku5JhCr/j
TZYnv55y5NIhstXJh4ZiUcDAvF/GVmdzL7KYPc4jkuUjOyARCzA0abuig0VNOkdy
eSuKYuniuLiOHeHh5hKO0eT13Kj8qt5h5LHmK24KPQFGArPHqFh/+7mSCY3nax0N
e979ALahcqNwR6itv4Wtky1seDPrLlghhxHloomuDBUJETmDgcesKZva/g3YKDr+
nlxsA8MaRY4TnCoYr087UkuX28yG87gSTz/5kZx+B2LiylUnA8KN2aCafd7Hbi6b
1vso68Wczz2OoDdhmgzf64W0+28/zvyQuVyFpFuXL3iT0rv3qCb+rhupA8XItMTe
voQ+xyxur5KA0I+X8RqUPlESd4nMWB5M44izy33+jI5gi/pM49XimYoL2TDMzaFT
hS4vnF9y84Z8hGHSv2LvgcH1cHKY+C6u0YeGAG2i19R3rUpGuuLKoDVC5x1NhxWk
nhbmCcE3vIOKP5M5y8QsezmfrQlf0FbR2iQyoqdCQDtzR8f+QCv9lltxzIIO4Ubh
VXI9ckhoK8TwQS9u84OnxnG8zJrnJ4ocGFUCZHaYBGZAg4aN10HYZBmWR5/4y6DO
cvOBoxOZ5Rb8hQqaXrKejz+lWMZBmdpHUiECRuSq39NX5RGvfl/bxSWHcZAKAVS6
0x9GIDZoVCd458kSK3eHl4xtGUiZtwrybdbe2O35ncT6xzQaUVrPhgUi4CSH8Q5M
aJzYp/lveaUDHpzgypARSbopS+sjrYLDBlEx+lsJSo+aXTr/33knwKVQZE1JDBN0
gouDj/FPTVDcE9TkPiYf2I2fDVeWkeDVi/WLR65QdrMz1T+aBAvygasvCGssb6XP
GvsDqC+8QCjbOkd7jfnNQjtJpgl/b6wXfR5P66pjXrrS4M7079PPesc3VDF/Kv6J
fZ2fqCDpFK7DbOM6E8r6Kn41oKBVybLEdPz5bpB7a1p63GLroFJ8w1hS16WokozF
oGcn6rcfdugJS3us8GouqAt8WW2LeRtMxb3pMGxSJob2p1X/MoDZKhzBhFf2cn/a
I7YNvzEjZw2Jyveo4m4paOKBj0OdsIe8Uw5Jbi+Oeleq5fiMBdOyshS5Ipg7s5jM
MixgR35ZwseNuCIaGf1j7J3LfFj1F6eWhDSdO6+DM6jZw/3GhXhP5w9R9aGhNfIa
4bmsxMPFMiGWAmnUn68GXef/hIZWOOjUgIw9PPTgvvN6BVwoKJtIO5bnUdOpOfNt
vYjBHP5cK/mas5utEe7foAWSCmMRbSifeGL4Fp61xC7t5QB8g2pozrERs8NaQQup
JJJlXNitFpfDc5YWEI7ICfESg3KoVpvmo8731b+B1/pzVoRimFJYpAUmfv0hH2jF
uderpOObcEguTL6ZwD/UTv2NGXPQMqv3fLQGoGhrMj3jj1th7uVOuUqH3PXmQFa3
Gy/jccGDiL1DdZTo/qbQJ4CTmW+vO6QLDnCBRvlmIiFxSg1UtimmWIOWCoEYCN8H
qBMbY6qsNPbDV91bxqGdhkDUHg4A8XpVFkv4nfxDj9Yyyu6xJEnlgvLfaNEZJX+W
9YcesNl1vXbCBrMRcOWZ0oGgXj1JP0DN+MP+Q3jIPhp29HNcgl5qyM2x34scbUBn
2S64UOutVhh/6XLsxuiRY9fEdfdbyqxA+o2invpUvefUu8hGNPOublWbf64YPQY3
HLWnJmVkRBS/0T/+oL7AUvxQGPh9Lcf9hPmW/t0Ew0apmq+rVrj2m1sUVxCK8jy9
xmBjiiw4BSzxFZAYgUDCsK4kzgMbU15h3IIpJezxv9+xyiOiQtJm1thr7IwtaqLW
VsK9jD7RPJcAr3u7G0f1q+FSIcBIAqRIMNR7rltG6FLhOvanQxcysRyrNUS0f0NU
feDHn90MeX1FFNlnTXGWqWL2t2yTSVExAgMmNd8IeqEsvNs0/rgbNpCAENY/Z1sl
43BsAn92i1hsBmGGu6LO4Vw1KpoGCChmIRrxIO+1/j506RVl+CgR+PdpYp3AVeaJ
KAoLE/FnXB5uHwfiRC3oOLqa1VZRmk9/Alob9lMWsTbTv8ajrvj+H7kxdgpxN2/8
9A0pq6XAPefJU0Yu60RoGA7ItxuOe1uq7OlrkpFoJ0dMafJMAAfSA3LJ4K0SGlVu
zPAD2+nEE8jgIueyzmv2LL9UA8GLtrVOFWPWFmyYczirqiUCu4hbrsG03ftKqasq
qj4Fxfb/xdh0i4BiHjXOQir4ApbJVjX3fziv341O0p8aNGX7iZ7uMZb9RDLI6Ec5
vE9Z14Pqps88Pt/7Qh32k65NLtTmdDWF5jVkpH68QNctWjsyWSwGv+BgGvE5YTk8
QEX8SPfD394eUPK7W1gNfrKhKZmi9dJuwXjI/PcKZ9ED6+Z/VYggKU46EKu76nUy
VPjUTQinmx+PueKOPhCXAzILaOuLHmC19sCJhmg1js73yy44SjlmyiOps36bGfGc
RjuPhCP/a3yHUkWvyz+l00F9nlYoB2GRhvBc7RWJto3jTCzdP3Ia1o1Y5tcfp3QX
y9XcxLcprQR8pivYsNFwq6zCU0P8Z6uLpypY6FOXkzfy9Ru73jpAclZEf89PppP3
ISfKdyAp+ve4Qn6gOzY930XXgqPRJwGM+ERyb4JaSU4i7yMkXWQQq2kFY2jfijZ7
fWXZjd3uM/GnAxT1UYLMIYMp59BrEey8Nnz7PI8vqHY90iMxhQ1ieyv8+sw3D5nW
xYWm2UwO2TOUcvpAx1XdxAOGV0IB5fpDmNtp507/pghkvRpX+0sMzEd7+eXyBvfN
QIuCfjmMRoX9szpAwQ+R9YHT1e9PprkLEd7QJZBOzebB9YdgZnMfId6smLnOXylk
/NWnvAsMv7kw3AtzVCB5xHr9vmjJ6fudt50Mf3RY6Ioyai59TbCy4A9RLXkxKNJj
EkRJ0fdeYYCrP+dPtAHvbdvWEqHyomGAZCslvWSo1wyFwxOFksLSP9J7TmDdmBMF
FOk3CKFxly8+hZLhlrkV+3TZGrso5Z7JpGkWT/FcuqJvd9/6wxAK7kZreD5XmqYT
YEKTYurojuetoW28rdN0gKBHLBwuBg1A1cDTH+1T6ogHxq6+6JKR5WVDXS2sDG1u
L3TCJRA9A5pl7VOQ9oOxZ/HIWtEPLg7jdE+Y2FlyrIGe/9LcYtBKSDUYLb3ZY8UE
r0IxjSHjN3CAnHlnyuCZ4H1oOP4ldDrWD4f7QNG8l4UeXUFivO3RZRZw60nu8N1l
/qUmH9RkpYkW9zRn4WLLah2uTvNYB+8fptMKRWTPQRN+rdPC/SP7bKMPLZkGyT/R
hA5RfdqcS48hFRtEmy+dDVCfPJJVMd9jUGpGNZXLJUGGrG2+Dsq9LfU33Tpra3HZ
dzWFlVPAopYj/x9uYqRkvRAV4Yg0m0Nak6yi8BeCsCW0wcjKa/zJdQo5bh5umgI3
byRyimw3xNzPGbn1QC6zhPQhUA68yOUOyYRQdc05qPg4zrWS4iqPPhb85x40xpzq
aPdLNF6P7UenqNazM8wecZ+yF7htSDYBazxDfOxRCDRoITS2EGj3ZDTt5M5XYsmw
f28HqHeGQB6MkN/8n6WPhne2C6RusPZCY7PL+Rufi9lyy0vYH+5Ct914A3Kw/UXr
a4ohKW+h6q9kYWW9Gasb20+khUlqwxGpBeos90SQLkBvTr6tji9ZbN20AnQx21An
m7eq4mGCzRB0L/+xoUSQgfcPCan5TX8a90DONZQN1WL0Hv7Ig4tgZdWBcd14os/C
SBvv47/20P0z/CAKXC8QdYRJDnNA9QeNHd2G2uUdLAvZa07Jo7ltEJw1/fUA+Duk
24xm3Ct9mPXi23irfMr2+i1wrx0bRMH/baYTwJ3fG2QQ4ZzwPH6OWID7z/M2U6SR
h8fG30+udtHZh9zyL7MJCsPrCsMCRMDVDWM4OHDZwqXYpUTKXVeKKg1PdMtsVoZm
kkzwL+M6FBzZr+io0PXX1hJUFqEP3YXX28V5VF4A/pxzjF5Splcsf5ZUWUTAhsrC
fqzTtkU47z3IyNDa4xSQWmYQtNuDzxZqjSgWT0fE8IAu3iBVxHBUXtOjj7TFeVWb
IExu/Km7sJO8Ygn3TlI8q8UiOqPmIctXVpR3XvBAAJ0T1S0peo7gW3Mck97/97ZE
4gQltFBytjjR8IoFmyajxgMd9bzJplaCLUmonpdonZHrStCqkP1kPYQgRI0X3bPi
nLg6Z9144h5I81Opmnlulq2QnKvMdqSagFFydKJP/uHi960T2JPTkeKRdcmG7hmm
L7D9w+jlDAznKP/j1jlI0Eucqhp1vWyBtvakQQBtrgjGAVSZarQg6U3YUoSiG0KL
ma7S1wrpWvTW8HhSjAzLv949Cyt6UMtior3xn2JMbeUQE/puCoyu2u0oqdPPa/Ec
rQc0cYgrAFr2P4s6deJMREMaaU0+zQUJZ/W4m8sLgWnLm/jdnvjWxx3jyH/7xZX/
7WagqurApE5R5qh9NfRPqzDF3ii7LRka0t0qiNpo0Nq0NMaQtjgZEtOeWlge/pZ/
iW71OJbJHtQ+hXBtX7loisdn2W14GhK5KNloSoKWK9NtFKvodzCOnwmhIamZ75VQ
AoIaKhA96dq7KMhz8vPEyEVUDJhzC7kmOH3RNeig2yAHagItrAYgoohx4jVAZi8t
JtUTHKDsOogi8mcgXIM7Kox1KXQC8J3Zpu+ruNVE7yrNvnNotNMetK4/gpZdZ0tg
y7V+cHKTp9Cy8vQBS6SnF1tslXAVi+t5Od6byjCuo0nkTDOh0ktxH/092vIsAwHX
Wl7b81tgjuwWR++3cgrvLEP1vcX54K83n5wkUkUUy2QSUR4TNu7sK0tW5w8Q5hie
CBwHBW3opCtuOu+aPzFS80mmm9D02bQUtjdgZpqibDJHZr7RzBsJEntu2egNuOUl
kws59WjSbT8Z8I1F71HI3VxZJLkohi0DADBH9CpVYKJJS51hVNtM6uGXC7pSFXQn
NXDcDt9e1w2SteledpINGSIvehK9Lu0Ez0Y3lpcy2hMhzaHejpHCBviCwVnnZFBg
4D/gdeJJG794UGuNa+wcuJMHmHYeWmVXvOYHLdAcwVc+GbNXg+wUN3DFuerW/+bv
RSChd852/wRbyfrOqS9CA/46s47QkUogxFHkntKT5ZsPbaimyTPDbhasqsLbN/Ot
Z41yg6a6QO1FUjQCRfjmqp37Q5NTr0ZaSzn3nsmQ2HU5UcEo1Wuz6NYk7+ttHsga
HN9GSLM6nV62xp0P/SbE35Ag4u8eTJNeGp2n/GFJVpSHJcCgc3BQi0hz65zDNjA2
/miFgCSUjfRHpHoKsPPl2DjeUzuZqbEZWv4dH52wXv5Ss+o2wBSXQ+V439qkXtEy
K6G/50k7Eh7yT1sv+k/1r77BxZvIx2xgovW9dHIoTk9MaBVqgxijOdlqwhVF031L
Gmr6gY6fWEM/Fobb5eS/jkARfOVC2WFiwg+a+NqI9R6E4Kwm8yqOVKonZIiyCxI1
MAUTNp54uCqP3UnHAXey8/rD/jwoui1SUdeK7S+LF0Fdz2DgHh1fvHiMhiBT+5tQ
YsW1gHAeSuALMgn5n0Fd0oCY2pKvP4EYMH+gdWaTEIaqa857ZpIx7iq5US/mRWhA
7zVukIWZx+AIAg5tg49TTO45wGxPT4CwGigqbae+p+kzsS9OZo/MxD1HbfAgjt5c
C6mpAheFbYzQqGto+KfX+0/tcMy62BN7lr5YbJfzmpU0WDYQGjJ392pJVn80Alnk
ZFaDfwsLoZ+4eOG7VV10uDwzb+e5iqIkpCmN6vvtgP7mLI1C9lKPYnh1qc2bi4gl
vuqyCo2jsAUAnmMS3zuoHNMdPS7+kgcHP1sgco6FQ2muC/kV7j7lcEko4VYemorl
R9V1XAFygtp/K1DJoAoeKkpp8geY5R8yvS3oBTB3o8MFz5QVW5GvuEkazhp++1T3
y0HmYHFF2At1QLq9T4X+2K6R35xLfgVR/MchgBtJHB21OwECibAgqG52CpRHCr6N
GZeWHwdqaaMCoAhs3Ee/yR21ryqmf7be0LcKPjpDAPoMscGFuS25j1KFh+rnuyl5
ce02rm8ymHfJ1/ox0aYYxdXqmQev+HeUzsE8bPly8ii/gBSRp9lmwhzxrnQt9gUH
if/LGDuN0YWitVzVNSNyMLRy7VcANYY1L56aU2qi1ExhndLYfF/FAMYJzrBEkDMv
rfY0GtJt0MUcMr/rge7bVoEhrxPCHHxii8u8bhVlXRIbjzVHG7mEivyuYswQlRmH
zyUDO5OcaYU6KKxCU6tJDSoT8//voGmmWJ86LxvcE9E/II0ABhW7ExxHwj/F5v4Y
3/skYCU+fwGirdA4FNbnUiUaW33YhT12SxAUO8zhLFyUh7vs+aahEgBGRK7pYrWc
gvwk1kUKfse1p7owrdbMm1P+kc64x5LRtqRl0V3Vf0NJrdYOidsPwBnU/rfR2H2I
HaB+SkkNbWqnv8kXr0oSHZTuhGW5v8mxu6E0CqpP2v2NnYHTZLXxiIhpE6wCq266
nzM668/Yv/fnRj10C5uXyDygUV+bW6mgHqrTUZemRfwKwLB7ug+AFykab5MmMjTb
cVBlYUeVqMy2mizzSIehkliVD2UEFbdcNPO426AzIKXyClMrvL3Za3NqAnA+ntcE
na/tns+wqCOpSe7Mz+BGgYJAeRQ2G7Q9TrJ7ioQiljG0Qq7QHfQh4IkPOPutE8iU
w5CEkiL+HuWw5GkJXLX6MBmMVg2xciwFugpicClwb3D2yg1ZhiHXmC0LncO5LgA3
cdkvkljpwFEsq58lXH7U2CgzMgwRYPEBaSqjed61F4rMmvK6Na7j/RnZvNPg0P9L
gccBh6zMrEwz9wXoOBXBdq4i7lZhXI71ZQAoeodqig0HqJ/QMBxauhT0yKdln3Ma
Tyr3DDf4Oix71h9fcToYL/Unohd5bpTrwZJELnX/mdbgazlM0GZNdtEXKeVZyOsI
Yoznj1qdptUQnrqCQ2mcmB8Y7OLvpcnxfUZIW3nNLh2Ed9acEZc2E1hUynTJKeV3
9K9NmtHn7KcfUZbq8NiaooHIKE0k8E+6hx0TUzydpfPXRw4ze7S2UOGbrOITPUz1
EOpAFUSsY84dlE4MddgaI6C7ylSrz84F/dD/JYPawJtGfKY+lNqJ7TJzu46bjznO
MWlUIp51CcMZcF4yodtFsQDJK1oGy5N8QwTlMPfEhxi/Ba1xL/DyFoKB82eW/wX4
9O26muYMniwIVlNFs0i12RB07S8IEleM2ndwlZNkmhohKuW8zGTajusN8/hHe86c
JRXtbTz3dsii6RC1bd9ujsjCIgz3jtRiinMXE0PpGZwABc9pmcIPYY88miF9/0Fd
yvAkeEzy05Y308BtT/U2U9GC7Jp3eV1F5NaAIo2jTN8sUn++Snr/FlPJ+a8P8X2W
1btkYGg6l18R+CCvsKsZWy6QmktlrBEVn9cjCPg1341thFvfZsIVE71Cd8asx451
AFGyJucW7ko8Hea+lXolTTZAIr52A7SSXO9wkyzBmz38hiAXubm0aIKDV9tgjYcj
EDQeyJz8Eupp0e+C6kMMwWSCSJdcK2y9LTOk5zc1hrOx4/FbsoqOI+Xhi6F5cYO4
x2xl+VLlcaWVBml4/YBpjU3xC9cbHXcYTSzH/p80pQ6EOYGgzWBn6f98Mt/BqsDf
vXb+40cKKytKGqF05uEWIO9ds4KW/SjDF6XtvTm/gicobUBc+2ZNp5pj8nckQ4G9
u/99mLKqdCVIAqEPjmg3fw0ptkgpQWrEGGd85CG+SE788WBnza6BufHCVaiasQGp
RmK7TxYFrkWAL1iNeYd1FeRdFiLYkWiwDHawISZ65GVsOnpdsOhHl/VD4wsjFyad
MInd0bfm3Mybf8I4wswATu7N6pKVzpxTmIGxg7xfxHhVsfPi0JpFONCfD9/oX6on
xThuDsptZWYTqZIyKWLP+wgnBEJIha2goS5vUziT3yikfMP8dKbXTTYHclyayP8N
tLCJuQpC52c4yM2mpnRAEyfmSz0377VJAs7TvZBNq1/KFyrkQ8bYrlKhW9QkxiVC
Y03tujT5CVQV1wJSF1oH44nOaUtyfTRsZG1GE8K2B/fXEiN7hGUbPKyAxK3FCZs3
wt7kn68/wHO5bEt0E1b6bX5TrNJXmd97zPqCr2uN+EX5A9e3GcXk6N8UPp1Db7p4
xAQH3E29KjhSAJPOzZCrF4o/lMnjLVehgfcI6wRXueZPhM/zyuWO9ZER1mGIzoVt
K3KccZz+nMNrnWGh3g4PchVyTK/qhQcDCi30CKo2rWLJep+V0Rtw1FpCwTnsRJQ8
P5jMJLuiKGhZ0kp/Fp0oLi+hLSNIj5iZf45bQWGU80AHO/JfOGB8/Guma7eOW/5t
+vGiHDYRclzgkIPoTExdfbD/2ymfLEFvuTNdIw2ln9L/fH/yKig+D97sMjc8UAof
mJ3ZlVJXdC4O+OroZ6JTQiT0KIMBt1dJwmr/azQOl0knCABZ5jJTtmh1ai/HhKLE
Vjr8zj16/vaYtQ+VTbhoKM8Q9aS/QMEyhFo7KDuOuRu+0kxB3oJX+4VNYNZaKrz5
OWqzApqjWXYeuXcx/FS0IygKmMglaJiaqvH7NsmOjXptuFjFoISXibGxXNTBH4xP
4hUv1TuaS2qcnt73DfM+7QfaqV3D944rEHJRHWAiWouMbL9tenebg5nzZoD3ZjXy
jMGeRbKF/v4crk4uAIbo/g0xR1MUYrZtkln/L1w9DmMCubMlUOTmbIFx8LntCg79
x32g9vI+rLIvMbQkkZeBIkHAoi6sCOq8QcVcRnxR5L+QU9mbrZ3rD0HfEmyIVjuw
8imDt2bztbpycc/71UvMjxa2h4wy8i++vv0Yn2qHnkVWZM2jp5hbM3ElQXULCQYI
BaU6RtzTbuhZyiMaPlXvJgLW8gM7ljoA6gDp9Ivp4hglUBeL2loDFSVj0M/xZvbZ
2XJn3bQ7ofNCmdd7IiuT/9Klt0ioJsG5NbUnFlYDyviMKd/T4oc3VjZAh6fLaEKV
FoOvx590Tghgf5FrDa52Hj7y8k5i+0lfLFIz6TvqDoFtDei6Z+S7T9vH+1535Vwo
u320Krm7jKIOExfRb3Mb/veVDt30HwtB3pXDBQT3MWYHRZbPN7SecDAH49TZP8jE
u3BM9fLYX1WoV4C/2XSBWXsdDvcMVIi6W23KC1sy8ZbYSldbiO/Vzti50JaSaLh4
5tldBUmKeAHVbi8qcyTi0QIqOJYRC7ysI7phTRvhCnlA7YF3LSpMjoeIU+YhtWSR
HpOXXDiIt1lzpQZZo0elRAP1argv0PRuj8THXJP2+qxSVMq4oxsCP+vBH3Vet7Fy
d9+tGyfp5yfA0Y5rNrqnp+um/omqsYlJ98FBK97d/WkE+Tv9aRX2G5o+3FIU9HM0
L4h9RofFmkLJ17grYQfAFhIEfOJEQbjXawWjTQhqMbP+BTFQ26d9ulLubIDVec65
iUZ/0xG8SifBui86ytP18sYBTdYZOouqPIli6mNRTHMALUCUOOuLFhzcDCZUIbum
+FlQ/IJwGWWVadhMz+S22OWGR9zZKdmErAlox4M7SoxOQgPzQ8QDwSbTB0kBqFyA
UtPuEJERodOsU9hApwdKrdi1zggsY3RhVc6Dw0npwbT3qlpw74mXNczBQtmHPtxV
P1D5OGE4oGLELiKJq63mXpt3xoUYLxVo3qEos3V5n4AQT7V68Kk4fXHgPBPiVSc3
dpll1/47oHOByyNcjRRJ/QQZ8rYa/zD82l6SXJnxnAtWU0zMbJB5sIcserT4pWST
/jaW9rbCjqExOokONoMqsC2E3B2pL08wbB3EStJxSq4hF30wnNJdt35w/m8hd8TB
C/YANXC4L8sVWD2Psm9RbqZznlrnnYqe8ZLWxpoDD3uTMFNLNtySmy7MQtMBVq5b
v1fVNLy4Qw6ZFY++RTjBL08PbbHkNhD7eZ23sHlEwX1ELaryenBGpXU3wNdrNKvw
BKBpHUwJ4gqL8euZLHcgliHjCeOOvmQ5xSpjp2UJ23tqQWuUUHHVJEAUvM5VcreG
FnhVytkhruh3Fm3GCyKNHIVR26ucvcH+gHiQzKMw3dLIDhWVA4K0vQZOpuoSkzfz
QBEnxZ4D3U4ek06tg+Qbk5afYr39GjRIVa/H1jRVspdYHvqEB9zl+Ukg3NZbi4D2
ZmpuVajyygvrwg7EYzvSOUZb07ph37AEmoZcEiLb/iIFnvD+FTK0C+8EPpinXEto
K74npb2COiZPC+VrjPpoMj0Ex8G7RodqATUGp+1AbmxL5sdUFAz3PsWWwmt5uy/B
JrAkYxdkrWa+cyOHaKeLGci1spCCFq9qNKisi5dag/uc08QGZCp7y0nonDzK/XyI
NPNEvhU8VYagGk4/TMSwvB6vhYAkSH5B+qgMI5dJJ/4mN2A/RWq6GbPdO1UJqvwD
Mai4rpC90pT07vXqvnnnQGZq/npfelcg2EfDDJODdM6VSn7EjHZojGKGRtcu/u8V
IlU9A6GEtzalV61UBZWVecNgIHjyniAQz7qgIj3iRpfbMGdowtKxbH2zP1TEv7Pb
+Qi+aTogMvjsfCs3tst0KDK/lzIdMBykgWP6mMdJ/whVxrxnU67rEp5SGZLzGODv
q0YF6j88beU4uReoOdvZycFLFHYXzOsBnKlQQtFTpYDUjaMkvB1/J6J3QNt65RTU
7GUvcpf0sTnud6JRS8om6ijRBTxVJviW8MdVse1jeyxghyqwoV4C8dOqGo8jjsZy
490O5ffsUK90AP1Vf65twRxtXMV/M1sl36ACssdJ03IzS9oZr5jUsNFXCBU19UWd
26OQArfMcKJGhOlBeeQ9FAqZYI1w+/lfVBIOpmaOZb6JYbtCaVKKzRpvqa5ugT9f
YCQBLROfuLrAKnriK3nqGUE5pDSkHEA8mKMsw6VdJeA2fKKv3TbqD6EGgtmm8Tlg
SfERx084EEo52xsJueju0QSHPIWZ5E6hm2WLER+4NUNeYbtD4jt4E3+MO4kCKNx/
U96wqW1q+9w9MhVKEBJ7o4xJzqWsQUQ1R/DScPM6/w865A6gvZi7PHjOZTqBM0T9
eG4d2nc9pDsAX8FkPEM0v26b54IxHhhLbGPZN+HuWlQzYPMVdY7VjN11/nBeZuDS
lo4d4EByupIDcJqd1eywENqERT7dY8yt7XbF7kSDzbEMp5L7OqMOuFdWo9eIqWvr
HEO5cYpMLxm3XbE44Sw++FzH3ya+NTfYl+3UFXgbeltQ9dk9Km+rUfxpJa7nB/zi
9wkXciqI5P5RosArUbI/rTspuMh0iV5v8sPZUh50Z3nIR03+z5Lny5vmZm5r0ocM
3TcqVoKnRMvkSci1KTieVf+wmR1bgLtZoxdy0OS8GVkVLW8lQNpXt17V5GcBzDxr
VT8gxCfETaXEOhupHRGX9EfDl3XcSx1L64O8tq4pYrnLTArQ60Pf0ZAjGAj4jMNi
WZvURAe5Mcs7B9k0q0deO8SLrDutDRYpvwWoRB3jR8UY2hwjtNnJNJQSxfE4FrGS
LrpffVQXPClu7n6NfDO7uLHlYFCErhYM078gHYgBtBJSA4BVYuW3xugd67KuNF55
9yT6jb5GDuC8+vfpvOorHZJD9IDu4jfawsd5i3Qs8+lYYELKEefcb8QeSQEPy5c6
r6/RmSGQ8ljizW5uExGPcuSDJnQ8x3l61Yals1UOSXIibpiyAkpr0fiUWi2KsP4S
XljtV/XnB/oHVPS+INzdyxwyMO74Emx9rDjp7iCxG83PctFfzYzd0HnSyMYgHa90
h19VPMMwm2M5coLViS94ACbBCg7pX0JJRamzD7wJmAN+2C4Km29NBil9BWNKLcD8
xYp4W7OmwM3+fRCR1jXoVpo8kGkDWti3NpPTsXVEBHlMcSeFWst6oih85BzUrRXS
kLQP+75w4JWGTHVFmSdWGmgA5iAOKcPQ5em9EH36X1Os6/XtjF4xqjjIrVsIn/yV
SgIFQm/zlbuPWBNhenZFWGCriGsE7WvK5O61w0YbX2B5B95BkPOBJfNUaDFCasJc
B4QXMenMdeI3J5TtCZ4GLHw+vxAa5Woaw6uEEFD1Vr33dgxdtoF6H6+EEiWsYJvV
UPKrl3DEpNvenz6LJrIV5PQjEn3VR2Pfbzidv79JnumVGbcExhBoKzacpIiXRSGQ
ehNn56xux/IObX/nnJ+EZh5UrVcm1/eiyAQ2SFhEodqj/1h0vtBI9ke2iObNOuiM
tpwts6BSePBEIpxEhyJMP5Cvqs8rJb+6p6fzZQOqBwaP+ID9mjLiBNsC1Oc9z3Wy
b+msoo3M6ESzBH/M0qhyQ38eMF1disb/UaTAlZ7WhnAwckmFJSAwF5RnsMJ3kRCU
k4OOo0XwdM/utIwWIVJIuLwfkZnE6vmVlVLM6hM8G0EMniXFFrYVSwDCDED3z8oe
bOs0TYfznzJhm3DMud79O5PbHwtbuEgeypLT5Iv2b2nUPbrV0d0fHLvXfzA0qi9k
gW3VIlLR9UVIRc5ftG+hJNzjFdF2SwxoxCSt6lGqQvvqXQRX5Y5CWGD8ROJ3fJpb
KNwaNJms4PYD+8jAUPOa+c4m7WUwNP//kednmKMrNKsqLKhGcbgZ+g1ZZCKyngm7
mcUs13zxz1exIqWfQP1sesEtHQfBHATRyefk6+zCDb0pM9/QhAQRiY7cfasJSAPy
ybZO90RGOebjoGcaSWJgjGcNqDxyNYOY+VY3Y0m9VGJ+cFJUoKC3QP0IE8RVrUre
xsD1iJZTN5fAIuRFp0uqsQZWiXdBrGf8S5Wbyo11MfnRELGCFFjIAiO2lpSC8rec
Y8ibLvBD2+nC1etnbF1kXJOeMVWc+ZRBHcfwDa0VfQkQGFJ0gJNUpOrpw6M3DAKs
DbY6C839kABmj5vp7PYHt0U/nHRSD2kzoKR4ek4Nyw89akBNJwWmkgJ3HsveJ9wJ
blKqPDRytc011u2yJbBLnmW3oTIyUivsBqyxh4/KwMnD+SN3eZ3C+34+qxMiGvGj
VuPA9FLboMTK7Jjl9FVPfARQxi6WbFTZZaf7bDFonExprnBhs1F8aK3g9WeHrZDN
tXTiRgyEwuPOFne8wH120u50olK2iE+REormLxCnPbBBNWFbiXw0hwXqgr63/+Ti
PJH+F2B4YbhBlK2G3cBH3cGTSyMqGfUaYElm2uSiQkiL/7JCjBoxQQtopTeNf4t8
AXDz7wGKqkrpbDIXLh9zwjnOYdIa1Crj2ZNZUXduHka8uimnaNUwO7JzJPCZkjxa
yJC25jT4qEpCqSYoneYfrzOXZQj+x9rzDTNex8j24PqXmXUCz7UeMAkn31FgeZcV
+kspkoiKb4IHp7jnVAtQby9JcipF7rBKO+eYfyAid1RM+xbQ/cm8k6nR2GkBVr1C
fczvqCiNITYWi37tQGZ70KtIur6M45FOERW3P5fHrWSkVRzpHXZJqdokapFxO0/X
6NkznJ6CAf6e4a06fnxkpHNkaiLM+HNgk2HRukVHkNmoSxjxkcm5ff5BHn9Qnr6w
vcM8XIHDjeiEHvj9mpVKFwJKnENgrhVZRsKUWibZuUTUISaeeQxOwtKIcO2eM6fU
k6jyV2bPjTIG1VYf5p2l1orJYHX6GXf9xTdaAtd2wpWKS3gai48E2wxPgHm0CIDH
4j4qAvsaQR8EBKyev2HLyEVFBDMm3579AiFIER0OWRDyKANCJRYRyRS/N3ZRyQ7F
ukWMtrFDhAOnojEkQLp7YoqXSrsgnRY4Es+6BpCpVbyVYpGQchhGDPNWYNs78W/c
odyWbMEar/Q7w3BAuty8duNzYPL56vg+ljbCEpGgb0fPAoqzRtKfDrb/uxCvWr2k
eyiLF9XWDfF/dnr5YHv2eZYjIPJxC1Zr0R5iKgHNK4M3YH14VQnOCGPLS1ACNHxC
nykzjowiAThSLhX8EsEcP/vKUIUnPdbslQ6dsLeEev/G+2vNF+ovqseyhvoj8/ZD
UdjZS/Qwo/k37KNJPECTk+AurQYhKyNZE9wnOb/021Q4l/uu910lNFNJPMv1wtlN
ED8nNHBq5CT7kT1yED7TcBQPL726+4nU9cnciGzFd1OOwOYTMvakpNqp4VjsUaFv
ylVOhJJwnknqHm0eP0ZW5r5cN2ubdio16+NEjUrMTV4ZOmtahdXC7bjZ6SwCRCYN
khWK+1gL3sRtPXpkgk4NLfKVrOfti2rBM92tg1S9JAOLWSS3WEcyesr9KgMMP9ZE
ELkGdp+nIsQW/w4OoEGYUl80JVIbPhlBb/V0rpjrr9Iaj9x7ATILN9juyLEJJUXG
huYlurApX4FrhWJvZU0PBdVi61EFkuPbUYxcXns61UtyTmg7RXtywtKtZ9mYv00z
ot38oVu8yj8UcMgb25TLOx92R4sR6DahDVmaoEDR2dYPWy/ullnAesq4xskEB4bs
fwF3gTKinClywjNHQmK1ZsOxoDSs0EAVRkdQB4Du6JS8cVJQ9/M5/miplaJzDIWm
215L62thQp1VkFigXr3Pm0Q7/L3Q01yZwUyLw5VA7C5r6+sQ8SJX5JvlbM/nv9JY
eWXiemSN+7Tl7q3vJr75Yn5v7ri/rTWltc8FxZy6KeWlvdvdU7ogIJdp7LC3twhA
YjyL6MnVyquO/ehup3zbI5BmPBIY3VMTp0PoBp4mQYs7J3vUa2gaGhmE2YLZAEml
zNNXh2unDN7aovttne7Zr10c0zDngw8DU0LFvf4w7y1H06tIcT4e1tmHASt+xpQ+
nHf6sNrgLRidAqmysFDalk/nXKc5Ilox38U9jwTWf1icwfCdO0FaGFqtI86ZAcUH
hNv5rv81V0cbjoTg4Hdm4rhzQ98iL8F4E6Civ2yaeprnvBOSdwnI6m8mx0stEEUP
xedZn2L/gM77wZDJQEjKzzQQWDPUJer07hnJGaYJirYZJpaDAWTY4YmIQOGRyu/I
ZTnS7AgICrURh0KDPyeEAOUrHsRJnAXgm5+sBACvg8386QaaLOMJEMLultITTkOj
5rZFi6ViCdkpDgfXxhcj9qrRsO+MhYWyFewKJsxg1KMbhvPJbTLUlM8FjeiTvcJj
Whfmu8eJDV2NVbMuuq4TrQdNBrXQnV9F8+2pgzGMMlOXt0iX/c9/mJwMma8VN/jO
ugD5eifie7dXE5pwRMXUlrCBgyE6Zyy/is+wcgsCXvRwSL+36tY/5rbSv5HTx0a+
Nek5fGn3xDPelaBoF/Tdx3YlxFbkvf5RWM823huBx1n5BlOydwSdNf3niQ4lFQz5
QN8l/Gq57iVO9BKT3nqEfz3BQhr2mZyD3vmmHb6d4IsnpLwkkpejZfneW0saS0od
NLj+YpZeVtbqOamx3vmnUPVcpFhGzCaFVbvQXbo5dPKzZ+MtZo87wSU6r6KgzW6+
wUmj7/nqzWXw1Y682pVkk0NQ9k4BzhZLFvikYfSvm3UGXuL3yksJJTsaO1qVGjvD
flugv0tIhasiIHWIZ6lYTWFgCfjEX450osOys5bEE7XzICt8SL3JxNCVR2pemJMq
zhsEpI9m/JIWewQV7EoU4Kd+INg9oF00RJS1qgMrp2X3zQDwmwq1GyzbA7HIoOrn
+r9h9nChP3h5MGgBI8L4ekqHaskb+uWThUXxe4H83ELrBBjBQRgsp8ggtDF1C2HR
F1Aa2yCauvGYt+5YJskCmrF0MGBa8q/yazgmBoIkvyU5UReoczwIAvgXjm8T+HAk
SuwrNYt2Eilor7UrZtlBwUpDNQrWfwq9ioV2+gIcZ5Yz+ZuMINxY+oa930Hsz6P6
52m3ZYPoe8mT2Ieqt5RwPITgl97aegneiWwpTOVimdHVJHeXmEhvat7GXmEnic4G
t6otKRTSoBRDOFsxxQQBGGlAaHZv00p0n+HPas5gPM5skckmPf8zJ3brGs8X+F58
LW2zxYG2tzaLbdikksg3F/rU9mvl4p9st9n1RHlAtLHoK8u/PGbr5wghRmAFAejW
HwA7/dGP4mUTOTbcbkeeOaQknXRGYWYgdR1d53xePkPeqNOMvsPS3ygcEuE/z1Dg
v7jEhn5VH/jemwRtLOiZ54OdtLzJ0AGYRjggCat9VsaGNZ6kh6ujO609Q6XchtRB
43wXCWSTF1ZABdX1D+Q4V62HgB0Pakxv2h1cNK2l+pmDe1Noszf1L5MhOo5mvs+P
tyZMWGffNAvS3iReZ1XDZK5IwBIA818CJGWGkS3mRsjqcuZRTOfZ4DOHBC9Zdpf+
ReHwzi08hpzGoOfJAibcm4ny7jroCIITbR/0hgkQPIvHtSGp0wOfWjcPuw3v6YVn
mjuiK3CONIWNO2UXhAUaPekt0GqVy8mfdh7b2CIkANSyNczZbGh7gx0ln87D02xa
8+XNI1j556R2pdrqnwzeI8suXAi05kKjadEvRfT9ES7dyjmyCCi1hsTYhknzjNjy
4nuCS9sCdI9PlK2Zq2cWXXX0EFsYhoc5HhGtmN8GLGoqJEbydjI/iq082DpiHYGo
Xbv9BmqZJu870zpE5ANE3IH4L7vOsCR/TKc5/+VkFnLaz5Npjyd8ag6uGnjnrnYa
lhifTrf+xR9CXkpSSV3ll7sz9SeuPQieBeN5j+bP6yODvPwlWF67/kMxLplNpDOe
HU6sgzhFrKZ2i/Ueqf9TjGG0ncDCDWd3pyrMWAGBTGn0v7P3t7ODtlRi92MGw0T0
haf49F7DM9O5HPSIXKIzP9knSmiG6ot905v3dzsvJ7pvPutiZq3ZwKvkR4WcLAnm
nBxnw3cvT0BODYTTdTzxT3laf7pWYPMMYd74Xus++irOENSsrMZqAh8qJtQqMHrc
qS4t/8MK7LAAZXAAv56kdJrDhCyAZEF5NXX4Kmw3P5xzGmmFRP6KBAwa5i9B9HO7
M+YJGM1EKKXAs429t/dFEeF0OSBHc3qgGtOiZ4Sc/f1mZ0ACCPrC3urD9bnjs2Y0
l1kmo/xPSIAw512hOyey3cBJBmhi55XHx8BQt2+Iow8RyOoUkdckxSFRMva+24rG
q6Ld/Q9/JOLHXNjaTi+DZ0UpSO4kVfj4IUtE80x/yatcw8xejknV9k7Be9988wkD
vJUOLjqwgOHhTMIOREE13814RzVTBvtZ90X1ip+kPWA8dXr8/oKfm6b87DVK9Tl0
jLlicu91eEyl6J5RmaM+vC6UzMM2MQNsB8SdAOXtmkFqYtssaUG0XedW4toFNa78
0KY5OKv6kq6EUl+lwVXgtQZ8IK7YiThJBIV//3zi9gjfOG10jCHsIAKnK+YCow3I
h4ZaAPDYRV6I4ZWY5abr48O9YBwPcedK0DBvQNzXyETTroTwztB7AZbbjguwSBHi
tyFQQMce19Bh0Ln0nl2xD0sMmX/udAHq+DT6vtneg5wHwzEhMBGC5WDL4xxu6mW9
Zlljhc5DV79XB0YWCf9AlzCN3XvWP1B4Mp6wFh96SFUmRD9Ezb+bqIQ2hBBTd0Uu
cVr3nblnFRSs6I/Ba5Gi962vU/1oOQJ0kTCci2sF9Aq/VtUUvAZo250vua6EAIJF
WLRdi/XAQY0hxn3JWXEB8e6o6/5x2wM0Yb8mtjqWbsBqALNaAeBhhEicTPCAA796
a9tkJ6emfsxVXEZUW2D/pYvJuZH4NpqD1VxDW67os9/x96VSA4htd5+aWADrHAM1
b/xhBu2sbHjzfrIbQot+BWYx1cKN7XMUWtvH2SSDvbB/y0Sy1thAzg9YipvIX+YF
B2jeOPO4a9JwOUh+Lmc6YZVpQjs+1zQLfhHVo9LEPQJbp26IP8p32pX6d771XzR7
jLqqbera3BssCyjkEXDvZA6YlyCHd1LDjUmPhhYCyOqHHqWgRSrE6UL24tEMM0MD
u42BQybwj2K4PgLkRv4JfO7aQvPpH8PKbm151A5CKNMoRdhWxpL4JVUEtIn8PUMi
Z2dmkOgD1RE8IMb1T9oFT3+tlLmmTcPacteTDP98sFj4yEHM+WFrbfiDu/pciXS0
BiDczh1A38iACeinKxf8sqZksXEQxwKKPUALOKi/05KSh4xzePfKla1bR/ml1+c1
WtCJ3uvq75fEbJiSRxfYIZCs2IGbIVVuMJweFU9vg3as5tHjY7xJBrvG9VoIrFOY
GdIEIf6RRjR1T8zR/nn7X4sCrVJuHFavfsxCYilZUdeaTcL27tGE0YcNxrZrZvGA
YKWGlcTi3aaJpgu+z2THDcVgSi8EMmC4K2zah5fp17I6khvWI141NxJLGjnad0Uc
Op2iovyHjKHGihFlcAXXE3kUZ2xYLkaQgscT+hd8/7cZUOLisjFcg1Rtze7bH0ad
64ZAElezF0PfMdD53/GUpVFzqFzNOQmipvB1ZB8BN/95iWPC2PVgEIbIEHAYJFic
tpt6SsZX8AnrCSGGAS0JRJZnTYH1gjKp5JG022/no3WWUn2E0rBaGS+VRv9gevwO
0O44/3p0gWrIfkG+1Ub6oIs4F4TX3NKwRWnwbkmKxjtAaaMNZ86uc8wkBQRxZ5WR
jpteyD3CR4GyGUAQejYhy0vzVemp7I7+/f7tPAEXD9994xozaCwTSz3G323hJc9B
KVub/yWxy54NQe47f3dqGAOGP9W5zVPEHsifVraY+BoFQCJ5+eed9XSP+wrWKgta
aTJdsEsW55LPvJL3Sw+HykrTMIMSlZvGdbAeJl7B5U4rgbpREoFQfyVwvfi6LW8u
imu8ADDFdi8HLFbNfIbLH7+vr+8wbMamHXfQ/luqZrTDw86bifWVupBDY2Vi+1j6
B8GAc3QZwDfL8bdUWLwIWGEtcqFHoGtfBB9CjCVUoHYKsK56OZc+QvaZih4MXt/M
qOxbS9u0Dj2QodVy6pUDZMIXi9cwOiJxYcOhPAcu7T37VVnUrUHvXItiY75lC45Z
f8tdideIqYsb0GUFYvfPIEhPoAusdHr4yWbcdsKwJ5dikrUxIWc7khMAFAFngk86
zQyC9aUmu392D731l8RmQD9q6JIfZRtwYXm5WDyOjCQfTYbUeP/7ZEAYLJSOPNCd
TDTm83KUzrcPQVy2KBzFgi0JfQiz9yhXE56WkNn0MN8JfeOrU/69qYlSaE9WVj68
XEpeANnzhN+YWX09VJDQhgIGJhTHbu+XxMiRsTZlqs/ZoZ2I+VeWEnrpYBY5JZak
VZqR+fd7CkTWurTSnBze4bLscj1FbHOHwap1DMQRW6cSDMpAG6lrtIj7YSbB4IeY
x7wBs8Y+23V3DhJAQJdEBm2wQxn24SIBPFqP9ca8ZPycqxKUSv4l965BAN9XaBMU
8/Sm29ZzMg1MuvsacYYvvJK/RlbqHVbKIl4XH4OFcD36Xv88MlRiF3hACLjk9c7s
t45SpNnOw4EGsCzlfuJIaCb5vOB/C7cnImxdtRoxv1XAAiLphNNrOzMzIjCT5tkj
IxUUrIr4rwtvg+8RFErhOYDZb0uEuPToWL8n2ZPxE0d4samIaU/UcV9fWzx4WLkC
zo5/BGkALOscWBCzHDQdvIhEmw9DlavtDS3ItpHCqzwFzV1FJr7su18if9BoU31X
vNhHY0KR8aAME9w5YS2js4tbxVfIUFBnLJMhmoOPPmUg6WWHhdTWJUONpVIZOuDZ
26IshlP/b7wxePDuZqemA6nDMQ2z28cKq6DxGce4RwAjwk6GBr0Hy8ZLKSOiokMX
vJnD4zejxTv37WACCwgr+g7rw56cqb2Kvs+VX4iClhC13qy1PEFxwK0DhEK/RfSE
FucP1RX/u5SLgq3tQrg4o3T5dU7d6911Cb+qtTqXq/vSKpfvTckRFaXCKKYEdkTE
mBedO03BbYrVEQv9HXMhbGMsmARaqok5KnfHDhXJ+hr6O+guer/VHwKQHlUe87VT
aI5rs3ryBSZb3oH1MIli/dYrYSwnFvQlwCEE0EczbNjCm/hrhFRk2P2ARi/TSUBl
rWzu4Cf1n6K8++SBp3eKRD+3/ObZHEWXtD1mlw1/dhkqe4SXu+Ja1pmlVTJNDUyw
P0aOjWXQbpusyiYhmH6ZUejh1rcX4qzdwQiz0aoos9l4Nr36Y63MvCY+HcvfbHRY
2XDkfcaDJELs/QntM7s9mDgpKfiKyLvlbNB1kY7WqNv3HNVHYmvWmjfZVgRQi0+R
AxZBTk5Hw8tQiVlQE1XWnx5Hy2aTFDq3lUjZi/vnL/BxMsmjytRD9fy98xKW+sIe
73gP/7Cx5S6oW3KRqZizjU8/48+HFjM9PDtvA7EgXpMWbUyO6JcIYiqQsDjmzHjH
cwZBJ3fXKv1sh45ndS6Hcm65c22Ey4XSjrrf9zSXvaSUbHBwFAQaz4ChpJDnt+xt
uqI9jWHwnuSLRze3hZWkx7vE4p21qPp/Fwwzu5JyoruGx7rcqNvtu7A4xXMIuHYF
hXDh5MICyR4ddWOi2Y/ecHNe6mFwwW88Fey+e/DRZM/zAft2W3zLMdsnkcXQo6Oc
vmUEYMugCA6F9AXRCEIH+yW9N15P1kOuC6R6FXvHUTE3Jjb3CUKo8TjWDQMoOGV4
nDnVBCdvQN6XD/uKilDEm49WHwkwX1rpscnj62LgftmAl5VTtR+MPhHlzrIuU+qo
wyKmwohJn5VoI965XI6wZrKexuIXXODtQpl5DgbUnJ6JzZB3wq+BdzFEXQAC/2KY
K77ZNfP/57tQOAa71OqLJ1762p7fxHXInsGlMzMXn5zvUS4IZRmpKtmC9RtPEVxa
yYhHovxyi7CUp9R4yB9Iy5M4jRIAcUXz6B+mfO9ZuQNyosgA7SAvElsA9Uf9JaHt
Q3H5UREKbFuQYfTYm+bTa/4JI9EoBjiGc/uB9cYw1fgNJDIcDOp+20LGdKUiS/QC
DQWkAaYfHUnmvRPdSC2fTzGYHF/z4WnP/FoQaACDRkHWfRk1pas3WbMmKCF3Fh+y
mKDNbrJhPCt03aZC5JNB87nvXyDdn6luYwCJ4yq71mut6wE1B4pvHMSss/PfYVoc
nG1JRiAAbgNa48W9iFP3UDWoC3A343UXs0kGcpNpRDEspYFW76X7NWuBelj701Ql
+ebuL35Xxrqn1xKRZdUgJLKkwmLwI1gn8NzRHrxgV2yjhSvG6eF9LvzsUuTGhdUh
JurPoEXFpv9KamS8z1flwe3ruPovgAFLRN3PBdy6tKDgE3vvf3gUrPWP+J7+mPGQ
P9tRvFHymfQjuup1tu2qZtZwwlgA1vGVnqi5bfNq5i5fsiRq1TGHreg6T67mk28S
LA/gXpjTH8u+ifxDYC4Ly8747kFiXt4IkKS75m464f6oBwp/A6jkz3U3hDOC7NRn
HWwYtlHo7XxDrPYD8Kqt9AnXhF0TSL08tA7wlfI0VeQ2hqaizhxkqyOpvAMGFk89
8lbm6HTK7KTmoiEh1PLoySS3giDxYiubRwUjoM8I6Kim6m0x7Y38/qHe60DdK0xq
eIttw8lp9NjbG5lgYmPwgICiWif77gYrCaWTRp6dq6UZHoCmJFUTcfiS0UoQAxMI
UbHhJj53/xyUzWIAGYmevdd9wIxwAmfHgZNxMNmJ/ZjH/xtsBOli+VGtHB9R0GP6
7ZJpirOO12H87fq6702mrfzdpRliwLu+ATbxDVar78GLJOmlyz+6cHlbWMHwS0oB
EFG72wC1I710ZwxjhEWR8xm1kPx8KLlvw236a3OBC2KTIKbu4uFkX8avvddpMDYy
Hq2ET7E4ltcn0siMCusYT1us+nhqsM3+sLre7CKtlXWH13MBk5InX6RWVQyCOZfw
5AkJ73FQI1ne+3s1tsRjznaZggxjW4ru6eWayD+a4hxjTytNYccdVUVV0dv76H+M
lzHq+yNVga2OrDeJv68TVzgoPESVS6WrmRopwd/k1tEvNMYfInrLqTQ/oOdiaEkA
uhuHiZvLNdrGMbGBTYAYXe+mIuznPJ6ZH1I0FVYS9r76CVDKnQSF/ma4demwpMXa
yQykQUZEKMtvO5LS1JuGZkTifZq3lhmrZnak0WoeHP8AnNVS3BY9OVkfcsWjgQFq
bcjFgH9nPbX6RPZjWlC2ibEULwHpmIUaN2qLTqgosS5eTqm/IJ+KwpWlJ88TkTPU
FVAZZ5IsO+Ye6lhSjEcT7QgxW/CBjfzzVtD8qIKtXED3aotlTbKF8v/Pt4hH3SH1
8JJ3V3fVRTpGhZVApqBdU14hp+X+PLN3YFiIrDk2Hnu6Sbr4Yy215wFEsTOAF+8E
JKjkNHtNj55bzc+UpoPA4bjnkdvH4Q/8j5UO4clUl3g5ijip8cL+ssYF4S7ntist
D1JbXCaRpIV4ZZ0QGPPMIwytLQXZ/WL+OJHOx6miznGeKHnE530NpV2uYNAgMlw2
XCFGiamBzoSJ0Ar2h7P6fIXlAIglwDennxKo2BJyFvBdZ6yxk26PGJ+eVrXYW5eE
nR0XHJG8RsWpsEkfJs2xWO2QeLZryULJB8vPKMWcrVgS/qAkPduwKBNEmLv2JSuc
kvmKhJTf3FecNCRuuVKIIaj/o3Zqx+LN4EBmo/PPDtJ4Fts5LSKqTWhVnU05DauV
VJ9Yp3cw6iebwoPGcctSDE+l9Fj5ssI8/ex88+a4w+A89l6mBS2SSy9u2Shd93EQ
Us7nM8RhtjkwONqQPf4nLxMXLqM0/n/LZ22/k6+Sks+yBWhT9fbthuVGf06+9sXp
RKS8GYm5Cm3yTqM3qi0Nn7hZns/EjbQIGAG9mOuyRr2zg7+wECd/T7ym4o7l3h6B
4r/8xx7touDnULNC3Ad9Z7tUg3gzXFqsrDeHa9Ru3rbzvS9KC3wcXDimSs2IFA69
2f/utj+5OaTI0vacZesbWvwAqjM6GlX29knQ9aRmtVQ/VItVenr5AFEMgcUJBcDU
hM6Sb0mHQfxqrHsGgPj2keiNNYHuqMFJkqwfNUAzj9MxXEwa4I4PGB8wcepIsOU3
IiySj6pxk/IaEPZJv1IFWnhi8EB7brkZ2osoVCjBQTXARH1W42+qD6+PWFDtNZ4H
w6KHBhScNOuo9SlEr9n365toXtfcARE+Q71swd+jgrjfBejc9PIOUmy4gmhsyLJe
ffeIrPT+5ftWiWMV5YNAGGvyYcufH8StPtqaHyB6j91M24QuDMXe9bAavoZ/gYjK
E90JwJ6Pr5o+T5lT2ye7+P+mtj8q5v6x74VMSJnU+/IPDRNfdmj80P6nY7ReFcfN
6jRcIJ7EiOg9BPHYnAMIQ9daIk6wxOX2UMQ8JDFGesKOj8zN5EZ3iYxf8LZVrtt5
w1VOveom32AxPLeLOanBrxtKELllpRTLpz999aCsYtA6+7xgBSvCPdkg7CrgfuSd
CNO74YJO41/NwTjbCdkHiSGX9eL7aFphcZ6CHjhd6pUqqAm8IxMCw45woA3nSp20
T816a5xXfz82eiFAvMBUWY+wdl6tFM6HfGOt6KWRDdK1E5PeU9kX7syZt9pt8stu
sR5kGnW5aiRBFfLumUEDNv/3SzsEfSfTVBQDftmfhQPVHkb+DPO7fUJR8BF9ZeaG
YYGdqEpucI8jH9SZyAtQ/RYYqjrIqlld/eQuuVudA/aPpNsJwRKFYVfl/DcKpMjf
yFbmW+CuWY3q+0qJQquiMjcFPwD9r3isbpBhGwckmMWBOAqVcAzs+F8VWag5r9i7
QIj0Vlg/QjyldhiGVmrV58++ZYKLCphbsxrKv6IxAGRmz4J8hEhZtcKG+/A+3Fba
h03ipHVRx29yPxal0nAT3pbDLPtiJsKYm8kSb5GARp8J9e+/FDa3XqzmgWurnpT9
QQ7fkiz4bJTtntI8KqfTvVgcHXpBay04Hpc9xWBMg2mkKxgO/TWGJVU0jU6dixsV
VgF1R14uiigg/8QwBBjTnncIGgOwNSYDrk7nMSSWSgRDNsteFgX3ZZTXwiOcT+h3
XTTu6ZEB/7sMXRAjI5FwxKieGeMgyJ46BHojNjU0NaMGra3047yDGXC7Q8y0/SgX
kBQzAHQaARmTg0nUdRpAHEMeH5C/EqWcM2y39q90Lwdre8tg+/JMvaC7OYUQuqmZ
em3Jeq+hqWQiE/2Z+OPJKwKlwmJe4YlmYkhga3lsPepACzw02z7H9/vHs9eceSrc
1XhAzNo7mExzYZikYJEoXXugC+2T94HQubjE6dI94dkW3P9IhCUPbnMZ3Bf8oR2M
xJkMYb27/7lyfp3eMk6BOFkb5eAqMcoTLFcLPQuR2a721FXYKI+z93AAUO1SaJ6A
zaO6edaP4LCk9YbCZGmQn4V9zB0IGeWyzyYIbTdAV4zoiB1M+0p6S43M2DWHpzv4
ynQrmi2MtXCpF8vTbS13DUSkl4bFIHAd79qTeQ7jbklP6PQGuPhtYxaR2MLBNiJ8
zc+6gIcLYZCYekZsOa8wJscIae4qK8P1yIwx5U1780m0dJtSIptlVzaD3dc2HHhA
I0CfieXVl129Q2shVOY287cL/uuhkle1ymhqrQ6GbpHN4e0GeDi6sE9fiLrZ47Fn
ilTvwBmnO1uj+ou+Mj5sgeLH2OuGzpjqjXxHPPL4aKz6XBt1N+X6jRwVsjmq3PLJ
HSzaB4MpXmn1A4P0inDkq+oEaFNlLEfuDr15ILPEQc/1hsWEQGwPrkt3fWXhM0H5
qOD/v7A5YkUTVT5mQMG8pviT4LLTNvFcgwNzmkHKzzXkk4OR7z7qFb0SvUo90AjO
06iHTbpoYPFkjQxvLdiBMHQOU2C1nhYymPRgnORlIZhbmstWdnoRSsTTJI0TtDP/
B3NTcol5W3EvFbJyglR38rcQGxWm9VJX4/qHMNif/njAx4wDEnHKpdqzDEEAnT2F
TpePx/zuILhAT0bRmtbk74OM6xX8gjTVB8AG2oyAH8moL/JvIafGibtzH4uSL54c
B/gMWG3nfvZWCrPYI7oaFWKE/79ULCZ1+gbXdr7Hz19J4HAnpMGd19y7hC4anBgA
b5wW6GWsRagshX0PAiBCvy7G2zUCyhnOLf0lzlghjzO8hpZ9kNEWAqLPEsztRtE3
wfVi0FP/c2vjFfR3ILWmpE5cgrPvYUjweYAr/cjGSDgs74EJHeClQ2m7peRX46ZC
Lh9+aDe7cSYciJTaMR1lSPDwlz+rxc/JCCQn3mlihPIknIcHsfbDvbP+05YAVJ8J
zQHQPBsf8JFt14XFDMPHEBGtkut/ZiUUACdo92SFsdB7JEeciqrJzK5HN+Fbc71M
tS7FazQ4ujMf/mHhwjkz2ICbmTy8iurQVI0BMbr8q+t6svaycB7ieDBdR6Cy10fW
4UbfnlCMtpl6vm67WRQeRewIuI3OJ2xu7ur9VZcbTN9XXv7NP+ZUyqdrwDI23YMu
Y5f/tw0q2yYgojomSuBrVu80TB44YMd8KnkO1s0CUV5ayn8UvblkuFjLdgBxMa3G
fY5QNrkj9BCvbNZhk6IEuCwVYZT+G+ZzOmPmcPLwgI+SiL+QybPecZysf2DvKsCK
f034IrhvnKEEawrsuUNAqVoYMWwFYl5mb8kf2uECPwHfYOzMS5+cmP2Vqz3sVKrk
Ve+CABMOQnvD5wdFxkrKGy6jVp/5SVLV8Xsp5RpwD6pdfgJLwwwmFSOXrBbFGwoi
Xr4aObc0j/cygrPd7WUxOThgDqKBglI3lN3WFwIuFLfskn6bjZoOqeLxYOzgBFV6
KcYKblgX3XrfG2BpltNBTye83p7vgWqXomMGb5Xwk3otgL52HaVZm1IRSSsqtwhh
J+XjLjD5+oftbZwPakWC5nJShmQ0ViMgVnl5adQ8ZptPGVeHTEGp2WkAVKcn+wUF
mlmPm4UU7jfXL+/zpifyLJSAOW8l7Czh3caSun8s78Al+tgjqIBv62ePSR63FCAU
Rz3+5P2yxayGOEDN8yWVgsi/fE105vsMVSfz4/+Xk/EVuNlQWJyH4C7EVFhBZ9O+
DjOc6A1mvOqQ6jjdWPnmzR6+jdNgOKqego/p31OG0tOwgDwin+ACx3nQDoMkADIk
4gf5lccDL4L1ve8ix+8M5yu3YOwBEDBN3XK1z8uarzm9ipOLVUUUwXeGjCWqAwrA
IenB7Vhn7BXdwInKvN0UOkoMu4oK1sW8kQG/prjy9i96x5lZnM51Ww4K522KPdI1
EnASUOV/divmcRpDVte63SPUTLEN2y82uYNe360cs7Q2kldEbA+DnjBXYtyncvvK
OKmJ4nCakpvCxCbG//f/7RTymThdWpU+46iRM5SBPVmiSvmfY3NEgNUJnD3STboZ
gCclS82TaedzaISszzzc/aLncrOiqaciKmzQDQ8cmTovwk0zvKSdMgc6fooi35+g
2xDeR7S7fnSd6kKz72HmNFoCAvzXRGlWbu+7p9V7InL0l0240g8+DfvY/fBPmubG
iuBuqz1Z/Dh+xEVGKfKwT6DeYddLAQQYO5XkkAekX9NAK+f5BBjb2XQZPGozVBFW
vduWzn63MYwrYgtgzhlvdj7Tv+opFMuFtNWZ3HWpwNMcU/AE/+PYazfN7HLtMg5Z
KhCvPZhTDdTHt9A6WunhejSjCyMmCeDMzes3H6XNQeUvd6hjgQ1Sdyjv2EBof6ZJ
jVtGl1rD83XMf23FN+OTnMUOn8F/nY/COv2Bg+HwKpQwXr1ZcT1agX2Fpsx01ooD
X1ZUrb8wc3orXzn/m4xCePCyTc5nB6TVvIgrMGqZWXtAShGMEt/UHwd0cje83iTI
iUpL6eApTlfyv9g/waR+7M2afvzlwzIa6kbwJJ8rv1ccGeyZ9ASzkbIqIViebzVO
tTxLY3d8+QVylPmv5Qx5Moo5F2B3vQMy+fSDJQKxWPT8lOU9CkH9W9hW83fzqhUh
RHdHzucda/JTm/s98ih9t0m1qwqmSKqO2AutT10LldsiWIRS1M2uDXQBkgBOKMG4
y/3nfVjA++hWqDBI48GQNvfWxfgdpqE1NspUw3XvhOJP5o/H36ZiykpH5IGWnSlh
Csvh4nuN7zcsRCx7f80zB7xFHkjttF3fk/TKl/V2YPahkx4D88ncxtW7MXdT1EVQ
qPlK2ZheTdwYDKR9npqvIEsAKPZhMmyWgpMqNjyIKU9oJrA7759ysvlScihQmhhX
k17Y2AfF9fmEmEuxNLYwi4ss4/fzSaW1ZCrVCCNQG1EPgT679yzsL35Un1JTcwSu
k/fB8JDymRhopfXI4FyjrorjCIwdb0nbizY57Fj6ku8jpKF0CaYeGnIwmf7737W4
EDyNxuLcE2NYfIxLbspdOU+zhQuNiNGYU+lXkkrit+gFscRO1xQAD5T5Pp0N2D+q
6vC8lceuZEo8nCQaTRIY+DvUN3VgQqgQswMNtWM2dodKncYGWuwKKKyUdfU/kp6J
s1D1FYaC2rgO9yU8q/bHO4EogeveBnAvv6etTiqzanW3GwVba02EEAj7qg2Vzu4x
9ScsZmfivh6ri8cn1VCaUAmL87HTx4ctQYEL1+h6w639FfzWs3cFHrruRpRRyYjL
7D/PDrg+Q9H4VJap2SEbGyWE7lE8T4hoM2L+rOpFd2QuMR7xyK9aILxg9WgJlUi6
ygWmdTGs20KMCMXBMtkslrqKOKqQn9olJLzcVZ3i7W/yiX9C0Umosqyq7T7ckZy4
aXyv6e0iiczw9vqTftdFrGrEo8HUrH4zBD2MO33pdv4ViyBBlOpWqZSH/+4zf8OB
+et+znv78KhmgDxurrSx2lbEyhnXAIJ77X+ZeNe0ELAPmOQLWnVPCA2dUAwjSfzO
yD7srhR7a41LOu14324PL4PgNo7inDyY6MhF5dlmm284/mqqQm5OjDPBVDOO1WtQ
YwrdRwuS2RBcgCtP0ohb92YXJVKRBvrT+g5qMapSh5kuIIB5rkclzDdKZ4A7Z8a3
N9NFu72tyL1quGRqvMc4dhx2jGiHInL4PI9BymGDnzeBp5GEkZNwW3Yb7igbtg4A
kkZiuwyBMehxZZRVPKAoD3TKENbU9a0LLesEKFVjzr0KOXubYvkLrMjwXsvJkz1p
NI5BIIShphgms1ZJG6yLyWQ2cC5dD1gLEIVQWEPDHqhOUd4MudV6jALLRVG2dRkZ
XgzBZmfC/rHvB746dhDWjTxVuLOGhyAKcVg/ZzWm/UuAGK80zKtIACCOWFi/dgys
7x7lLe9qsEoCeTTr+7h/QJIHds+PooTgtWFX+JQZ8pkmSdt+1Rh5FttPZ8WUeQr2
7E6hXVOwYPifD7MZy41dY8Pdddk43ObVGA+jt7wSZdOAI5AdSISUZfEvPoBRdMhC
b/BDi5c5nlnssiLgR/2GhNEp1mgZXJ2j90jdt8NZRUXOfSoCYjWCqDVZ1OxnIvFF
PhM5YQ0LQXWx16fINUm2yRTfshOGRvvZgoepbVe3ZWzwD3GWI8v9tRPWYsGndsfS
kHLWyD45Z5PirgVShfqjDL6cdNqGWhZmKy25Rmwo7BUn+whRR14L4vFwAbKcPlu9
Rhyt7XbgyEEkH8AMEo9M84bebEuMgMymXMHlVnR0GQTKY2jNdDuvLIJZHRNIC5HJ
ZJxfmDaKdz0zAa4Lj4zwTzIj1ay4l5kdrhRZRT5u9BK3+3Hcm7vG07rXS0BThXY7
f03WlcRS69QMoB+EMI2SKOLQ+fiwyyh76dwJg9kfr9+7hJCWvTmbqUn1U1egJYdY
259mi2h+O1sWF541gRDG21xjTl4UIvuyjFKVq4nBDJ3jUr0Cpxow2nwDvNKuMyh6
sAwzOPOE1REnxzWD6Db3j3Ea2A+m8x4LcZ/kWhgIMlhOXrl3JAz5dRvmFTD/u4ec
VPos0s40oQTZ44lleSyibmBe7/hsNVoz0rC7dwqsJNHeWiSsVgih8fQnXX+tOj9y
3UBl7dpgw/ztI0iPFfo+4kANB11g4V73CWW34TEAiI4hToPb+tiDIcWATpvdLtGG
L8bPHu/BfY/SRThsOj9AXJltJShpWHBarhNBHgBt/qM873R9D77rtjAyuc9A2YIE
dvaL1MOMYrm1ZsHS9QrO9TgsPMt7gv63xJge8IX6CiIyNKtJgWD5MT1Py50/s5G/
UuWmlcT1pwj26TLeGFLPeIMBCfH7kUPqFG3L0pX6y4WDgA0Ko7LuYMraiyBVSIap
58clDMNBpgYJwYXuDxy2Rvi2tjkGBUzKH6E8iP4qtkepgU/I1JOvK4lRH7KCY3zT
lqlNHEB5wy6IAo1jdnuTiAhskxFhWZIXs5whQl/EV/qxLpz0YRDrBWCbvS/vmi+X
gv3z5nQVe068YJB8dPdisxt3pyi9Dq6ikXPv1t1QT2WKFONrjeoL/ewSxOxIrliI
UH4we1ZZLDnZPDc0egaKrPx00r2ffy/X67JgFyGjThBWCfI1C3hDAjAZ01zRqpRb
c0tyiiKTzliu7/B/PW0SQYeDgfbrAHGVxe5f51OYBVNHQ4JF/bVXmoc/e29jRF6l
PNXphQbj91T4FMj46bm1RjUbp7EnWKsm5XpXtysP1YZWi3F1X501SmQG/KyLfW4R
MQbbeq7KjTbdXvqXkAMRg/DJmwtKxEbjIr2700kQ1zd5N4fqzJMujqyH1V9Tn7ZH
p0A2+rytJiSEoux3byHsPLJf2AImw5N92vxFpu0g8ZPYqkwqWTMV0uM7lVglaJeo
3oa3gDMozco/vun6yBUumtCA7REzFy/ZnVG37DR8gh4CpF5Umochz595jQ7RcdU1
4JDDdXKIRavrR79/I3BlJfCd/MLy1KCv8hHBnx/0os0U9T1ktxulTwXLi2CsGWvy
AoNz8Pm8PM2ozP8EF/ipxApBtinW5Vz1uwiuk6EbvntosuuH84R8nkNdoNVsz5w7
e29Z+NHLnp+Lh3d/mHlmAw99/Xr8PIkK7NimHd8clVBpJlOrr7nG4cnbNdDlaidD
x1r7c9JN/NAb/GGqAO25dMTMGXwl5UjzMKR9oech/mPapVq4N1XZ30wKvZlwW9lS
okmShtQcwuoGcFKpEyX/3VqbcFKt3bVerobbdEDUFToEoBnlQqXlQQ62UuUU8CqQ
eoS+Yzz+q91F8s72Oiq9gnrOhD6vM8MEv1nTSuRLxGrRXVKdcACjHWNGkbVvjgmH
QQ1LPg0C3bmzMuJagy7F+H6vZ1ChVf1RZvNixDwXdGTkyQKTnkWA1XeoSd5LKz2e
Yh0oByRwIwOnybfxvQ7cJqMDXni9OD2DVZXLuJBXeUcQrAGWwZgJh1+MriygX2tL
iwQ79gXqECQ27MBZujdHdqw50WRNk/4TWgdylNK5iimqFjWdhdUL9UB+yPKTyEGC
x+UEXaEpiLGD5GdrRI5wpbYp4uIqADONxxbRWNze3TMBZ9z2SZflI5Rp0W2x5f7+
dE/qVH343Qh4xmg14nfBPodYVX6MyPAQkodj9BklrJ+gGzIKWudzxC+OoyTShvYD
RfuhRwv1gxPyvOnlqlXkYaxwO+1C5InK33yLWA5KCebQ/vUSJo3vgqvFJu+Eg6GZ
+KWaZKEzhVSHZ4JY/DIUwlof4gdFRgbzz/KZu+OUjBUHQZ33e8pcpnV7DMxhCMnV
2IyKO5ev+5G5omYBTwN6zTKwI+LmIPz8gK3Eu2Xwv+OjitV9+MRb461f7dGriYXN
h31L5OrcGLEbKFjx1ALFtUbj3tBYTMItKd8UAa8V7eSBpjdI9FCNsAiZn7iKemrP
GNT2Yh4oVDJ22Eew6jSrStYjbwR4mvhQdyHfxhcJVEcSeWHdSAmO0/DYpFro/qRQ
EI30qkF/uMpNLRlE6N4tRPbMH8VqEjVut6IFDKpKkZRScUijw2ThiW+YSyQanwEz
UkYhMcYoc2NrlAmWs0lXsKl5eTeDRzBnzdaGywNvQ1kMvfY7NB4bfa6mfmKF8HXF
okazaLiAUAdCbjc8TTSPIcwdhanX4fzVvUmZ8qTBpqpqXWS1yQ0Kj1nVNTMnjWPV
oFBMPAlJQgdUqV2Fjf7shpY0CCHvJ4e8EqLYWvqTpo+THmXNpude5RvuSOFNEqco
KSzFDNaMnINf9U1NCEuR/19mRm9Iy51ZeaWrftv6613Tu+sjYzHCH6vucJq6PRBE
pEnI/6V0l0BsV+UzULWLOUYMXZdbdTWgJZXFC8FrS9l7x4d4iFHzf357jEwdsVmX
ftuZ386cX+g39a3BS2aVH4tCzNCZfo1zX5wPFPW/KXLVv+LbEx1epaqS02SMK86Y
P6qwRwXsCHqal4LO2+EBeOVIeGmAWNIAKAquuOEzPS2eFaNQKOZewAHGxkENMeSd
lOu/4e/pho8NIRXIe2TxaG1+UK/195APOdCLLsAelUz7tX2koV3PJjgGAHWIht4x
pbg2ytgM9+xw2dcnWHD/aDDp1GYnym9Mken9rDueolMJZdNozZMTGF4X6eiN4nJv
JMY1Op+my8SltF/N6Fe0u/yzMNRu+C5Tw0fhDHuIjyiPSHM/oXvn2/zG7xMKnYTz
EnutbmP2T0DN6b+LuPdsNgMxX8r5A0BvpvByLJ9Sn1NYH7Bd7bYwsZ0FLngd4Xpc
8ldoFst11XZOPYpPLcIrSp4wVcM/bhLTSLYbHCe+Ro17cr1QNMnVj/IaLLO75AQl
vALflw2KgLD+90cvm+75tW+ydawpJe9cQcujbKgKuahgVgF700jWJsqewbA037pe
rPniuGbRH+3mpf6U3yaVbxZHR7lbB3H9MjIf0/eg+o2D0xTXE+06MAYlXxvevhdI
LHENFCJpLnfTkm5PkR799gmP8Pt6i3S8hsrukYV5K5AEmeMPSwAxvTyagoEDQJnl
riVuYjznyex1G4XVnqg1MiFJ2+EteLkx6AwbExcOPWT4BQP4ASKJv+iU4IzWoLko
Z7Kp8spDFglUqze+X6wmvygqYbN8WyWfs8yaAapf1wNf9ydI6QVx0p26qP/nsEiu
qCC6ELSVm83IHlbXZqJUDqnR+z/tO3tiOFBtKjKOJgn85EMUlwHR2BbcHSjQBDxv
tC0ipo4tBB73n3RwVSWJCzvqiVeKqyoPcIpDlrq+XHguDD7xJShEfk1VGVLGOgWC
uslAZus0FTxWF1QoGYSPEJgAOGBY8PeD9hS32mLC6EZeNBOllinr8+qLDKQZKARQ
E70/ca3826FxUT/T84pI7BBYNDvrgjI2syc/uPDLkR2rhIbUYZed3ktYmGFRDeb+
rStis2/NMLXS0h57lPTHZlZonIx8vN+z2szjxmhY1tlUF2jGuoZxeBPIac0FfWou
cBD5SR0pKNLMWSOtjnIf8vukr34h3xrpLYaN55wUsWdplEWbacqDR7fbOaoyajox
YinAsKy5doX0dEnALxorDwF7602V4rf3Q1iux8hNQBja0CMC5oV3yPNcHEdvHvbf
PLZA51oOkNjysjvxdzSrYnwsaAaYuRxviBhPNw414vUlZTbjmGymD/5sF0OwaENL
s71d2+tLvVn5MlJeP2UtY0TKeFjX4/4aJTFLi/dEM8wVTrZEz2UOtCZXILgjAipx
ZkvvAH2Aa1tPFneMLs3BTqi5s+iY8O5LfEzugfSGE9w7m1AZ78m8Ir5qPmyrJPal
QNIkom6BS8/+o7hE9nHf2LCMjk75koCVWL04QTG6ZJTO29dighexva0sZGs1M+pl
Nl28Z9L+kb4k34ujc03zG0lmWzz37QJwDuE6YkvTIYKuV8BXYaxMTdNXhBqXf+Sj
J+wldW/YrOVW9owtxGH2V2e2GstJv79fHxoA6U3plj16KJV/FzgRJivsmRjS/WGa
/gkhxtVFvg+R2lkbymyzRULFzPN4zDW4QLuSatTC54l98SdfBBqx8vrPJJP0Nr6u
pRpu13WAuiODEBhcyHeoVmjQgtrkOLlkH8XD+eLK62jbSgK3Eh1rgvUzqr6RXOib
BfkG6saIVhPGQXcB8R8NxhdA5PZ46Kqm6mZAhxU2uemVG5Z8xDnD/OVUIT9J4tD9
o6ZYoeN5CJbKRsYzH2+yJ/lEEkWSfWdVVL9PKgKBMlnkQUuSDh2Mp0RnqalUfPtG
KhoFrRq0EJn5Sgk8pyh7pzExN32UO5HicM3/eKoOxu7+3kgvXNOlXgVFBInAP/uN
Ssu+EseZPRDoMLta5jW8YGt8k9ucQBgMmPlMxNoh0Ae49yfSFe4wnZlmhugyoDqI
bFqZ20/fFVI0tH7IeOehW9l3OQgPn9A5gLvolSbHxjAg3Tj5n/AS/rQ2M081VADm
hBNcZ6x3UfsP/8yQD/LaMywv9MFakiatUOlO4jk8Ov+dY5OFZPKEaeXu694s6KRH
K3LqwcntvyNwLLJue0Y2DwJp245x08QRXieUzlcsd6ZvgFEebeslP/Nwo78IKjNw
OTgy4qAuhzSX1QuYTmnODqsPC1IjXYHOK/A4vFQjaICWq0z8Pz3gmnXuVkCD8IM+
QUM9NJrOM4iarjXWjiPFrVaALxM/I2qP9Bq4C2KkF9NmlPpQVMLqDULypS04xGAv
gpP72R0Y63Qt6znJfVqvI9Pg+aycXubZmEcdHoDbdwsDOSMJrPqt3HVRmp2MguZK
whH9OY6V29z+HfTRFBDSDf5OnJF/zj+ZE35RPGkAhByrORWMcxpADwpLCiLRNF5c
WP198NRJ7Qms2UYcCl7DJYK0MZytJU5yEiXf1tX6l58XT2T95TvS8o2LxXcgpM/w
Bff7IQXVA3VRpTOtIHWQ/MeAZbjJ8OjGOR9cM3dg1MDBvXi7wbHzc5ictgsECqJG
4kq3zFDh3Maz2QpkAveyAbOT0wMsnl8leBHf2FrhfblmrKAH65TMIfVOGcPS5QT0
ihvWPXDtVeTpn5pCAI6LF5z1sAMzOSMnv8v/zNYNZEuU2OtzGHAHZTnpn3h6kE/+
B1Ck9zJn4UcAUFj5zvY4c/r8m1sdRmsxXDFP02rcF0M/dridHfsFgZI4veTy1X88
XzUqVavbvNjUg7WRtEMQeVJv9AbXIjylBB0/VxZW5CYQtR3f6/sPJa2u9x46DU/n
o2C5tN3h8XbxTl7SHMpJmzVoRNYqw4MBfxxvheBpJRfDZp9fOQ+fxeogTPNpxslM
R0j8qNMaw+nOlJ5b5FuIue61M2W2dWM+IPm4cs+WCSJb/F0S1uRkVoQPnf411eqj
pzpefPuINrpzXRnpHo4DNvwcvq96esnyOEy4yD/qX6o7q0mTaeQZk5JcjxiHozR4
YWfamnSAe72VfyWK27V166Xphw+Vhhpq0QSVoPQ/vSQfMwx96hnMrYl4zcmemZXR
2ji1Uo4QO2C3qywifJuwc0PrtwmZyHRlB3Wmnpxh689XjgrawPVx/Lc97hiIrysp
KKXxTZjeR+0jKFbrGGLLwxidm1TiXjcSkSaouC22HRX3Kf8XsrD3FtPlbGeEIJEZ
5Ip9XAg5sGjm6TetslmUox29HIGRcarYpCtkrNIyDhwHmBv/Z49Ik6610Calyw+h
oX3jDwDY2hvoNulKLDRdrfkNyhOKlUNSxmvuHFyZuk4b1QPuUtfrdVuXAOV8sLps
aOy/y3W5XciYMdGjoNGnFI0ngPPBaXdZl1NeEitGdlCqktDcJ1OiY2khe+IaR/ym
VLUsU8OswBVoSy44H5FIz7jIitQfBGWA3usm9abP8ogUw+UL4Z3fH6amOm+746aS
XziU+KX/z7hEui7T5vtqYcuxTNA6NjywKXzI9wCOvgzMtcH1LWiI1eawO9lJ1K9w
nzgj9vpyiSKnR+uddH7bz52LL1phZOAZv4ecmJfwniZnTx9Xvpzui1QuK3AI1cyp
HamKqv4T6HKNRlaswAbAo0cuKsyQb5pKnir5hWfhNWaIDz0HVp8srji++DeRDMGY
ud4MpHPFb+F6ufvEdxKdXgwaTMTR4Y2RVIkvj/AbSdEgMFDMZjewmrdzbi19KhEM
7152ahzVBYszIjkr3x6OSXZ8MuUvwFRH0g93n0zZaXHMbPcJECJdNvjziRPVdXvw
AP0pF5o+i8Cx2fjFaCW3EXU77iLsFn52u2XvnwEy0LgCFV4fbuVwkHgVBjB7U6h2
kegu1UqJS3jHcUAbcDRI9x6EH/sZeXLoB5eLHDqmJeFSvNAjFW1wtuxAdT+RcpWP
yQ7y1MMqxtReNx7LBHniG2k88QAMfD0eZNFZz/yZ7+R/HGwnJiK4EHcpnWMOO+bk
JB0dzLi4Oj+g3lZ3eYdtSgECzkivMoxul1Mae6sdxNcMshwizV+huX0LXqq2oyWz
NNkrPG9cGJtUyRVOUtQ6EHSIF1Q7sn+xFFw4fnRbPFkKXOSk3NTSfvxsVqYZeGKl
ycGnqIDPTvei8gjwuhrbK98idRBiyKnak1Hk+RP4aaXzQUFuHeECCLOlx0HadJtt
r3UKfcI70LrboCXLCF3mx8t+BO4bgj0P+7iSryrDNqfLqL53pZTc3wGI4SPhrqzX
RJpYYkaRe+ZU5m8iH/N6KMBHqKbPIgdSGyq/xRyRoYAOjQ6QgD+3vFjpFqeseEuq
1wUFqwQ+dYp2lzxhgjAeFvh1bLVDBtxs4yDT3VfpyhNDWDpBx5kjPNyTOB1RI1vP
JygRtANbnMkYUxKTMxz6UM8bsY21wxZeSjkK63VogzKQT1vyMKc+oLulDIORy9tv
mHR89Sz0HPrqyov6vi3a4sHQEVQZPOur9tghuia+h36wymue4+0QqAD4GdFusyIg
rB8/AUDqe1tGugm5oc5O3NR4MoITM7RQpqX//zKuGV2EiWJPUUY5TvewDJfT+tp7
7potHFgoOoIjgjI8gn4wOw6MlyGKIlrxWcU5N055URsvPJlagPaPAznnDnAMXAjU
uaVukSs/7CLKhUTz6KfGUCX8UHUojlFRdiNDIwbdS20t17mODWc2D1i4/uAAUNEn
CVP83IcH7A0wDN/mYGmCXf6z1xhGG0HWJe77vAlKeAaSwYWPW6BFQAtY7F1kAt4U
fMOuNqntLCdgTO21Y9J7XR+E/9EYZ/mO8gzpm/KGwGki0sYfxZFTOHUDi/TBoPx6
UGnLBnYVY2sHO6x7/FanZVZlI4MilxRPSbsLXq+5EJF+hUYiaCWYw4dhSLM5oh69
oQlGxkInfy2lrMDGUlP6Hhn4RSRD7W6AzSpoIZt/ZMbYiTxkMZSZPO8m3lZNb9mY
p07ZaIoYLl6JVrcTjiFhcqOhg1e1lXnhdXSVV+xrznmPfDNSDYc7XyRoMihwWuFJ
HGF3jgb+tGuFdcwKnIwI+1SUwlnZBP2ChFLoO1oR3p9z2YP0eBQIcTTWqZR30lvR
Y1upGdjJTma/SOQlkWsl2E0WPyhEG5EzsLygmnQ0KvOrcyrHD4SjV6zVe92gJkE6
kRS40Cy2+mfYRrLreVDtIgxmbIGOuW1/Z53Fj1pv1Mpduxf87OT6wqGdcGCSygtO
as3ZwFfx0E/F5XqE/P2FAuMbcZhyYreaIpBtEN8IU4XFFIdTcJKPe+ixaq/jMw/e
tDJ1aq6u+tfuVSV4P5E01P5YIXLxkgqYfX5BNSa5MJnJHZAj4Ec89K9yHsO9kL5w
MIrUDXQBWP0QMkZOi8HKQBiBnti/Fmm58NBz7eui778ghHnjuA6qvixOTKoQG9RO
juRGp3H1MTdvDGMe8WUjPlLSNuy1TkTxlfKfjGJk5LyLFkt39EeVUWiuTETzx0yf
rRLgGiUuQAUdge2Y0UIliEGoec98/EWFj3wZ4rCxwgWkNhTGVjfugEejAVcqpyhy
Appqs8Zb5KvfjiNLVn3CFDtQjQRv/jjq1kFmHDSpBuHJijZPP78qaAGTBTtVbHSR
LKYqtdAxULm6v9bFsyiRvt1Fg+Tj4S8UCaNwsDXCkq9G/uEK4IpCb26KJUF4BRyE
8UyWTV9Ivy7M3MWWpHO8egn6Px+LVNgYLi8pcStoMZPhv/gcBgRWKzYRri6+/cQf
b6tBpKNpU34kb3qF3mxrumRMeWgrQRLchg4wc1YpYHfo2MLwVK9e5Kc2rBS255el
qxfXOPHjtby0EzOJhd3YOUIrZxXvT4rH1FcC2QkzNVC5FIa/gfPkTKjku6wXnzpH
dU9f1OD711XtviKke22/8k0HSrtzBblC8Urdh+oZyFHEyru/7YVlre30itYDLT6e
sQbN11IeN/zJt0Rr2mhQdrbHf22My4svYw35CWh6zfUZ8OKe57AvVcHfa6OS8wjF
eH2qsFrhipOndxWYPKLCXjALsetQNgdS3awX02lMF06y0w4t4Qpi19kLK57xU3wJ
3ooLg4cAl/3ZOjdcChNz9+tfJsH+7CBWyYEruoQCAnVgoq/phymRRzfb1v8wEjMl
pYSjytyJaLAqoOjtvDHmsCvvIkGuesoB7Fk/oOuTFejtFFcaxMIgkKqm/U1WvyYN
gIUb8r48i7maqc9YSw9FR9Bu9gSjPECV6Ff8plEhPEZkg5odi8mwPPn4KeC9gFoi
QQeVhXaUeSnJd6HcG4HBwv4S7JbhsCAiBt92iqf6bnZ1mLDthwPqOq+4bvU8pHpE
Rm28DHigd/lLgPZLCIcPshF7EDK96CSeQ32l+6aG8L/Q4aVUPsOxVSUz1ez79Cor
xXtj8syKKRx7H5r+ygcfQc2dpc/illOCmq7rHrfPjf6wH2K0MKMkfvILyj+rwJiD
Ca2qaPKXin1mRT/qKm56HB41kfR3TFlmzsT9gIuH3lX79O9MYIL3Y9s1+yXTykTb
YLE9lp2O1pQQE57/DdZYuJpXI+rodUCRIbNziiACFBZGlb4Bheq9ZU22NK439qyI
u9Cis4blkz7ZKIr9Jd9aWXEUPwkiP9ukbTctvU10yG66B0SXKWm7s/oPwA9nCvEx
2wAfWSEhyZ/aUqDi4xMR8RJm6f45PRP6NBno7mfwRnz+iBkcZ3PlWceHF/hNp11Y
4mcgys281mp4kfLSXbGiyPG7k+4m5bgF8r4WrRk1t7rUeoPwAhyqVaqrtwmUgDLZ
JRsOU60pJyXnajZ4aUwRuYmtMGRmgv96ReDvyPd9XXxtjkDgO1yJC9Kpo31wJ894
mcE1qcf/bTujCB5IkxL2q5/J73Ifo0ssSDlHFXsKN9ojUyDApDSXGYS2zYMciMRL
/C6svQcodsM53O6gGlAlds79bwTMAb5sFKKa2+3uO2coe2qxnjHGew0Fqehp7nCX
j9Ku/rKiFuvO/vt+C77by3b3EEeyp+NY/2N7JryClCGLh6gEU+8toO7imkVErt8u
wrkFQjcskfwVTvwNwj9qtr4+b4aJuQQGe90w3Gjt+bX7F8Voga8TE1qk5MjmdeoC
x5J1ZAEPpufJEjQqkuFxYOzbz+YkCSPA3qdqAPQkyqnZH5nrwaTMD2F2jTiuV2zM
eNwmKNYIlfX3IYLMDX7hRHMIMzKV0D6BIFFFwBRn1E/x1nsn6tBWVtpagFU++2f2
tmEgpujipuE+o7XlI+FEawP+pfLhorT37nKW3G6+CoO3NOE/i57U+MNrYOAhdlpG
aOspgCOtWAD8RdFaZ2d57fMi432pjJx+8d66uWxJhmjB4JzvmilwUySQ0kJ1hV8/
s9y32gGKcWOeOpPGheclX3lXFW6be6uU6jVCwc09QGbOE8iBxK2jbluUyoMc6YeZ
xCyUI32SA/S0745PuvXmpbd25xwjhc2LH7AYSFQeWGmLhFowaqwIaEBIKTGUKTjF
o+R9vCZ1721v2kg2FCZvMJrJvrpEY0cnnWOMiR+xZGshGvgpszhcHPt3Nj9/lFGY
fatgu0rqOdlXiUO4tbnXjKqIva+E2rQp63hwrQdE3yINK6wC7oFtS0Fz/8iwSQgJ
jGvHqASvH7ccHyXQZivAI+9oOE8Tp3+PSFCe2kq7ILrhhfdDfeLBKXLB10oG1Ls2
fQ/9NmgFZ7gThKWwGIBZKWbDMHmNUgbtAsp2jTyuZXPHW7Ro9IkAkERCMjPQyiTz
o0w7TPSQIg3XDXKn90A8g+25a45MPCAzze0ATqIepFhFftoQdpqX7yKi9QnSztvE
NosxRoTwYEdvSYGhSojT1sZzXMNNwxi1wWIY6LPYB7noMOn6GxJFPd0S0fpwWpnS
HdKK/ZEvmYtoUdgyMfExpXKxDAJZukIl0Sw6FweZc18Qyql8sHbIJ8tJdEymyETo
sM5eEcyk8zcW1nNRGRn/T94HgWMOF0/2rGJzasvhBvBkXXSc+lowbCgq+fFUEaI3
gx4JEhJ03+Cfgre2kVeAqZ7huPUkm5e8zm4ZjvAYKjGY4YFXgVI56FaZLOE1yAd9
C2zCTrcSSvfNwG8cu7BRYc79a/9hn2GG+QVfZT2tZ4kRWLRclbz5q1nnsmnHt4Xe
co2KxUHJHko/rY1YOtTOop/KNMjyWVKo/HzJctTNaCLe1iWiKPcLvHCzpv3sz4sx
qrHfetQYKoaTDAy8Cfq6A8KSimcNsaN+zkUTGPPDzEkEWIW2Ob6umox/rtYPuKhs
ASWOZxKX7xdpdoBte1BKLgTcKpQMQpn73sm6oA8C3tyYJ0pjnhgFrFKE6w/Z2BeH
HUzaHEZwwHvXy/e9jaATtdQSLSkpEWwmZqKz8Lw3rorPrUYzj4VFTBXuR4XGkpo4
MI3F3z37rFwJqCUUJ56mrcvOpU/GaxjAhAXdh72eCn6y1zjRW9Bc+B+DHn4i2ty1
k6aiyciIgDbXx7pXLbl9U8XxeG5rWkh/WpdW/vMEs1EoiIejH/4xPKPjYQupopTO
jPtHI0/seO8QDtpw3QkEN+Qho8ADnhZmf7hVhNGa+gOQbnBnNclvmJXZvYH+kS2C
X2ik1qwNlom3X8PWT6q1479S4CqgcuiInfhsZDN74Jx1kgoPjw5hBzT/iYc0BLqX
IwJ+djXvHqJ0XPJAFgO53Vr3dMXoySO7vSDjYGvl7WudYLgQmZ+dzQD2rXjkankC
XaX4vBrGcF0wprEzh8SixvuLCJliG+Zd11lNHmjaGi8m3lfEhTxNvqPRA84v1mMP
OeAdASBg2bxpkmLgvWqVIypgM15uyBvlunb9UWhx6PseWhqJrNsOt0fBK264kM/u
XvfOP6btL7JUcCfFnhqC4f07lEVvvQQDVo7JkdjHzeYRpWy2f1sLvCaSxfc3vV9E
zqKKZSkvAwcqUiVuFVkHprbv2tsLRrNLiKvuaCKk9TqhqRS1mdUrN7+2IM/cu8Dn
9CqQ3cRTzqd3IMsCE2mIDjcAgaM/fjMEaKSps3/PSX9GpM81GgYIzJ3uMQYO9hwk
fhcGIM+PFSbRDoqf6s7aYc0fhhV3FfxZ0GReqyWPYWhmsFuMTyFITcknYGarBK4/
P8cs/5K3M+gzCob7XvM/Acy2guRLVK/dl6dD8Bj+QNj0WCY3vwFaYq0cvJZceih+
81+s3Kb9swtrYrMRSVA2QbN/T430IsPJ92QfqNdXD2+IUvBejeWLiV/JqxHCA96j
PdLBDd1zCS12TFMwcAiSo07xtZGdbWi/WcIP/LeV6SZ+X5Hq4NbMfqF7vjDLfsds
RjGvPPYRLJysXcugsGyqulnip5x68jFV6lQRHZ+a6TbbK25/qqGWjRu4RKfOROui
wc1oOpzmGpWD80EMrzq4cNAwSx4oM7UAdkqVNyEESCNbV3G0UIP3tIAn4i8zm9yA
u7bate/mLXI+bwx6BmWHVphy0gIPefKYRyK4eo0xab/qcTI9rs8ShbkQfvbVIAb7
65V7Zymh32nmeapiiyoNk78az1T5Q7FKI/Z55/m69dTAuky5rxSHMUeguqOsA6U9
wioWvitm1A45iJzBo5R5BQGR7pL+0Z198UiufpmuyQC/QnMiF2Ct5a9tsCCZbnLF
f8sSx9QhoLp0ukV/3LivjPJT7BP/VESkm0rYA4mgvWBv6rM0Hd8LxDhsKCePUhUp
vZN6BmY2iw9/t1f1r9mYBAnvS/lt54lWOAHdwhK3Mwg8Tn+oEh8qXFgr4e55s263
08jy3ZmF3m5uwop6zFeWEMhlhdcNUpXSjD2FYZ1Gws/1NDw1ISDrSmtKmLBez4Hm
CgXK4Hk4Y4Z0FVhLY5svCuA1pZ3lPVh3dS5FPYkdVuBvkJdPaCKNC23hJoVrrs8C
/6DX8O4ceiKmL6y1B832NG9xoXOZ4rvk9Tl5/pT4qpV4t1XfTOizFAIgm8IDdK1U
6qM0eR54AAS+k/tmhrLru1dVJ4GyGSieUrkgGh+pb0Rl4zxV04R3bwHPLNirNP1H
AaWpOJqn7M4UkE7DMWVRzxtSI9xjpziDSjx4/YGdxYQeirZW7VLIhxvAiPDur5mT
dg267cb8TeS5hd+sQrhtmnsti0tweno2QmU44M5gLNr3XSLxIl/Xcp5+2Lc+wZVP
qNoWWierA6HyA0V4ZZgjsVoDej1AWZNb0neD97x0nL0n7PDa7k5YuITTLY1FeMAk
BEowF9yIP1REdUftHQk8wBdh8EMHU9yDcJ8xX8+8SyQp8kgVxU8JaE5AUh5bBThe
FifZljbticv0bzUIUJOFEBYhv+N9Y9KXJ4qocxKLM4JBUBooYiZKtf1Yely56WM7
QuqTAVPkAQIbP3OwUoc2UOaxxzKFYeTmR8RVj6FhXbaCyNIPKriUcktMv82kCvPO
ICucGBnEim2/A0P6eHFM5HFa3ZrwtYML7Hp1MxRZpEbwaJu40PibkgeCD7Uq7r2M
eV8mAc6GAiiRjaUShKVETQEk8nEfv4DpkVa8KQLUmLZcXFs/pZAgxSxN3ERDPwkj
F109jKVqo4mYr9q8jaLqWLBELptAkGe+wjvtIzQxHV5W4k3iYMW65cPMTRfda7Vk
rKuXb1iw5HupWIxYqdgvKSsbiZ9W9QkYndMvwunHHE9Y/puHu1A7nMZ/gZ3iKoyi
h3qk4Sh/Hlwlqpd2YEDPbN6sf+ctHFnwIOm/mpMpxhhlcDOsWOFyx2t3urcJsb+S
jB0zX9QEmqdfCrqj5iaWkhKV5f12h2zfRIb2BkRk742OllTBvdk7z7Vt5YmuIf7K
6nDuX+iesB38sf/AXUWcawb+Yr+4zf+vk6ttNmWLveo4c+eyk/thg2OztlD+xCkz
YvVfr+O2+wZoqjbbKIhBljTnRdOMVk+X1oXa5YpPMGZ7Wm29XJw445VLV4CESZkf
R480jCVa/NpC1kl9mcbNfk0J8Ha275HLSUQKGYu0JbWJLwyv0scUIr6dow/NPHOJ
HLHWPYahQfbhbTyYyHkYBHjEGukXdE5JSi5NgMq64V9WyzeH7OgUGgVXIuFTJeRE
P4lQTXDCFMl3Twcff6owiqnJC5OQAF7fTCHI/pHYd/TQXyUBI31wN5h8REUZW24n
EpkGREACxehdP5sqiJQusgUA3RFAPmaSOzxcJORXIb25H5YtGUtyEQuHP5Ryf5ve
174965aAkPI/cxnYytuVvA9DDMYwfCvVYkbOKiuCihvf4qRux7tw52UcHijy5uxy
XZ5ce+CX1FQldR86OoixY3eCaekQK/d7+0m1tCWsIUHvoIEqXjnnLHFwlXqkIUaW
JZh1CXZpbsX92/j3BHTl8WOqtjSTiwKP/OgCvgo9O7qAxsJl+Se4JcjiOlc3A6pT
uZja8NPX94EOCKixN5LNPZIH1vU99tuF1AgEscjpXqdQ3Jt/boktL/v/B541mCJF
R9XDRGBsXnsoa5vvp5VV9abOrRTvRCtyQqgY/yZ0TB2zXigAoWmJ+QAUZt1SYY1v
AhqqNCWZUvsx6zPVcOprNpjxxFwMXsS8d748Bj4K4f3pW6Z59M+0lkdQ+d35Pihx
S2AIBSiSlY1ZMoheG6dGYq80EUn/FviQfSa5YNsqAoeGrZMWeznw2CCiMYvf7Gdg
9MYZI7cvsfJo8/f/yO62wFSelZpJPm7Yp4Dz99ncwx/SR3/kk2SA+Sq7YnDL4+dQ
p3PneqxPGvqUfVSJ++ipRXAzXdlC4aXwjKV0U9Fson68CrqwX0Q3pZaB6b/IeDOR
DJIR998flsW0vn1cdO6D7o3WmLgx3qZF+1UJNHyYg5bpkG3321qOO9jSh+bfcFw1
Ij8w/TI3xazNjbpozHhSJCyLtMNH/MHqlqxhx3JMWHsCi37mnm92DDYTswn407RT
+Bg5j53xzrICvchUQxuBT4YH7ONUh74P5dYmufMmG8LDEnbp57qOf3nkGPOKLFKq
1pyLzfdtmgFuqJjRRxoh/e/Ph38gn3q4kdihYPSkq3AbcV0t4j7WwHNXeFQy1E6l
FUhOFe2RXM6Teb5EcVAObaBosG8PfzjcR9TrK6TJRpeLU+MA2A4b2NzsEC4EsSZX
M7EZN/wD679prSbp0rq8seprHKpB2IVkH6PJDS0hB6d/UUXu2ofkin91Wj9i3r0Y
blaZ2hRBWeEItb8BxyGXUtJrG7T2e0JMHSLwzu7Kwg8Yyd/BFX3l/t1j+iER+N90
rCoo+x2QRiAo6+IjIiG9+jRsx6OOa9bVBHz1kwiGY5qyY/OfnXSl9hLnzQNFiF/D
jko2TLwTolRzLjd5TTLGbD4xMt1MeZalm5tGQHsI3am5wMXL7PskFqIKpSB23dK1
vQdzQHhija1k5toH6k7skgZk1MpSA7lyYC48FR5cUSu1ovEEW1rAVkUC8shMtw4b
ln5X0ozqrlREM11aE1EXcRmf6XAZ0GEl+MJMJrq3H2XUpQ6hcc18CEdzYzCFhRaK
BTaF1G9r+g6T98pd/yPg+EDpMzZHRuy3WWZu7Q+xnUGhnYa2RH1NH9I0ZEgp3HJT
HLk0WYqsWUudBFuUnV6gN0oPvgGG9lxo454QUg7AOQCA9m2iSnF9tGKFrMnXMtS9
7OdkED6E3jGImvE9/gjpy2WaXx4MCrdFtbSPGMBDhc1f14ZMGj+Avt+OI9LLDXpg
RjwkSBtj0Iju08BoXZ4JWOhv3Xcxlzm3CLW3pMlFz9nMYA2QuZxU90Bi6ZL0Kqeo
xxM0mnjejn4VD15tjW0drl7n75+EYUCi6/DE1rye5W/BH6sCP6aI8L2WzMP/EKYk
hb7X52msAJSMcvLOcuL6LySD3G77iPEx3g0dRwgFnOvG5rRernrA/YTBauyv+J6W
RPfJoLDR7OlRvSs7UYDJB1pEA80cdzVt0j7UmcaDuMJC4n7xZ3wlZrzDBsUJNeXT
YGpstclJs4TXN8EmYqscqQaYDuGA4PFIjESPL9bOjP3Ncud9JenfjWADQZ9vxR3C
za8zke61OKCWtxQC4Q9Z/Vkpr2cAGXjRmPIpdYZSHuWidaup77j6oqvVNbVYoi2v
HbAEweNuArepveB5S7WSlIdWsAHE6+9YLeHxQp1pzAiGe8iaa4h8DvTH8R5ytiOb
MBJj4q7E1WqMFReUH3nsK5Ml7hdWRPRjsb26Q5qGpK3PH5msEvY1t7daoZdxRZbK
eOX5agEAxAhu1vCAafP2VK8e9d9/RRcYJDBEKeJ0EX3XJwr+Ara5UBccBqkIwf7o
H1MODjc5qyH8JmcR8rCsEwA2c8K3Z4RZKihkZ8gHnYbM4bVitjJpDDPlrx/qqlKs
vFoRE7PVt/YVCMhT8PKNh1gDRv0Vj+c0ZQpUolZbrLhzOizZYhUlY6niQESFoBGw
PLmn0jaVEAV3q6dM7RA+yyR9qNMnt4N4M0OiLPCqXWN2V2OvnIKtUqlMoZDixO9D
mFzMXVtkobn76/wuBOLOGioQ2s2z1YKVpwT5t8xO2Xqxb68FDKABgRCOYZX+Tqqg
PRs43QwXFG6fMgkQcY1hjl+FdEgavijkBVc5i8gvZi8zRItPpyeJOHIS+lV2BCpY
3AAF6lMJvnrhG1L5kkUk/Mi+IqfHi8188BNGlJNvoOsQuRM8mkbs3XVbT6A5Vuez
xwPKl3jkDPt62rxG8jyqKkw+EWLC0d0JhuRUaF3oixXoGZG4cFxhcukVhiTHUonm
/5a2UJIsSaEItRZSaj3zMV+amm8jenQ9v8GySKFNm/q9fYQM9RDTsrQ2JYN+T6OZ
xBCCi2h4YsmGKq01DCdgwQNPnouSRrplXS1q83R2pYD18Pd3cBCo6yRrKrUgVw+/
FVQZJ1Frysjij6YfZ7tEvut9Ql9Ca1RUls6YtqWjZ1qB5vmr3kv4KoIGRpuRA8mt
sCG8DR1HgBNp7lLD0vHGF7Tz4/Fxg4uQqqqc+dIqteMt1x8cEYheAUWHRyOouFIR
GxaUVc6Z8NSB6+CxZcqkt6IgLjWh2r/jbEI7I7mJRfV/OarsEcvwGdH4NSOZZ3aV
c5pZzXYn8oVvD0dfJjgbAW5RTqSErV8EyPvtpq1g2bM+0YCkCRJQoCHpqHNKQVaX
JZP2XhTlZ+pj46H3qePPnScCHgcWOGawwpxVZ6oYMqW0129Ckztla5yGlMCwT61d
WuCyQIlYdDyAoKBlK/mxmxJ7EHJgOasYUTqfHEIyC/EHdukq2+0wiAMMe80FqLQo
73qPfN0WU3Y7DseNY7FzK5k8HlKhbpGuOAXP6xzMR4effPqh9jswcZhww+GdM4fj
ff6Ine5z2nGJA1G1C8p60M9cUcwMmpwlqerZmempGpV5jlihujcRIp0YlLlPzGr2
CTZUu87ekEwWy2uVpVHnXMiWYLBzBNOTxDt9XbyWICrJiD35aMn/j/ljvXTNzYAR
gHOMwHu5kCNEwmlpUSsEMgA7996xBj0YiJZ3avOdPWkZfHdgHnIWbnA8Pc5d12Gb
wFyH1WAWUdw0nlTDJ66NYXOSI0wPjW9U2I8wsh/BImivYtexWq4daZqlmY0kVyVM
Z9x/pPZ7JJjcKG/dzXdyxrHVdRvUBH1i8VSZc4dWub3VqKpntZY1ciSY4zb1zs1G
+vV9X+i7ybprqIhFE8tmkBmjV5YUoPKhRtA3nY57BrjT9rsnsVwuqAbMnEq42pvm
WIM9ZspvqpAlCX2hXOWa/r8b3yUcX9QKz4W9jr7Km9VkHzS/Wx85Br6najiuAC2L
Lh+XjJP/R9I2bjO9BhooQZ/w021On27Q61QPuvk6pbmY/zeC8NKAwqO5YxsCM0Bi
oI82FicAp8h4n5VSW+mTBtQNc25slHG1737LAypKQWc6Ox5zzAuQseFtGCJhOr1v
tVgHHY2oaxKx+OC0+BrgncbgReUaIGRf7ft/FDsHOGDSoaCKWlhB9oBMZ0S/q5s2
KwgkLggfMggjsKtx1Eh0SKCtcMauoVyQbvoU7FRvSLwtqM/FB0r4IUZsC9OU4C1e
KDdM2An9KAiZ3vgCevzS0zmxGCJwAOq7trioYCBDtRyvILPVbnmZ2j9RqPW22p00
cI8fDpsvjOhevoZfXe/kc/nCdXluTBOkey43k2Vb3BK8rn/UeD8nh2uKUKsNZNqd
8X+3wFMS3cs9vOPLio2XddIr78EOghtSLFSLjtfn36ds0yuIdvh/VCnc5bMXPvUB
VJcsaHBW7r9Dr02hTorq8dRKbEBmDSNG+dSI2z/4cA2s9OZVgXFGRE3EPRtWLlW2
lbG0rVECCrbmjdWs6meJKUwjx6MYBwN3svUK+YhpQiDwIncE7NZ+z8SONGaqikIt
4LJn5h/at1E6do7GoKMNZ8Yc1OXI6pkXWZRaY6L/DC389b3yUMhXifTlyNkc9Kk6
pPqbCuSr9x4pe6PlN5CBhB4PwOX6fOPJywXhlkdgsWQqz8zJjrmXVNaqQo5FB24V
keEalBzgxScp9nEXuCKe7vrpJlsLYqS/PtLBSF3UneJQ/ubaLTMf+V2hF8Qrc1yL
FAq2p9eCW3tbRlLN+VyCSUziW6HRQAFc6lukZ4IdhXihLu/FmxyNWIE4ZHHuYgzl
wHDYfAjFD/HfII3/TXkQyHW89/CBUzH8pimK8JdijZm9Fa0fUCu3odgucAfyUIbe
SR0VGcUp4rdLxnMC7zCwBviBSlo3WETBAZSyU7ypJwqc5yNo/BNq4o0v3J/7SP4B
+Mv1OfqYWZ2jULlD/5Nod93PwCwOM37e6nSSXC4VsOQdN+sWUSAQhKr/q+YqhFPE
yVvHjXHOuVvy4wcWhXw5jRnCPfJ7VZCVaKwLrTLlGkI8WXqtckj9rE12ElHFRCsb
VzOg7NX6IzzWfpuJyqfI9sQhPZFQGG5xd70JXgh1f63RcpNKyTqXn6dWywiuaRZ3
WFBO06t24otwNTRf/PwMux7fvFxsDnomFk5ocvXDvIlqs8mmVoLK0pWYxHAGfXni
8bmYWezgQeH5LgEnHSToAFF0ov2wpv7iQuMBjPq7bDuJFuk64hgMaa030lItVacL
F/jlM891imIzwDCjDlx2Gujzs2KrdtDD6Z/PUdzV1iesgc27jxdC2Au6qHlMorox
qTRx7ClkTwO/1LIp3NqA/R7LSB9WOzRb2A2iud+2PZlXI1LNDmj2fXDshK6nyUfy
5saOreqV2idn7SmyXgiIkwGUPo+30IoY5Js9vRTVSN8dW5owDaCbRqrK/3GkSsHw
Q1/w0rhODB25cBMw6IcTZWnz7+L1gbhBGLnZJmD5IyMpChaY83q27v/joOY68UXA
XQx9A8IWP4ixHnkTSzBMpST0PIbnu41oeEsU3rU6BkOZiO30pFeX9PTLJ7yjcPRl
HbFtxCIxbm/m6vzjWFjneYc9C8EOU+kcRDOo0keIX5TQgrXRksDd/Ci+3eElG38i
dSfq2XsUz3se2MT31yhGta7tDImUJhFNPndhaG1r65rAVmutsB61dYZUO22rnX9n
Pk8tRjV4ycYTPTODFzp5c7PDGSCOdsV57+3rfuL6hu1/gNN6yvgaDSYaiRXClr5L
C0RmdtmewnyOk47o5YeBGnuW4A16EhnI/youflmrWZCr1DxrM+fBkdkiTx9p8GvO
Zw2Fcyc6YoVmd1PqIinRttu7yrkloMsaZcXPYrlRk+0eYrejE0Aa7lzvIjKQplaD
R7QZgZE2vAVXyL+cJ7YspYfuaeaVQT1egQtcMbVfyWMic15Qat5kJLTw9BVqXeTN
4TuFvpoEehP+7VLf85kpFjh5g3ASfC9xwqhiIjf0+Er9xsHsdtZfALazpTv425Jw
o92dIy9qc6/7FrxJAEZ5HRLJ5BPsSfedYkOm4WGBQv81STjS4E82ZLQmFHyzWJXL
V0bwQSr+ZHCsLIp9cJK7DjC01oi6/eLKqWCUumygXyVL04BIQJL34OBjAZOWPlfM
9LxiA871H+87jQMJOBFPRCxTUDKLBFnXBGMiObzykCXsJ2b9vRYBoJowvpxeDVeZ
8ZSjGtll1dnNNimMs85H738UytN9G0RuEl3hF56XxeYkqBGLStrjsMzAMqHLoolg
OZbFmPEZjcNIeUI7022BbzVs+6gdQGwuu/w3bBae0Mp2G520V7hMUYNECZ0T/9Ju
z0waSLUKaIfcArzLtz9JFtLLucDFIyS6p3RR1DbEq8JKyuJQqOvHblNXKJgIBu5C
v7m0/u5n8WeDrJkADDMf6q7P4j5jtP23QK6ommskSPecdeYOeAZeRDvM6uH+880+
RDkdwXZRAkgI8Arko/GRt4F3t6wa6X+uLU/NH3+EeGmdzQHluvvHC6qZpgo0IIUU
PmYZ9slQaIh/h6N5agApi2ada87dIGxheKoJonsC/cr+igDI7iPLvkR6FR7oAZnR
1+Boy01h/nJRiHAH+FWewT6jqJVDPHlUEznKXJHqHKq9EfRew+SW7EdM3idncbWo
ySdRTClZ1WPoUZ1VvspBlMGEGbqtHSWaTKP2GHrZwjviwgywiALQdQ7gKUb27tLP
n2rTDS9LfrkxkIYa3VAhrUyQFAUSpcpVjWO1bGFp8krDt4uiv37rFDQDEBWHv2Gw
sBMW05P2nEPuxf0sTs6aGd+fZykUY2+aAree0b72SmwYuCpnhACXJ4fbyQvBVLN5
KvNiNL4lic6Vw/YC7aSHOfI8Lb4Mf1QvDfBtj6NwVfLNzugGVIidx0SsvXDAQpLh
/gROA5mmCfrUGhgwaaU4EBQQFgXanJk3zpYP/ibvp42taqmUM/hpvIYM3eZN67oL
DhL9HlfhfHHrwlz8u716TzXBUZCq1P78sHCTno3GCrpvQIda2J5QchcDt8y7grdb
hNqKzaB6s5wZgjSOXNooao9e8MNyVZBPyQ2rAg3K4PUH44KHazLk4vo0iWmZDSJU
jubvJPIUMh6xIavp3LZNSy9abxwgknp2iUP2N36pLjWcSHbSHXx6bBMbHIBWDAPL
VI3SHmomHCGK/JPfAJ9wPMkEFJ7oBlaPEQ5Kq9vEqbRnQ4PguPcSYY87zOmrBc5Q
uMMYfdBe87h1Mutg/EbARruHXjxfpBRg/OPN2oIdZVk2m4h3NTWwAXjYhh/AqXpI
dF2hk6a+NFdMvOjlBT7NAQUoyCRuFMOLFpFhAbEp/Td42vigpaccmbZu2QWm+OWj
GMUQWWAL4B7GxSXrJ1jMT0o96JU+u03q/cYkiEOPS5iHNnAtCcipLDs5erUlmnYl
2jhzywGfWBAc7rKfMzMlS3ib9FOS0z6FPUeVKf/CUe096Ir2TSlxcyTD7a21xlrk
RQAKvTib/UDJJOQJWUEjSPCkHjdC8ioCJ7UwOonoC5EQnYYt6a5QZifpQ0Bt4XNs
K5cWkww40yQ2V/TbQdxXTvKvICkqvayNHnsdKNM8sXYZ0pIG+ak+d+NLHxBZKvVL
6pKBbcQJLHDS6o2UDxJ+g1sxzXfkDLvkoE/tr2rKxz1lPTp10/lO3Vyi8OTUNfqt
A/wc1SqNHJ3lyaXc2MN1MAEsc9V1PN+6s6X9JnifJ5cwIZK79cNREdwV9wMTP5Yf
XyImhYjPHsBmQonxiM0btsslOcYcGpAGjbhZWYt3tnSMJFLeC63bFP30JMkK0LwZ
UG8py/cY0GHPAsawRCT3QDnl6kbwAFdx6wOsVo1Fglj3ksFZk5cNrQlHBmwLV2L6
j38A3dDdTIbJsiM3yr4RHrE739mYoNrluarraGZddEZhPvPh2hCzdQk3m5VWsQbQ
XkFcIjnFIpyUcgzjBNhW3BMALtNeNgLCrrso5xOUowObPQzB/9kvZiJ1rB26uNJY
Z8IQHs0dRPnXam0QcXZqTLKVspWwlEMEbZwT+aXW2fGRZSvEzDP7fP/1Jeux0NB5
hgWZPuvhcjjE3YYSQC99lfad+7/4wjB4JvmaqVb9vSgPqq0YgUlWiohRAECPP46c
FJJ9TRcgBcjh27po1j9dVlUewWdYuE0uE59XLUL9+1UNJ7i5BTzfm4qOqLt9KmVX
LNdbnnbgwJetUyn6rnEihXb9xZaa5Yc9spkEcy4TozWxjB9mqdL3/n/2v6pc3WaR
pmQLG3OxtjD0dD5HiWlElSFrrOiEY1cm4l4nbHXf6+OEHdi6TJIM9MoPsPy1IveI
YQJvcveQC+h/CNNweJV14LP6Z7c/FKC56dGdp+GNCHWnHPEFtfR5TNfZJ3I31H+W
WyNnHUNNNjSpN4f1z1usVR0ae7r2/eQwrH6wf7bQc+bV5CPwLLNZvtqrJlJ8ZsQy
yB5wDWMdKR1bZz6nzmaEKcOPAmcwzeIfx6yS0bJAxNc6azOhIbZY5KyX27pq7G2E
HIUnr8yFrUCkM2KufHWxOXpsvvXAj7A9zI2i1TNpCCpyKSRxn1UooNfXE/SNUoBK
MeR3p+Ga4un3M1alb3ZBnrM9vY2OdYHrTNXBl5EXOT1g3flwKcQETaqSIv4+uwX+
bLleXK/fCL7lFihk4i0srXv3m6QJoWx5caRmR5KHeGJ0WRqrIB7w3/yYSWA4HUoA
0tNIp8BqCHi0C/IaPN58PWTm3bpc/KtW23f7m+kSDfXvaHcs386dAB0RztskW++0
DoajZE4otk2MgSvHr7u0LoDFnAOdnbYEWjRwkNUR9nbqvrQWb64ovmSW6Ipsabfo
yg8rJaTsszrIErQWrGC8CP7sncobTaqh3wyZoRbavTvoLMUxTzYC9ucVxafSHveX
h8gRxHgAAp/aorwQmY2EbMqYe78NIO3tP0nA8E04Yvyboro5K/MEvcJ8oSlFvrfS
BN4t2EXWsJ5W5aimoU5+82KMzWL+mAQmbaihgFugJULLgoaIeE4e6FACz9iMY6f8
KeNAGw4tmJLDa3TvPFj+J3PFsLzT3KihOZzD2agF0vNxEs/8tctOOnsKVQZt9oix
7MdOYFywdrSSFXnaWPozxnZy0oLRLAF+AMSusj3AMEanrWE8iW0V1ubP0mZNuphM
oXzNc+2aDpA9EsMexWKS7918Xne0gZ31zD/foPgh9st1dUnAMSXQF8IS3Onm/VyJ
LqySRcwDd6Tp1Ak9eLbxJMvGHDWI04DKf62jS03Qf7+zb8zms5HgHzNsDFilnh77
BqHw8P5zeFeq8tn5tUKqGP7hIwPtRdxOca3Z1yDfFVw22NmbDRL6hdftUrTYn6+w
/NAgspekA0VQLdxm3Ohbca3Ju3LxCSXYN1S8HIhXPa/MvwSJGiKycpkT3LuXqGjZ
fm2mgqB/kqJveUIIoQuOUTkYYGrxi0gG3z10Gs0ZxHDs5ASAR1YZZBdezwNUH3Ir
RIdJImeTz+4IobRwJlL4/0BooLqkP+OH2bntZHICWaWOKDgYEtHfUyQfywDrN4vs
rcXJ7A68+qzFe3rixa7JYy3SGeqyTbnQejKATTCr8M5V7ZmalT+/xh1ZdjZXuWqK
OXJIjs3XfKZKbaTomCCCcwcOGjucZL704s/hKcW04dbLq242B1ibd41/Uvq6XICw
6S6GO+7vRSgB2SuR4KuvxTdGdpIO4ZGpQ670OyqwCOEMC3oY5Vyx4xRst2v7hTEM
ziEDm8dpTSb5xgacot7+Oe+FnM4wTctUZYXsLMHpsieYXt+8HB8neSwB3FZia/DY
uZTaGESDO6Z2zBTB1DTv5Y/9IsTQF4GGEf7mUUcC9DUD/li2gPUwfnAxykdB2VC0
dNKYD36hWdpsZy/T5xezdSnFBUZyHlnApW3OJzhvPczyhKxPcTM6Pw+BH6l3y/YH
bgJXPJmClhmRxhMX7TsQgotQQHrtdhB5mFafkO6P8kYLnESpdiQiYVrSDCJR/4O/
DxmHHl9CPG9tjLeQLsu7v5dN2rcYSbsSFJj7cbw+As0U6c+xGblNb0ujmFNwvTYj
s5mgfC7kseZPDxRwDTJhhbJBY4YEWUEzC99oo4jm7zbHyHG8hJ1pID4Y2KeraC17
YO/xnJwr/i0SQkssqkSEPHGP4nwIfRWZYdCaQmvLXyKZFSNs3XqvXBBtIQrfvUio
hoTWL9gh3vpxJLJqrV8NkFBMlwn0nYUTTo0kjL1djL+geBfFHoznYH8QeBrwF4k0
uF+ovEVIhRIz8/IfTGpgKQPDPKzcx/kCtm54n5f3V8KJxq9aMqGw+8rk49GUdd+b
LsDQ4tFHQjh0ymRpADHH8kXxKUTBS5gGikJcH3Gu3rV4ffdzQT3QilOJVYoHJFYZ
qnBexDy95ytBpwiHVNpcMDtsL8zyzrO21dc6agtZNNPY19UB4teVOw4O/sCQdzJH
WPRHgySyK+G7xmPgsAJabBxuWDqAHQVs50A51lKoctU4UIqHsj+l+tP/5zaQhrXd
tUgMImgiWYU1y5PFwCK/Z9SgnDHiv612yuHtFTvyyUHrpZIyqF/IZKfkgS0CjSxC
FOiDmEiXVc5LOw6ZpmnOJHNwnfgo7Z1e+JXPDw/O/ddtZ8OL55fikQWHHkCl9kuG
za45UoXvHUtbeicObCXjk/xLgHurDAwOhJ1aUjvbubXZRqGu4ZkO2JfRI+wO/FAY
0wxd1ihO2ibhq2JkDtc/dydMAofQV5GFr9kH9Sydxv+pwHnLSkD9dY7or+/Pg3yg
Ia+kHWBH+UVmsHRH/lTU1ID4sJDVJ1G0hS/s6HVGb7kkANTR6sUXBAKjTIEdnZH5
4q90kxpMrJTM2fh4kj0Z4oqMiXvBmJkGhS1TOD+0yfnxCN0MqSeGJw9qQS3M5VPZ
Ox/ZwjybIwgD5XVYwpTpW0lbSUOKhJH7hZpXab9uQaWMJqHudp6iRkSO5D0jPtHb
9zXyztXxPDGAh3RIPdmX4MBPonIdu9a5G8WiLz97lYSR3g/JF87KtG5QbWntAOLv
3CPdm2cAMri8DZ4vLBirKWJ1kdvkN3nL71k8AKJf7YR8r9KO6W8u1i0Fp1QFVqYR
V2v0B4RKmLd0djSsu7rC+7suAYnho4hEMkrbIJ9cc3I1jR29W2yu3b0mIBLLYJi9
qOTmZQOpLheODC2xRrQBb5YkUSVehw878rdCuJP/suEmyKEBsYoRpVVurNiTMWUw
joSlay2EHiSw8P/FSGHcNhm1SqNV4KLzcbIHHi5ca8/BJH35aqOy/97/adbjNgON
KcQgADgKId509eRhXzF8AMuE/UMQ2AW/ANuW2EeX9rYVNWQj0J5Su8QO/5+XUhPx
XFe6LNsRv8H4OPzOuQEdT0/5a0H4xwKODnO5h19BN6lHpHsLcXpyJm2jExJbVUup
ujx8XRtjwW2bzCeFS2iliCiqMAdD17wxAdMxICgWVnEUT34bnNDE+9hqFDygmAsw
xjdxqk9dUDAAzrLO9syUO9CIZiMn0PRJ6R0UGSoLp325hD5CqL9nJDEAQNcRmowi
uJ3njuKJjI6/f+ehMLo/AaJR8uxm+kRqFZ6qS+PCq+F7GtC0chmKE2yxEjEqRI2+
Gr5SeH7MXEKiO6rEvgKAMr8jE5LOKylg0BP0pyCVWgmZ1loLeQa9+aikzXOWOwTv
4rqnGwb8VEwqsiryGeBXF4f8sQ7nEKjFp+E2oPQqd/x3dUbCmsMciWn1dml7FXRp
6XOIkl0VR1eoCYfQqvsMwOXG5Nobr8J5iRT3JM4gxTc81Y/BHmmXYoMefXuExqo0
BrFR7NaRYEQ0YWNJzEMbkt/3sINAxNnKnX5bj/QgrzCGduHypxygnNQvg9a79tes
FZDuFBrTJasW3aB/cegX+fZc6s2T3dUh4q6Rl/569+W5oEDro2nTPPCCblJe/Jwp
8oTPzJaJL5eF3UjoBMDnbfhJti7iu3NS/bBKEnaGEfoEmVvJeBFs6VTrHgdI6wYk
+/AegFw1z701aPmPq+tBdFGNx8n9cF2XsiIPolaaj6gA+YkBI++WbN+LDrd/qTWj
aZ0eAJt+NIirJBluYCdnDG0rDnVegb5qEQA8+9Ps5uBJqWGIVYXn/mtlblaMBBFa
eoRD2zqWhS6OicZGdm24qSjIP+t8ZxLGzn6u/pmlXscPb7uJiPLfrMmBDNkt0/id
EcF4EgNOXhZOYWP3IEumW9eOLEcg4W25JsyuNSs5l9pbaO6EBH4f5vz/tTVaR4u3
k/VamH8mrudNP9elnLk3UglxRHInkNKm3TZOTkQvu65DgPFNw1q7UguyWuoPWhY5
1g4NwNdTdQ00Pigi0/xee22LtWKcrX8bzHLMtxUdEgALUdWBJ8mwLYICX217Umhh
7S+pvnyXRoW+W6U9zaDuAkcd4Mos/RrKnvMEcBuOFHwofQvGdqmQBTKG2my1HaWT
UTSwLjS9wdYwbbBnAwG6ZJAFAqz/E5pGOnpIekw0ebPMcNsunSe/d3DNwmH7zpeU
QcaXLiCEEC9Tzaa6ZAS0R8M62TKJkziTDBUuVZLTpJ2KaH8MPmrhiDisA7fi8S1s
y1l1BbaTC4qI5EHb6+ywdla51GROZP8yuy4NbZKKiGsq2jhbABfqqckF/2mRVfud
/oehcDSWlnwhODcMqhO11WTA3Wiq0ooIIOtSVNIKlNpV+IF/4rqHKwJodOz4xd+H
Sbio3m+GIv8p1W5vkfXSvXXhuZliQD5ziF8Mg56PDdewD31SIeLnOFBK7qb0DMnX
ti4N+0Dm/ls09bG/3A3fpB53L98ox35UUe/66PulhJ8BBgMka50PxdYvfNOSw1Mf
W9i6SdP5i4AOOVqP3skiYrb27hQCt3EdBdVx3TBa5C2R/19j3bR+67KPsa4cLJm/
KwuYl244lkdIn/G0e92O9xmk4qVtt7dtOwVMPgb5e+mIEDdA7z+zy0z866u+Ku6j
62lRA87mnfRJUEYbnR7r5grBk9ZDrZKWAvS2uAiodpIifx4vN+YGWjRKNvA+/hop
8ZJlg6jtrtE2LLMXkXzc3CbWOXJGJ/skdoKLjXGbiP/rBVyefnWki60OYByJhu0N
nXiztmkCMvqPY6qSj4ujSnJkAitUe4dhorssID6uUh2CfkK1qMYiDtNsRlKHrVwg
v4OJ/DPlwE6C+fMQp6AVL0GP5ZTBAM24VyS7jYHP/EBb/qd4k71Lh4PD8yRcPKn3
3PHTnQZX8/scTHoGLXjDlq+g3rk3EQsR32Z/lnLrVvpwr7uwC5ZS8ic83/8Ilvwl
8Rkd6w0f+M+ns0gpf+322Brnd4i+sVpzZabJCSUCc7eE94yPkaMy9D+csPn1udEh
Iuxa7Pd77hd8VdIfezehS4jIParQuFcXf+y+2wxzzwsp+Zr11f//H0fPFjrsbyav
pvok/g5bxDTk44/zkjQXJuetfcJu6+odR958oLFn+mXI5Gl7gaxgUJqT7fVTuklh
uF5Qxd2wu3Psjxj+cxupbPkMc0yJRFE/rp2bZk0kwUseqUFE9vqDmiFB581910xZ
iiC88SV56Y9lUWTv1+AyGgxYDjlwoHTho7Xyj3hEabq0eKbgPyKKUwOxn4U2Xlao
oz0Cu59VFiSqY90gNMhNNjQVEOj8j7rdbFllZGXojUAtHMgyt4jjV/CwKse0olVy
y7oZNvasCBFkcmbrEz9n4i5jL5bHEi4rtboajRX9mBMAtv8JxaJkDUxdEn08Tx9j
EtqoeM4YqTZi/OFocc8WWzBhHu5U0Q7yknNHIWjLKVHsHRT+QbwfGYBBObV4GtUs
91BQ0OQgta5tKBJYD7mHx6QuT8oRqsoFs2N0f57Bhx+sGcyREOQFOj/DqnjXpczR
f4wvR/sEwAbGFKli3kL3IoMvXqr+7frCDAV+umvIY88AfL9YLB9Q2XFwWsQfNatL
ouzzfKS3rmQMOwrU6WgP3UXWR4eUIAfwvz0FqeqWtLQeokggue18NQlo09PZSs9R
SBEUOlcxOGzCbNRl5gGraiVgExDNoIW+nad9jg5NDxA7eJKl9AM5RU6ZerhWnMSW
OBF5xI0fcAn63HWqZLhO/FTq5iz3kpicWWh3B7hWbrs3pSfKqR3D1IRHCceV7xRF
tSim/XvTIcz0GkzxW8alfsoTzDCaL6QYduLL1SA0t0z9N8E1hb07Xw4T4h+htVrN
nKyfS2CPLeZp8TyL9qFhZzoMlZ8FKsqaUxTCDVhCV+3DXw17BGXqR3TWb38V8Wlr
nf0XyDSlEkTL56r+loIyMohMi2ClHAAZuf9AUmTOes8J+FiEp+usCRSgNRAMDFPG
9KHeytNF05nXdqR64BAMI62rJFCq+e+84Qta5lJaOEhGKJREt1Xed9oPo84R0bAz
88vBBBzyz+8P5KlRlMn/SDOKNOTX9SWUMiAxByFpWO3nVVQKLHvy7Jue8up+MA7H
JClW1GSgdOee/+ROPkERZIpl8tcNqVAZc7NPZ1BEQaktFT4V3MNm8lGUFkB0cwgy
gcjuiJbxpZJRuBxIOooxSwHvXZKb9p237Rprj+DyURMUkBJ3OW2U9q5MG/xov40W
XqrW6efav96qxDRXQpjaGk53ASH4FwhVYvlM97Gsa+ZVmkc9kDiBIAnk6MK9qTFz
WVGqK1WSsQd0fuFpX8xBThDFIInGGKI2TXwtpq8z5afBqbQcft5chWDcTCkCTJak
iN8q11OGDbmGqjg7vXdEzLAY1PBHumr0ApwAu3zz4zkq0Z/TOZJI0fLiQBU8yuYj
qET4+xuOf8EM5QbS2XCoRyON9lpJatvAJIjw0sa1nuYuTSYjVgwXPI3ZL2NoJLhf
pkn57wlD94DpkKJoGbTv4smqNUl8nOzeHec7HePaDHqZSRGxUcS1I25l9k+IKRl2
cbT3sCbIQO595gTEXSX04F0oMtH7pRxSJL04xI/ZWl/yBA8j/e4NuiBsLSk5lPbk
Bx1zyw3qUuXDLoBKIRntCEaV75xHolkiCzIL5n87Ux1O0M4odVH4wvE5ugWu/taY
/xxzdFeSrkz+XOOqWx1nZAVkBZukMqQAn4L+A2ALtZmloykhYLsb/jTkappC2lV2
/MmjRK/CCDtYGa+DPwXWQ2Tqb9NhY7oFINjeB5QppPloVrLQV/7I1EDfhX1vD5JY
/V+2Fyc5PD8zxQaIyxKVFqSc2cdyTvSi0PRxuYvRWzj6+TfS1/yS/cer3cvLzw/4
vLHytYAkqwJ9L/2gxRsrgqKpSuf5+yEm1heglMcf3U4kRhJreOirP4ShQvE0cFgU
f2/3FezEzUVKy8PRcvWMWJulSyTev2LbcW7K3hW4YFJWyM9FYWHGXC1+4L6tzE1V
P1GdSdbwy+usUwkkq9bG/dCHVmpiEic+07fk2bis5jrB/hkz2pMGN5QcieKF92rT
TKDP5reRjSTtl4UBzx4AOCVRJCxsnvUGhAz9QFus0E7RE4s0DanWtFCDm/xZ75TP
c5j6n1ojocAl8fsphIJsVbDYOnOXZeMo6s+DHA3ySSlh395pMJVSc9avu4aV+YOe
US6oJQGGKx1uCdFQ4ABKnKGgcgmj8ovThoon4ZYrsfh2GG7MVoDqG/JIDinThLsu
TjQhW3MpAxuIz9Y9omwCzc8+urjAT2KjLJ/xGkRlvajf5+S2/DhgF/1OKWIrYkUV
EI2LiXcr1Z5bOKmVqVSGvD9kuotVAmuZIxFLzBlhgD/XS+uENhXraincMyUtj9zA
MR0garOWgreV+ET1oB+EDRf5nc4l2bFeru1oGemZrPW9r4n+ATG4cFzGZNrM/Ycy
IZvrLP867cHAXhAF1YcOJRzK09s8g7XN+Ri8tKrZfYi60x+WHS4pczhxhlZnctyu
kMCFb3gTULQ3wP2lS7yr/2btqXBZuS83AC8YDOVLJ8FvK8253DlJNAnfViAzvEEz
wUFrhHs1nzA8H1rgJupbCpC0lLpnfTODbjB9YE170/wkNsLwSUahxf3hC7nu95CW
NOiMF4Erw2AVQ5/FWYf+m0sFclq/QRHj7tdi2TzSr3kELpIxHKGlYfryWD+aUBgH
PUikf1zYWKfuN3mkv2IOVO8b2MjVzrnTesZJIR5TYmaFCrYoc/1StwhKRKXSB1W6
sxeysdTkPKTiCgkMssU6o+H29c/2mhRqldk6tygTVTT1F/aNqU/bt+KSwNRBLVHv
4Eqp5i7vHLstAAGN/dljNvEwrmbDkQVLy6o7H2K/tnJkWCKvGs1K+s90414zT4Hs
lNI3lQGxNfyKxP+P7Ifk7+pNbru8v2wthQQclAC4pQ5thLRE5oUa+kOKnfu2tc0M
Aphm+uFQiBCa9WZPaiwVUewaXj14e6R031WCOFf6uvwp7Tauq+oFiCM6BLFny68q
rQ8Qzkeb3XC6JuoRuPTcEgqf+01dQYBJ4G1jHNiqphAxuEsPPru9MqSiYDmIIljI
SsgegiAJM8t6BM/aTe/38+khPKn9iXNp/yI+bZJopXrKXLBy8iig4rmansQ/df0c
Ey2/Ydn4MuTwPp3NrdR/lNmzkAt0kQOC0w8LE+oe5GiICiYBTB1XqC1M2tdeR10V
C1GYpO/2qxU7whb1C7aZQnFqMpTNhHMo9RDvyJFx9NsSYBmaEO9CVjVA+gkp9jo8
CKV889yQPc1efLqFVSu4EW6BApRnJ0AT1zPa0u8BsQKOFNayk07ArIlRaW+Aue4k
c/OgcIZPoIL2lL2HaEA5g23N4nRkt0/Ae5fKor49Veh46pF3TgSHRZ6rr0NeXiMt
586koQIJPpRtfThEILb64fcDrkyMyqDlXl5KHiBiyb+6tM6Awp6/bqdpAuwM9lLP
9kEvM4fVnJxYYV8Jt8AtlwhedYqVOVCbdg+SF6sdRNrt2oymLEGmgXMBifOP6v6u
6UgorWpHMsQB8akJwsg4a6zsQ4SjVHA6RXSJiGTV5I9RfJ1utMKg0Ey5Qi1bNDja
U8xzUgDkjz8yKgRPLG1fDqfneowVp46CJu6TedZk+2Wb/Gka+xIth5cKti4gPqXr
gzuf1NVAIP1ucms0IfjmU4k2RDcKKTmhBXoSJp5u81v+TU8t6roGikgF6yjS9J+o
3yThSsyMJnqfCkHU4OZkXeo3luLgpTRmi+ogblmZGfUQ4LHYT6x6oTW6CBnNqIhp
AID80EqZu4RZrmfgI9rbF7ldpgzCG0bi1g5quehYCUIjpuO9Nig2bM75NCSY3ecy
kUmou9BwFNlGsULRkLL4ZdOkX+QEnhM72IBFx0qpzy3PCmCq0soBdUkPyEDh5DrQ
AV3kLuYnvGpbIB9QQOR2Q5z6CBNLO0Lfxf6S+YKE7yHAKd6OJnrwiVB0SW0bYEYh
iQbCIDNiuk2DGHRno2cicGTtNuh3709NFp5OB0S2ousleQaTApZXF8T83pOPVJza
zSzjmor36e5p730QkXkEehsPSAOVEYvyg2+IvvqPLlaKxHQd5McmthABOh66ewS7
2mRwmMzLoPPK05rGL+pFpUUUtspQ4gQy18d5Lfb2/MG3GuP87SE3C+PhMHNoOnUJ
uSKH0iuHsePBCIGp9S8Kzf9xYDji6VvLFado/ggMIb7mxHo1CcgRG/C8v1LxBr3h
9I22aMB/sV+EHUZUWHeCGMvBdveceUTmGT6eMTE7Bl58Ex/arVbpqlQ8Ab5JMz0F
vUwZnboi5ev0Hygg0S3p8xXjxJB9kx5HkZ+EeJYjeqfKpOU4fZmzvaYAdvPMJreB
yqucL/2Lt4u3j/v6bdQkeOm0z5SOn72s1bUpuSDK4BDmXkNQnAwSRdWSxe1J4EHz
SP4KSA7wq0lIdwLqzqOwA6M1wcZLOMLPxpm9N8QXx1NLLxlrUTEJHX6z5Hs205dW
9dcUYevpCxFkZwiaxtF+dsFjzC/u94NyPAJCJZKdrKLs0QqCTGarjfJ4tYmYEyU8
aP7ZcBkU0A2g4QGiopHHrCAZWx2MUgM1c2NeZV9KG5hzQO77mkp1qThN7V9VaPXm
P6UutUXExZIsIs1dT7kKvy28FjUrOc42rQqd9dvsF0D89cEq2836ua1YxD0lupCk
bz7I0qVaRts9AiGXlFBEUBxqZxh0C/ehOC7K4myrCxd3fsfNFBSmrqS+7iD97J2P
2+/8+6IGIu6eum3VixYl6K6QNDLthf8uwJbkh8hfRfydA1OTV8hGWzTBhW5P6d0X
CpLx4NfYZeYCEn/gAYWckBqswOO5igtDTj7gt/0ijRzNqnteQs18OZEYBlQbtoIc
JJVvwqcA0j4e4Ub+HXOaiv4R2GXtd2nY5sDbFNYkFtmdSCIGEkOw96sy5x+Ywijs
uukqeGpYC6m1u5Ldqr2KTLj1Mf/XxSyZoAOaHtdnqJrhPMBcU63lZG2M4jQLKcR0
nGeaUW4xjy+/lix4i20U6TSIQ7qqubnUg+uPLLv4vidtywOMVb3mnTmeeevd35Y8
7Cpn4v1DtFZViTwo4UmrlqnnyHjUd7fYivCxTXQmPHMIxzgfyO7+G16a4VAXiPZK
y04XmVF4iLaPk5XF5qMmFGi4h1UFJfBje+segdcTBsWk/KBzHnRD7eJ55rNKsn1S
g2WsoPI/ZBflcUthB1cq0p0D9tqc1yc9Df6OT1Tjyr2HRYv+lvONVvia/jYNS5r+
QiuhGcGmoNOQuOp2uNimG3+o9Jrzcbi31pFoA3T5SNGwwnLXF6dwDPsNPw0fUcUa
lS/60rG4T1LYoWU7/lrEzwzdmCsYeSW3HDAvdY5ipkjlRuBjLUNbuKIZyOnRR0Th
vSgBUUupbnFzwrFk6KDBMT69NnM/gTQG9E3S8ie8P6BuiPr3pL+iIBqwU3qbWwdS
rOsgygfPwpkPhm5nNaxJ4ZlTGJWWwWJ7LDaxxFICWyooyMZpDcCf1ArL9oVRISPc
PD0UhMiUr2P54QXGdPDr3xsAm+bMWqD5Xwb+op3Vg4SbF8ID1vzy/Tb/qw0b6vZR
lqqvBG3GIkMja/pDC7bfCgHi/JmWtyMRBUzlMeCXRV25x0neM6vJJ48s5StCegQ6
ZkAGfUt1M28bkcy6ThLlBHoOXLrC21qndePqEAg74wd356jgA53q8sBkwHBvMMRN
h72xWQWLH8EQc24QTbai8b5nTyAhvDWyra2O2S+AMwyCfyyEuP0WSSqslIS9W4lt
cepoOMy23GQME22Ptv8114TfosKRWA2lZO0BTAgT5NoXqli01kC5iT/Rz0lr8KbV
Tm/WXJwOW1yf3Zne3NxMUsKL8zdSPdF6jX6qYC0b8L197ESkMtIKt5yKKtNHJob4
fvEi5UaT7KzFn3jWgmpsnLP/jqKpmfYN9kK+vpeomejCv8VBFLGPVMDzT4pYhkL7
06ogbzEONIhjzx/27N5wivTfaWSYU1qgMX0QgfwVKo9FOeLljgcdd1GCCAnxxhXv
S1QytEXcHR7ixY9DkZrztRVgQDQ9gTisUjSVuzVuqsTbH7Ii+Afy4PP7t7wTTd+D
Yz4iE6PZ82dKEaVkPN4RyNjvSTZzYNTY2aw2yEpczFPSnkfxWZWNTzNaseW9RiNC
tiG+DnBEKkAS6q75DmGPsTUztJHJKVS19rBJzEcKBEkCv+xFc+9tEGPJyHaJEePi
vvwvhZrfcyelcOWWwi7j9SBNwehhs5FWVOXNbjdGUi1niQbAlTAP0CA8kh0/vGH7
glVgQFjV6s7ATg6Oy80rTgMgdNa8yEP0oa4h0AQRIdZZvQdS8EQZuy0JMPGe77Nl
rbxSWbluddi0eihDI1M+9WqrNjbOAmG3zCPawcd6TSvOVL9/0fjkq1NLAxQ+3XGv
7M5F02u/AybpVW/v8wjLX4BuRI9xqCuQwa4zMvLtkXtPa9m8j8i91/jNRRBgNsED
2S32nuK/L9CesDyvGel0tznjm4UGJDpeLVzz+fGPa0wftNp/1eBxHP5AR3r9hP/F
yy9jOQds/7mBwsma5+0iJntxQ7UpCBkvjs5yOBxUQ+di4vnTVHNK08ZiF1Oax+ds
CdlAmRrhMv43YypEVm+OYp+kLnblWSDrgQAljImnsXhO//WQV7BPZVEoEx2p2LOA
TACrvLZ0VDFCzXmoGZQXO4Ed64vQ04WIbREzB0YnfHHHu9G3gqW0QL6HZm2/KVHm
/dGS5owEIsgsCTCeTBA3OBZQjK+aSBk5qrY3s1DK0+gORBUzVlaBY9Vnyq1bvqbl
T8v2HUfCCKgMqb7N8WsGvT5utaG3QOkrHkj9NLFBFPTPfD8PohsMzMUp4nGRUW5t
2J+vB4vkYM3NleNOfzxHgukuLAgTmkXYOofQheqDCIQzkOHN6b5EWa5W4JAxujqO
Ipal61CI169kZ3fHjM7tzjheHOqa6MECR3+BrZVvTW+Lrfq500pSGAEAbu/V1du9
OoLchKCpEYIpeCk0WT2mdiN5E/ypdgNN2k4jl+o0Vpgl9Sr86rzrCY8RAToE51MB
xZvHxdZ7XAXC0QD6D/cFCF33UEC8SlgSkXoqlBwxt5mVinSgQA/tbpFisqpv+a5Y
qdkWLOtGUsecsAEXfgxdRyYPRBRWTW1IrNxWDREDORim147W0/bk02zsMxQXDTMW
S/OAlGQsCvpszlHtJO2QsvX76R8lK/z4WJa6dCgfSOr7oD/YnjNhklDFANBeyW6a
jwbXWKHD0pbCXaN68yvK5DFVLqvFNTcxcwvs9hFKE4eTfcQ1Vb4LHFjAUXKoxzky
NUDloRjjOPowk6JWJoTlQe9oCqS/r/RmhYgR9g8S1nNeeLTjkTy8wN/SuGKTSw9W
pBs1as2YQoqX24beINeyMtE3Y/jJpPO6247rTMK3BgW4hi7GHukImCdMVt5Bvw2r
57FNp86Mpdn/d5iTiGEoseK5gGu3zdkFOVBSSHKGq9UFYfxvQK/IzzS8F4IKc84z
XTV/rPf2TtB3N0YH5SFMbmRoDk5hiMbD7i7ot4urMNx9l+L77bm3HwF0e5G62iZd
qYh8n5tL2MlEo1WZ0C5cE6h4dmj3WwxZy1g72NOtKHPFmgF5Mkpg4XuVl4giWrU2
ecXvtwt6+TlVx990HjbHgLNpzPnr55pXcWFMb+aGS6wbsmFOFjcssJ43qieE/o+E
znOBJJ+WlyEAzFtsnJIBjnsZsX9TVE4NLqBhjWY5EKPQoS54O2clKIFe0T9vYEv4
Lc+PuK89z1lbydMgyIiNZ1JfFG51A8lgOlDHPJMvszTnxyESWJInyZ3kfAyKGbfT
nGAW5RwymgWmet/kjlhsMI2iTjjqR1WDdws0jY/GftGhBVT7IXWwcLkljkXEErIP
0+R+FG5OtV3VrVoaEL9ixckzM8vizpgSdiU3XiVx2IKP+do7h6AVAvqkZWCdhcCM
hoUAVlWCOAGOFsnkPSGKtxlVBaMrKabn0/DT7OD9EvA3DjkHVGGZhddqFWPahkXn
6qPhQc8bXOfgpXLfGcoAhAF211QrolseG6SsqlEXV7M783/ncSsneEtC0fG+tx+b
2Og3RlmuYh9m4wj+MzIqMBX3kO62FiG6/i3cYQ8HcUXqVlOma4hnHcZxVU6jS8Al
Koxn4G69y1Fz40hzwcUpCkot12A4RDTZHHCCYblB6skcvFchFQouDxr/VoKs4ycY
o7YLbsPCzLzzsn9NWXBeUvJ2zAcaztcCHAVaEaaqmo6/4fVzXmePt3mTYIkTeN5r
YTWxYiKoCZ0IzwNrmYKjFDkcv4Cz3Z5oUiMhiKITBNVa7WfIuUc5JBPX6KecCwaH
eeT/5X1h9hQRv6a+YhFI8sVxqzzPeLlwT3o97V45DhmWzO1xS6knRohLFj3xfK4d
VPwSS06fnDHNss5eUBWM5fOeuwprDtATlO0hBAYi9jMsPIA8CT9VzS9c7+H6MXgV
4RUZiPGpmytiztIhb8/GM/lXVNpyBVo1WXP8G72GaWjVKRXnHUpKo6Q590gf+Qkn
Z9u8NICD54eN4q60HYzOIeC3HycII2n7dJiZpN402Y7S3kkqOOxfbyKCvuN+wsmz
Ax46ScuP1CPfqyrVzDGoP/RXzeB8ViLoRhxGRl0/HzME6cc8EtapmV7oLiIzi7LO
s+jWfzKFGm49/p/TRWcyLoN/m0CjSX2V2rNA59VaBMb8UsG9axcEd9Ym8uO9wtxG
+yAfsVTg0yy7Qm66amAmYJRxpqkaeIGBVnbA8uNJHYVuQa7PMX9MAyBIkomzxs1q
RIUSBgyapy8rJYKaBo3+/K5Xmz8uYeGndA8Rws0RbVCX5ejjkg2ntIojR40WZbaF
jHVfzyPHUPrI4VG9B8MR7cryA6CoG7oaqiSS9a9PKLZjGkD/ZwVGCZs22Djnm+th
14hH6QHqK3dd7/qKRllMxZCwg+wp1OBaWIX1rcmckyFEKED4K31rNLDzR9yRiaOp
DPf1ZJNuU+wBt/IlMsNFP9HpVKLN3XJ1Gr43PCCWe6bdow5SCeLQNGHakiUGQj3o
Z4JxvyJmClaGgMo+uHvGRtCGG1okMUrAffoYtle/hasQCAkUD5QbrWZ4/zKRwzna
niXfMjL1f5PwXDVCGVBbMq3YjrXr5ICeXF6KPPwCiO82JdgaWYc8qsgj7E6bcZrf
G6/EEbcYi336fIVjtJ5ATh9X+BwA+zNQpPRlanS5OzF5SHy5YXcivTWlSKU+nnzK
smHTrvekQ4wCpRZLK+7L9JT337/ZhadMzlCfPw83W5KyO3UTsu3utaPcqDG5NmDX
34qd1K1uzyngQAVQj1HQ2e1Gn7W85PASS+h7DIhorhn7BI5LHINqyxjM4f3jdOno
+a9suRyMWUGayb0Yil6I1k4jLzCTGC71dIbWfpGVun23jbxcZtkSmRziWdsH/gz6
D7Q1Orwfnl3gMNHI9noqmrnIB3JQpgcoRhagTOx5lwNEipl4mCvs3qWDkJxMA6em
NfW64GY4WooeODgDFXSkQSAAZfjMyTbQcMzMHfob5pD3cROAe+ISbNiwcBCBrfCb
gG0oeQPTBdV6SApTkoTwTLnyYPVAO8MHAG1F1mZ0ntaytuSZnXYIds/qBDl7Tr8C
LrjqsVLD5on6pYXLOqmqXe+0zdhMhRMkRS3yY/UH/3brY7rJVY++LIZDEeEINZEZ
rD1zOo80u1a6JqyLrmwtwTZtLg4dEItIpNzUiRhrj3tmgET/ncvSvhr1Mpa6SGLx
9KZ2B1FijNBxFSJxAmsfdQC8ES+B/Pjpjy0jE2QUc273+suD7QyJIzrBl09xgRzU
OZOxLV3BxOkoqAYuvX4c4KtxQ5ilu06lF0VoTfZhSKDcycxDncO+TCfCe1uf5XuL
o+hkpG5Fnkdi+BnKjNoZSRiXw/TNCsUvSWhQDb+EGeE39p+t5YQdVaxVtYVGnuwa
jaQpVJXxUj01XmsTSqBRKnD8G3Bqvzfu+HWXWvMpMntd1CiyEekd6Q0UhLgT/8Y6
NA9qWo7z/zXSZ72y16kUDBSBgvis1DrL8+B5HakNmNbvJshjny5/eXi/NKP0l7zT
tKxHCP5apEJMJcsoLpTn1mlkye3xzLX3YZsO0LsLjxDv5iECDtwwRLqDt60RSYjh
sxpRB/hN/W2kURhVpfK5iAmnz63OSk+sv2i+41MQEQd9prDy1S/OZqBlkEoXYcB1
bdNCwP7iffInyrk/jRu7d0pQQ01RptQWS3egMg+MU+JZ0S1abGeKOA92cxSSOylq
LAEPAi98/Y/R+5BtgAi9545MLTmgLO84shPFR8qc3hQzfZi+BRWbXCU9svJCauUk
iiFxLMeJpEn75oa69XgcBsWCG7sYfSf7Ymj5HNRhTI0ixliVAEyoFDBtvswBCe5E
y9oVgjU1IGEXYpp33Do+mNVD90q+J6cTfofXy7TiBqa1s36mZHMkQ78Ba0PfxA6U
2h31FIRbb99Wor7vr5khS0+PeI1bx7ZN9PoVhyqTIDa3v16q6F6mqI9JgZP1gTyR
OA/Pw9OHNfYHzrkw8BBHkHLxfNPwnLADweABoieeFZlZnjYKre4v0Siw254VwI+b
y4r2mk3nY7Cn3Kc2m3myW9+30vwYQRbNEO1HzQ+ePbaGnd3XVFPfZ+r7UB+Ti3Pz
yBDYIF/t5QcVRwTsoSLbiNmMarfVtLdrjrQkIQ3lAYnoFF5xwAIJeB++0wEzNpj3
9zrqvfx8d6ocU0ncnkwq4sprKrLoFaKNf1JzL1AtkhOhKrDkCKv1+yiVzOrhGp1j
4ohNPxbCEL5Fw4Uy8cJvyMpuAqVLYnwxBMto4dPHIRa8jY7omLHoxzVMYf9Js5DH
KZpi9roDCRg0E3TaOKFyOURWlMa5CtHdBWuvU1zXsraqGmdRpU5BlUdYD2NEMrHW
fF2udOgYra1BNKt1NU3iQcNg/Q5iKWn+5zkS7Uumg1GKwIVJI0C5ESWi9ekS6fja
dwYJbct/UO+oiXrWsWG4yqgkq/WnlrF3DWAyS+cYGJthkHzpOWHlkJSesptYdAep
T6nWW027mP9Q/MC4JNlWlh1HAZLtQPUTpeogI33s1WDjCnWz1SuJrCijwrJYjsNZ
uhj02F2uzSp0xgumO8EBLari7O3Hdm35gY1J5TPnipnwqzomi4lh8dfeM/Xyffve
LZ98K27PuPrVDfc4YXNaJZWHQzqojo9VO+/HRfeEAsR9cYOvYyJHWkFMabAP27ct
9o66kFfEomo/IQ2er+/kFR99wMEOEhxUVOaJmaHC4opSZ+tbFeJfqSpiRIQFf6tG
HHsZfcbDCXunD4Dri7ja5z7Rleak9GtXLrVjJqdfnM6ImuEiz2oRyp583iU4Xa8n
ihCyLJjabxbJc1DPXKOFqi8FvHww+HGoMzUvamvqZUIwn57b7b9iTI4MUgjpcO3N
g1FI8CFQE8ydZelIsoNdSF/S7VBM2JrU9lBQZwToFa6T3jOaG1Xfimx9HFURg3oA
Ci4S898rlPtAH/4f0u2qI8dJbf6JiH+p4fvlyUqma1KGIP7W1cxsItJXFziup8+l
GWDohaJB7qDehgbaqx1oQG9dTXb2+hPB6z+tCAD7a5Z9xFYAbpAj4Tgituw/TVK5
Suy6wPt1itI/7SB5b398xtx+XFTjGKBWh8N+WJ2kt2GabSoacy8q3vEWqdYE3hMh
cb+AGlN/DNtpsUaBq6TivPiqZ4tDXPm4ZZ7zoVHsEft9hYpzOQXXVBlozGe1uAbV
7MBUKexMpD++Bp2iEXg26mFtwzoIWkdvFywKO0wf1Fvy14QakX9obB3esD5H7G2S
k8rcif2H6BjWqESZQYkrXQeZKUKDk13HY9AEy+ZqkEWfavWmhYkLct93q6bIV4UE
UAGmRH3j7fZsw4/YWdJmEZD/1y3kkvh04LroSC1BqeiX+JCwH0h8rFNR47+elRAx
ctu7eXgkk1fa0wUBsDGujXxYxLrVenclnC2vjcyII8szY/p4mNo6H9otXGigVCrp
TPkUcFTTwt6t4bitI+TLhRStDlfl+rkySF/grMILRauzQhT8n+GSA0YI0NanNj0i
9sphHYi+dKSeTdDeO2hIbEHPrVPpBX8Kpdxgi0krp5dJu1+WGBa6LYh7WAUBBAXm
vN+VHvjqnq/kL3p9AMpqxjA8kGi6HLSI9kpTTQO4czZ3v/QA+q8FFQkyN1Pb9WN2
QRptPN0VUTqtdImlx1Gm3i2XhApN2qveyWlY9M+XYULt76Gbb2cs8ovf3C7BG7St
WzGn/jALHBg+KlwpHED+3Pf3vUZ2FF1VB3n6+Q25XZTIbC2KuvMZzH9TrVRsOQUy
soL19OD0LwFTjIRgUoId+nCAyvyFG8Pl0cVHzOjAPds6yt7YqPAWUhd4oBO36Kln
UykLQU59M1BdVlP80Kg7YFEnzgpAJjIbUR2oJw9gJ5fWo5y8PsEDivSYDqKE2gRP
fmAqY8JVF9dRpZAFFPvwvcPdH30T2qM47EhMw0nGAV7iCZTcn6JJZb+6eEfu8azO
+aBC3Xopumo/xeCmOIf7MCumGCnhxnBitgawXeXC1iy2yMnGytygruhE9Vz7dCng
PGGs2D5CRMVnXgjagSaqDDwHiGZ6wfflUjN9smgOyL19Pjk0pmLq0X5lYhD1W+r7
3nAzQS6rU0h6yIKMgdFGuuwAN5K77Ba748hQnejDb2M+PGyOkZ0ZOXOsjgMKeXfu
86Sf7CtPybQuAO6JmBi6RrDnWeuvsNvR2SH5XVfqHktgFanl71reLMozdoHLABTg
GCNpQvzB/roH9O3uUHCo49lDGdNZft+2CbULBAMdGNQYr/fhWXTA4+jV17c2ELgf
TsWwavq4kTZXX6qxdz4+m68jq5I2u+L4387USu4tX3yl04p0K3m4fS4P6eyo/MKb
OEj8hc2lWYK/cxL/TgT+IfI8fpK9eFIo9jRxgmJnhVzvhbcOlmffDIY+GJfeKbm/
gSuhjvHnMHASHVCJbm0HmghtFbxbwnVVadLGGg7DA/w0WURt4BuVBuIMCCwL2Crg
DxWfMtvQfdQNWlW1FVJh0cMx5ETNYvFqQnf5OKDf4ThnAnDilX+21UOktcq71+Nz
Atq4UVb1K+1lf1skUfjZqBO4s59HKm+BdixHch7YqmZpIAsAyOLW4/E4O2MNa+J9
CZsT7TGlWv1vP5qLz55TiVcGnQVJZmH/tZLXEZ/jgjOX+RJalV2+J4dQk8cCHoT1
qC5j/Vo5jdySWdjrGm6jBl2rC/Hr3hxKTp7XHLYQtVs/WUXdhSWUGl5sBGsd6cYA
BOFieLrGwrh15c8Il3kRlqtIab8WRYuu7BBDHnOX4edJbLWdXEDk1zBC9DKHlDr3
F4VZ4azuIDqGjR2mP+ouqZJgSRIoo1tOt4erGiWThvr//lDSuA1e2ncaGdh/I2ec
0To+OwQI/SmQqfTj89y2VjU7LJPP068k8L6tpXaj/dlyTD92tC1wTBVxDZq9he9j
trNJGlz3JzDAterXeLKTtHP5aHZDFU1y6ix1ca2Qft7Ku3F0h/LkMqHdDRQT9ZRq
6CCrna+tZDg6hbiqGfq18HFq+fKIJlxT0tRjkAi/R2rcwcittouGZe+JHKwk5PWq
rtnr8maaS6ZJTTHJ7V0iQxo1P5h/J2RGSLJuSOhssbpzES/FffBE1dinaU78l3zk
zFDc3xj42Bmk3WSzLPk7GYMU54SKSKQwwdWtzBYOn0rEyxE0XgvoCdYN8QZaiDjV
SwdGYUuJz5uLayQyDsZ1jegHhKShq2K3Lp/KPaDJd44xk1yVIq2I3lAprvwDX24h
F6etPskeT61b1ZCrZeuYEB8Wp/SEqej6P7P551x6ySJVbTlzU9TRi4YOEmVkJL/x
wK12zSmzrtIv1ESkDlsaYiTWg/69DL12TFw8NjzziTIdbD/rteWTPg+gF7SjuUwT
TPwaKjbtZQ8qS3wHO+m/v4fJuLRS2n4XgCQp9zFdLfIKj50nirY81lFbiPDQ6jWc
fIxI9tbLSBSlROfZ4zhEG5oNycEHKVryeLpDVr/HxYrFOGhPg2TowIeqnqZnJ8Hc
hgerDeyV49DA5je6/kd3Y+/XNcHo4gNNm83ddEu02IOmEWBdRYJC/sLXBpZu3a7c
RilqQe06HxFkzHWOs00fUW+MwDdRQVX4uUeJbPpb67VL2CJNnYMcDxV5FMxYTsZM
+YKgqXPjrSRd6wrs2jlaQzu32jnxsZocR0NZPd5n/M6xJ1JvaHkdAAqLa4hPik5I
iA/0Kw0BbKim0H7CHZXXia8AnKkdKdMVkYkY3yaQEqinnFM9S/iWJyOH9FzukAr0
/P1m5SaODNa/t2eRfKxEf4ulvAelZ6ucN3SFA/fGHwLTI1KJ98YmkLbsPc4/hXK/
0ljn8a35F1U2B9+cS3QoMjUsAdxzuWuE2mNbQxvsdDPR23pDYGN7xbqQeKNNezu2
iiadLM5avWics48uk8XxgJJJDHHFgPbC/qu4ViNLKZRFZR99ksDKyXubLOOyD18C
d5gEIXAKvi1EvtD44obwC4G93pbuNi+4jS+434G/XChO8kltcPwEOypeWhj4gdee
viXPaprgBYubVzoiGF9mz8J44igsyTKjVDe+UI++Uo1Xe8FMMxwMFTmDyYxbcLes
t5OSu532evAT6IsAiWr0D6A+8PTJPK9znAyGHt6KcYYbz43C5JtRuIBYcOgn5F8H
1TSQDtnjX8LnCJXzev3ZCImJNTROH7Iz3ktzNZridqd3loib5+VkeCobX63rpVgG
jNkOCIPGBVaexValczjvZ0opvN3Ylwq3Gyh3WUQBl9VkyulHcla6PTx4XuvH3NlW
lDZMkqD9HJLTfmdWgDH/tiJ7bo5Cr3ifhU3mkeLaYcuDgjEhW50rCcAVjoJCk6JL
td5WAio/iKTh92qd5nKYyEf0qEnOXCjZRtygjdC6goEgX8hctyP/kctt93FQUGBs
oI0FXxE/P6xlk6/x89Y+2TfxM8jnX1a8jM/PkVtAMClWixduv/90jAO9/5YBFnAx
nNOB2eOuuJNg4v16p7tpX+qZv/XsL8CBGtWBcqtTxtdSMSdVZhfQgD2TfGQEmbCN
IkNC1KozYaJ8FR0pfAn2fqSwfUSt1kgarEgJHeuSPuO3Bz2mNH1vgF7I8QPrASP3
Y2DkhNZetbo7wMZI6g4dRTt+Z1qYXlVDMNGBoihqlxjdA2MV/fsc39RJfKz+B9yn
pkQjF33PB7viCz4vEM69ZSKH4Dsm4kqrkswQvu+N7pxTZEKkynNIHsnikEN85M2I
8IQsSWRT7WLrX9iOadSttQToYo1/LqM994YrefXoQMmUmE2zYMG8iLvTHUZl49k7
6LRCAJAEk/vLQDUPLxbH8rucmlRwxPkzYSC++opzpoiZhU98+dMiPYPo/mpl8fVY
SfF38Qa+9eG9v36qWMevobxrmWH45W4i+yIQTKZ1RNmIiXSz1lLUPIZWIRxIqT5P
RF9zLD+kgy2BTfYaviMQ8oAeKDSowucuuvW4TFiV0bawkWih9hW58Bg+4KgRcsBu
0oXY7ue4uWgOWyXbjv8yN1vEtk1UIkxeuOIe9fp9UCmfrFRJsLi4ugTe+3T0es4w
Kh+6ABHihmdjj49NT4qnuCSfloUJHhIpBDxI+pDO3V6dYp4iUKMdgYtGyO2wwLAs
3eWIfedOPQMYdJG/JKTuOBYS7bCn7e/Zqgg51j8CjKIicb272XzCIIcdGo/51m84
K7aw+PQ11u4M6fRKJfD6OhpxxjxvNhQXnsJi/5/5fXPeNmsYMx77Al2XO2MQWTWv
IEL92j3flQRXqoZ4k38g6r/ZaMtXVV9DBOJldm1i6FjV+Ba5HQW1nOtTO6Agt1e1
YQr3+wFiW7Hw0oBvOKgtJFBESRkNVPRvxsSQq8wSQvg4fflSe8myeEqgccE2+11s
OLIkY7PChLUh5MxzhxfPVmksuezRZUI772kDx76yFCZ8RiPOJ9lykz87OSiE6Nsl
TvtX/rU9xBKcd/VxQA/5qUHB8COadqksELOjoWhQ0ZBmZbcffNG6rsX7O1yA9eLx
f/EC9mKRRK+N4M69elbhEA0JHPTgBX/EbdgKgtaH5hMryjp6bwRJcaIqHG91xBx4
JZv/ZmGVM7TFiGLpgDH4+rvG4mOOSeAl5pQi1K9Z74Kaz2qUIsxOXl8SYFZcFv9u
vikuYQPxh/ZWL6tWJtLuwAy3Uxa8sBCDUm1NIjZ6c0aOweJZL6LR8rtF0vfhMzwO
s+HXGYA/WT8QF4DDQ31PnHwR6d5KiqcwwmQZXh5C3thtOBwAifMsloF4xyhdSxW4
e4fF4C2QLJujWAb1ALGKDZsbBVOwuO6QqTTHX9JMynHKrMvM+umUfM/P42GG2BFY
dCidkkBw9LSLW6lLV7xxwxjZy+ybPOF0+I+R5MTKy0iGJ/UKrxwgOCiGsvu4Geh4
S4WPLS7CQDlErbAYHldqcJApPhKlL+QcVZnucLAP5jUAGnAHsiJqdntvIdlyzG/K
J24bRFmQFTAQ2djes/E9hLmvq9XhZ3rBPayG+kX6WLARphGhNjj8apYXMWyD92yG
ni7NHfYmafazlzk6oR8WLZeLkHFWNJPBdxGlU05HH9Ng/NYkX/5Pwp5OfeYhiKuV
WIMYpGtvEihsVns3Cd/HQOVnUqf9WTMiw5PYjnJE55HjAmK1xlT64OFW6NXFffDL
cmkHOTdiaRo697c9gTgEPFBbNjDz5bxomayAJ5I53jxDUN1q/ONolpc+QA9NZYmN
EIe/Afp769nd1kAc6bBFHNgOUP03UzKjIRQnUnfdaq4b+Xke178DdszfVjgPzPhQ
2f9tSqbkFA5+1eyn7QkOwAOoSg6T9qELWaSwmjVe9iWpMw1+Zv9XV4z4sXzywLpY
E1lzQLEQ7dOP3EmqlFbhMpKTvCpQyoHi+4Tn8ywthG5qR1fz2JyPJNVnkEJG91w0
aIh7x6Avokkc5jrX85M3b/AlXbEm/ap3SC8vp6o97p9TldYEc5Uvp88vJPUcWouA
sQd/7EwScpCJdXnaFp9h80tuzeCtHO14/dxG3VYKr8X28rRqsDmOj3eFcjtAz172
hf3yNru681T/5NjZAje/9dDzl0HwLYCEjt9y47/og8jOwGoA5fQa6OFGtTUaRzXj
I7lF89kFUc/U8KZ5r37DHhD09CGl0f7Fj5N2IBGBbmNFHusoZh5R6y71uWoCEEC+
uzaoswazmPr8/GIrFrMCliKQHyQSSVFz9cliTe7WsolTaSk+Db2Ta6uvMhllv0Mm
Y6hvBfGXaWWgVgTSmURpmVdPuwabGt6Ff2j8aV6jLrRyyPR8/59MYDZVMAZCIxY9
t7lmyZ9gCcLBLjVONXub4sR3lOUXhLLhUJE2o9HlQPJ0c2on4LXxTKIa33nrwowz
h4rHBz9+wSLZLK5ifRWYYDfJOKPGCOM6YMVz320pTEfjhdzQPvTY8hohuTK34SMz
h83gbPCoklXYE11R1rwz/ggKroqLTPnOhO9aQHsu7YIKf9+OKso6oTPzReNU5bnH
E1SynadhdTiOJms39UBg6xs7QJ9Yt2V0FqQD2n1sxhm6wrYTnRSqHz9IpxpqOzTl
XuIhq3OD3rZCiT+2qCQojsfAwauWgbLyeFfGeWRtU1TAXA8zEf+AUTy9Zj6gfSq2
4xlAVcUl1fBr2pMT3p5j7ZxM10JkR9fOq8t2RxihDc4cZ/BZjMBVtUwY+RRS3xOs
FiioSnkQvraptxhNAdbppvr5wDK5BEUJjNQrFlrt2UkDQbNzHKmmyR4YdNi3VSIP
ObQ+LSvpgkTlG6+mpDAw5gOxoTvuyIGcCVWPkW6Xe+KYo3jzbeqplEFJrM2Dj7JA
nM+rxfpwXxhM8MVKM3ayXEot6/FjjRftTq7/e50VsKAWLM1VXhezD+OIhY1Ge3sm
/5QlSQ5aPDmsXBQ+ZeBc8UhqjQsv5oW2oXttVlDJIohq1IFvnI40sLEvfvAtztl6
pCIZA53Ejwt4Fv4I3ASayTWgrupRi4WIhWPAE5lS1gOi99ZEBj3AVgNUfGvcXL20
8z9olB/SKOghUmLg9qBl9QwVcO4pbUjqTNE96z9NWdcZi1llhA/tyx9lqv5Q1+gl
7YZTj+SUKVVDDIXe7IuFm46LAG2dlekSzB+cE5BENw9fQPXKyj70AvwQKoSYJmWD
fYnbuJpsDs7CsHJt/6ZTVFok3LQv6yPe1bBA15CVL11P40zqDWs/Z7ZNgn4FRIi+
1Y1ORmNgl7Bb8c34qgbUxpbRy8iIptmjR56GNZkUNRij8eTodfkRYkOytHPED3j0
fTidgjFZW7n8GiCWPXU8ZkKbArbwM0r5oZIo1Ukb3OHxemwfYSe2XJd4fc1wt7kb
WbtCYqiuJM13E3Wh9/b905pylPLYTtlW0QGam2IE4mW85dVFOtP/SvJznB1VH7qO
7sVSOxRTPTTysLLAFx3Gpdv81jcqw3bleFNrHbDWmBDUKU6BaAdY6rt20b/Tx2YV
N9R+KeVe8iqKNue3PNeryTYRa/NJWFAZwiCn0Wy6IVmuQSMqzk8pXKW1Pv2KFNMe
H3EcVuDehIfwzflG0CWqx1n8PFTFryhY6lvWdNSEHxFUvG6GMQe2roxO9TOvt3B9
MxSd7ypaitbFnZfLZC2tUiRC55u1zvNH2YTaXtlqchmLancyWYnSCG3mM0T9I0BL
ZfQnPBwuWIXWnwvBp2b+2k+hkfD9+DJfVLiBXWJp4Bs6S0pwZMrsROby7gtafwOn
gI5KzDNWXNYJCXZ+A7h3x21+tNuBfnMHxMRiibZAT7cw2MHJet74zSuOG6HOB7Dg
1YcWvXpBlHEEF4rsnEnNZ6fr27Lti9UMIeUngJ8xhFh//e9SXIWGsM+rb/bwBzpW
8zA8sNNoyjoLdeAJFZJ7VAXtHSH13+JO9eC2/+IgqORWYboORMACxeyuDqD/EyeD
9X88VxJWsvBCyLno1VrZmLzqgk32myMNVdTJkIaA2KE4Wb57BmO2Pr1dIJVTNo+Z
EyeeG7fYXH+4IF3O7ayfXi1PXdsL/IKPC2sHy+G5k74eHB9EbHFt1WcZtgWmOZRO
TX6uke/EG3ODB6Wn//xxK0YLVZ5WQOLMJLgSXJZZnqxFk08uXgZtzcWsg666HFQP
1EPBnDS93luz6sRiKYliKy1lyBFFDYJl0gU5GoTpgb5HQdC4+yO/Vb4dTDpbtAl4
mJl1y6/MjwhtBUyg2SeF5TRILOF2rRRXb8236MTVb4C/7brN79YrhGiH/4r8Xuqn
42sSnykAp3BkhNxhDgb1AlDIjnrCZpP7+q1p7Hkrjr8Yw6W/jo3mKIQe+26Wj1Sf
2tfAarTRNcgFQRModnyqnnTvecdQq343PxshysReIdylNZSPEG/A/fp2p+zF7jfa
0rQ0dvfTP7KpkJtxIAffaL9zukvDdKe4Wd5AEGo1SYyfJrRXrkeenbApVZ91AIq1
oRvPkxVzSEERKRb3QhtGUctKDvMrDvPCVPSFUb1jTF624zFnAsCgGBxKX68d1rSx
4rvlg0dedoW/9WtUfFPuQJsjaU0PLi9TqUkAVhaKXQpsk2SRb8j7KPOdz24Kc1zz
Tl/B5M4P6wnjPCjolomVgaPDiuOVniN+28NlTLVEBxGksKyBZVHc/45ofMxAv14Z
+5ImR3DS+Ex4nR9630otYdTBey//CaX26o4CW66pZ8jgV2/aEBnwquHAWuiSWYbT
i/7G0tlLGNvUIqPHkkymN3PIznONmxe+2qm1E9BcNnwRci1VdaFOxs0zw4DxHbz7
24M6FIHIG7nhDpQLJDHUaTEZEX4iMoLW1uD31jg/f5RrdpDPPOmhl93SK9HsDKn/
YKwGzLuxETjVchrFKtS1e7wKX3nMBnl9yn5pZ5Tce6uJ9RjYvSYKQk7KGzn04rMt
R/Sr4gUuA8Q69AzbvbMBxGZ2WBpBp9YeD4VpkoSsZg/+eQmLXHLM8246J3LqaEO9
l6u7AZB1OwmWrUuMGxNrZt45WwDA/hY0fajHPlw9hGZckQNU7IyvKxkHNzdHX40O
RHFyuuRjKok0GEiM11nJ4oLiDjGBkMMvchbvIV59nNM3Owk511XzuaaxjLAORyqx
mA35jcmtdh8RWgst8Q0JaL78eabZoATZ4FRoe1SeqfcPC9D8kUy1W+ctg7GTEYnr
ix6o6rkJ+e6wjn0HF/jQiMHxMO6VyysrDgiyAuNbNUdh8WHrMJ7VzUS4dLlk1olW
G0F8fdVtl3lgmsFgLwGvjKd6lsrXIxRI94TBZ8rn6/sc1yXgXM3/m016smHQzlRG
xb2JobHDV418mzo9KwEy1gvuxrX6iri/Gu8kpOBI+jMQHDFMDT6M5oeqnP1bkd1J
e/R4+A/jC5q/keUNUxYE1toGKFdiJniAP8bOCH4OqyFzNYz6KjblEekqWRMIbZ+O
sii5XWuHWWSpDt74unZklj6UFOCzs39RtW17Ot/Vgwup2unkJl1L8zT4LBoyUExs
GgcQ1WbAbLicVRHUiUBAJFv89ykAFk+oR1iblK1TUhcID1wcl2bXhRKf47Fv3y57
af5qd9lYVOH2nFyExKLfRDIMZ9DWD9a3r6Dz1iyDGawTduVhtQszWKP8iUlM0+up
XMiQ0zN5fhyytZa+L2S47j91GzYfaQrZQMrf1xSmlPIsIdSKNJJ1qQI7dFTbJhBG
ZmDaEIM+B+USpxpPTLsBxWHf6otF4jvYtKo8B3WB8YB2VL+ypBvLd/2wTZzCG7PV
oZTtLRdOMjFUyMTHzRYPlrmPi8cvVCsDCnHFH19am2RYUYNxFYpXTuuogLU1fS/4
5aBfZrciqvSPxxBWMu980dj51twIzKyQg0zIGzUmfZOyakUQjS2NID71CIQo9YFB
eOJe+ISG16v3fzlE7WNIDWrNpNetD6KTvaDvDQ+IGwdECA+DZ3bdNZ3SblorlQlC
ZXskeOkdl9nf6gkvMFHphJqZCq/lbq7NlWcdbvC5itMyesdYHpLb1Mo1l4sy84O4
01CwAXTJ2ynyTb08kpfXgWySxeQsQYcxdHnKli5TpiHVfKF4+GF8X19Dkt6TNeB2
0lrgwGtORcMrNAFkNGDEDaeSfuf1aGpoUJlxNAzm35jOR7IPeeQWSVXfwJQXjVCR
3n/4pQ+eI6Wwh22FgfYUTNRpxT8hvzstD7Ik7469DZAsOGBQOr2EGB2DkW2L6o3d
GR7sDbtU4TTroEwiU78S58bwtZpM0VS3kGDKwCQ8pMgn+9DUOYeDoZLaiYyNo8GO
q+SWsFYmHlbvqgtz4hNOBhrRP4BgY+n2LpGZ0ZoF6kZfvjL4k26FyKdT2tfdZbnX
zymh3vEa8779WrkhqXza9MIfgybvhLWDsY/uiT3l2G5sH+k95DoEOJJ/Nq9VwDwi
PFVfdrcS9Lec7xyLzwNFPh/RJG+P3MyaJDu0fUvNA26RSq5HJ/Zk6QB2OCusCYCL
mffGjKKXErqTYoGQjjKvn0qjQ2a52946j0jhnVHOxsdxoHU4uqaxJQHgPfAuXpa9
o4dOCvza9Tjt7ljCPOl2al7/wPuov1pJQmDPMw5ik2Iunrbw+kCZSWYOwH3MLZsA
QVoNkahNFGAfwnr8D4Zq9ad1If7nkKYxei+gvwYo7v2haIUC0xxO7CerPuB5WuVX
3uW2hsRwBNROSNim23dNdpbRR0PUp+JrxVs/je2iQkSQgEXVAGLX+iJ5m03/U+x0
1wtf0SGpMrlAATmSz3+Dq5LAtEHf5Kl+W1uxzLQCqBpo3Cx9GrVRrJGtgIPK+ly+
kux3BOaJRDTkgN+ikgwDHNfhTP9BXfmfoMYEPmqwzwDHXUwarrLrn823cgceEsVY
xcQeDABgkIISaxA94E+V8CcGDH08NBKbI6XuoyFLr9FX2Q0gPdeuXAhhn2btiuL/
TIaNj2qq9GESMbKGsPcEAGOrvvPV4YOEkcd/VwfO5zW1Vw8E2pOkNpWoEgixcC0Y
3n5bcJcouglr3Mp4vSHfW1QHpa2ADq5uP1xz3Jnb27ttH7iDNbQHcEEbOXxrylgy
K6uh8N/T8h+B+47NRrd5OxWa5mdJvSbJqaBdmsMLE0C9bb+aDOrYVCJoGrsW+aV/
0Oa6h2PltjcwI23TJrpCyiWr5fg63f0clFujlD2rc+vQgLywNAOW3rXg/Ut0VtFy
VY4Yca0HFQ00PwTmWlrzacw5+1/BE0b+xjdfNvJumYEwKG4yHZD3YaXzGU6DZFC3
og8Y6EdpH9gMdtG1feezJPc6uJvFOBBqlqW+qycj3wjogdaT+Qnw9HFGiTGC00f1
jl4d9p2Oghnv5hSL4iFOrgGCm01ojQrPPYz2/gErra1vm8MZfyGZTw5MXW7dNVh3
XCqyIAcX9f0nGsOrRow7udxwMwKONBkEkHmRus75rQ8zCJHIdKgjXHKqRDlhDM8d
EVjS4g15d5hB5Zpqqg0LZLTiHZLA4SY/F3WD7jhH4hxIFK4SENhGPmHeL6YkL1Pd
TPh12UbacMZQm7NWg4H6bYZVRz+fAYxdE97j69CA1OK0r7FYbBuDo0bhgIdYuJRj
EqsuWMipbU8XXQ94uF/ifvOVUFIaBueMscKQ1neb3pNItp3oj7jUMqJ52mOsZlXm
6tuhFjMpc1I4Td8t/sHHsnedseunJXnWJm7yXc44vWfKgwROo27N/Cjt7w58w+9D
paQUgsAiLi331aI0fHIjPIlAg9MRrRLjtzLa97fRQvRCyGb98diy8N67XA4BTi8L
vrkf27ycaFP48N+5fYtbo9MLiPM3jCAs870MomEA3gO4TCrds/2YQ20CRrvrUn9W
c+Zj8YyKQ5OrPQJOgBdDRTubTupxxNKrQ8NTA0yIuDFF5zzqKd6fYzQHU5zxXoHx
e9Qu98sw5zOG9II8Jb6bWpUUab4ofM8DBWTLOErfgINEaWIuQxteSQc8Ql5zuQnE
rryu2Tx4SnFnwtT//Lft8qTvrzkBktH3IIfrsqsHVE82FJkVHSv8BUXjjbjHebU1
H9a083L1vkhoGF0E2pmjVzlxGvrCC1k4JJToA3Hu+lLI24EGgAKTkI4taLhNQ2Af
yxnhGc57tKM+y9tUfkZSImhQbkRSD6GVFKezpvg6s6YlW4+5eIv5BFGyvyl8pPUZ
K+VaIPq2E+Z0X8o31UCWpFrt8MDmz6u2V1akSefet+mivrwj0vnV/ZEXWWqhYZQc
qlCvMNbU+i7s6/kKyzEwvtje5MPw1SuoiJM6gWw/PXwMgeLhRygl8XEGA2ScLL7V
KDh39haxvPra1uNFrkh3sjTsIm02xb4bD+wzpUcrFYxqzebZepNpfrhsddnJarw0
pDxpHz0HONZzFvQQI+lc8n8c96rST0qOl4bXhRL97e3vLg+RlWNK5/zVej9hwsrx
8gsU7Cj9k7WRgjfTuKk1XWON7yUZFOlYWD1AMIOIT7JQY7HajQRMp1DvXvUR10WL
ZSu/CIC5Nrg5uQkTFBJ5MP5LANq5cijlPXTI4HOxz4dCZWqnkORxhpQW2iLUDtVq
GBcdn6aCcPDR+sM5qDKev/JAg97bMWxq+GjGGgyPitSV9w8D13c/HlsGJRqV+i+w
xQwnAmZLipvMlD5agMyeSrNUQ4UdmJUXE6boFD9kTH3+9A5LjI+XaIB9SjJE4wgH
b+zOAuZnMmdjzJCyIeCN2xYHrGdpb0qQI1sn9puN0dPACxE1DEh5JUPnulpBIhZK
WjINyrai/i5J2xc/EoFxg8eJfaoRMzr7/IyHJEg6zIeWbyOXjDJXE8OBPsJ3Ed/d
Wth/jZZKUcfw1hRqwq86JToZ+WzF1yePGYwmnfKAk+a5zvoakstNfXQuIM9XdnWE
h8KvBMVg0ygDYWTfdH/O+o94fU410XNERohVn/8G17g6mSkM5/PbT/Jslr8AZEHO
32ZSqfuXwKkB3POZuJkE1cm1A4Y0fZ2yTHIKMu/1cx8T3dFPu8WspNgNlKkKcHdi
9orWa1+xCKYj604ntD0XSSZrzOqVWiWwxfpMY5MBf1m976r7E81a/Ht9ME8fLjyy
IOrYuYk0lv8KYK9H6vM9/RaOq9VqCGUehbseL76d/xJ2p3eUyKt1F5ZmwTSSysgr
1Z5U50d+yK6r0IorHVNToEVWWUhyk29lwVlhQ5Wku+3fKYf5WM+V//JawoIrfJso
dSwyU7+2Xx+HzHMs5jQDsiaf45aZaB8clHeoObMU3f71KGWf5khsn+wBI9WjDVfm
1ZkqZ2K1Oc0OBW5z8OSgewvpchQMpJ61XgqCeW52r6x/LaaZ7GEw6z2XusZlSGn4
V1Ly4ORrjhAK1O0rO8niWlQ1C0XUzBtR4ZBnGVfMLcryhXRD0SYoL6w97U4Hm137
XQvwfb3r845ZkJ+IsYFuOaj/jFSUdbo2FQlHv+58WzT6FgHbVmNHPOYmYO9Yrf7q
XZxIsa2Y23V+DdfANft3ynu2BpZHuHbLO9LdVmBBWhZOBOl4dL39cZ3q+HtJeHHz
OUEGGPXr8LeEsYiRcxqIzSffuUxvM7A4/beLgD1otIb577qw5re5fMJWyGRc19Yz
QJOyRU/JBw+N1ykC2nPb3LWQXPT+cEoCqKpyBEiFZc2eQ/U664Nvx/NapD3k0W1Q
dlPoPdaOrna+A4XMy6jESJoAdmVACy5WRLUAXcljGSPPy3mMBPgHyYCAny2E+lUD
zK0XWDuGjGjEBN519umPRRwgh/cBYgNoF+mn8QQWmpRHJWvapcKAmV5xiChvhn17
uwXSN3sdmdxDBo81KbS2OJjba+JpIdZ8v5LXk/nuWknGAMOnIHHGDR8Tb9icumZV
6y1GLSM3dl21dcP6umJr8Tv90AAivL7x0cozwNCk5ERL93QgO+tj0qEGCbqNxOUG
DZtd8P+UjB+GtiOPSqV468TPJr9j6FB5RY14q+TcpF0hNSQNNZO2fV72STfTrGs3
/hmEwL3fXuidjPp8xhFYtxUpuxauz1+RD2jWjiIOylFa69/2SQ+QX9TRpMSkkcxI
8h/LA1yZvi8I8NT5gA83I4wBKLfn3bGFI86Lcnp9nyOgZa7Hcoko/UWM9rvKCl9J
tzcZr9Yzv8BT+KwhIjpLD/fwcIf5041nDwo7q/TlNfNBxFZu3eThFtv9lVL77vix
mwDZ1AoHEEnF4bU8/EIt9F8EeXwAGajFyFxcjWMY8B7NOovz0ku1zsMfnFS06tDm
DBT8Nwzb/cKJV86BHDwiB9mz39wIwPodAQuOrhtQQpMgputyVRobceARYatGs/4a
h457OF/Cl+eF6c+JOLBSd1DpYWPq5FrPuU8S6ehYONEHSl/KlKc4bLfoZ8GfLro2
fWLe7u+k+AgWP5qj1AwOvZyA54fUKfzAoQy9XQVF2+xC2QfKIKlIP92xeJyV9t88
tulo4vcUViaTJy3iHXL+OJq3sIL5i5LfNgxQOKoXq0rDhD94Z0aqRTOGUatXTJDi
MelQbcu2Viy14Q1ZNGNXUMl9oLNolE/aD5mNW1Zvdjew40gL1HpwESJbsKnN5r2g
N2ni/RIl4oighpCM7N7O4y58CKc3qitIeAseGOeKuiLbxVwTm70YjYpEFe+i6aEc
E4mdM+3YxEDTyVI3PZcR5O+vhMwRB3SML0EehdB9uHgQ6R+w43Elk4g6Z/fmqo4r
V+TEFicV1EuYwAMoY3vetRRXlUYsaEjquV/6sKYTokGa1Zx/b40s1ZbtXtdW5/gf
CF6U9O+zhTOMxWb+Ub200YQzyBPPw0Udi5RvLwwXLe82rcxTTvyOOQbnTSF7zs6o
s6GMPxKNGtr3Lmb9SapOoIneSV9Vw4sAmClnEQWIoeUvmG6fmUFkv+/g9Ww277HL
l2t0iKttmwZ7Ew4i8b1uqLLZ8oJASVI9Uo1JO7K+EZWSWErz+gemRsrV57l+GNGe
54JVhcnb04da50L9tlCCBOzH74coes6w0fcIbFBfsqpxvjPh4KO2iy6tnpiTUYBc
8ITUbNAqWdNqr0BVBXVo0gQb8YGhGMCVRDqx2j1vhj+RnT5Oy5+jpcVpGzjukT3N
kUevcejMinzFfMl4JlKZci4/Lch/WDJa0un0hm4Cp4NjhRskyhuLCo12A3hjtJ2c
lMFKiu8/fxzayvyxJB1Wf2Zn3AYlW4D509cKaxIxZyrGSzSbhe41e6y/fZlbvMGS
R6hEkMlqjSZOv5gibSTC2iCHvJcn6PU/0rocVP5AYMF5tJOC3dTGe8aJLOwEcEYG
6RNh2G925hIUAb4qmgS3Yhsc20xRpSb208ClNBfMI0+3ftH1cxx7DzC8NlPMhzFe
to8VqkLABX3O6gDMMBc+3vPiffQqFAtMt5D6G8WaxggLsDkxSanPkGFLHH4JWUMB
n/SlGEv567B8//n2xyjCwhV6djm3Q36XaCNCZIn9EgASpZMEKCJsetttwx9Gcjdd
JhQepapfuj6wvJvcS8UMT+VzTKn4oIzxFVVLlcYx+ZwFIIV4HdyNn2nI8bdmSe6t
IwsM82PRwJe7ir0NX94991e4XPk1sxzCFcba806TgoS5hEtWm74zLZYn00M6gzkz
UJKyEMcJeQ+v8A+HEXKQC7v1gXbng60QE+tC3g8mSenXsfyPyFABOT6b8kliQrWK
CyV+V2m39mQyU62gnILFAXJXAovx6LuN69S/y+pqnxKhkHWB4Zlrrl/fMZNqeYZj
qx3YFG7jpDILhHRsygtcpj27wADPsY3YyoOfv78pRMovbYTtHC7jTl2x4svqGANi
j9+aEzlJSap3WDWAggDu7bYf+hypwZeHmMWS3YK9w7VjaOeh3s03h4AnGLjnYtPD
CNkBlVSmPZrHhhjRyS2wqOma6Hv91vZgpT6PSqPAjKeL5Z0kAR4d1X66qP0s5JBc
+jUhiKV3pXy3tQ8e1BGxkIrtob2BbPS6oS0hUeXeHPmz2zqwpfpsxMPaOCpmYHBu
5IjHyos5qt5ZuiYYPdtvkB3Cc5nLhaTW9pm8YWyzCiI2xgV/CKqZePeyNZx+vwtn
hhGXEOuWox3Ngu0d1RIZTdCAc6HgmxOqxoz6O5xm6s94KZhG7Jq+GEHySpdATgwd
JnDKQ10ge9ZTDg88s7AYTkv00G5BqdL8ItcwTfdO5+ISuJiGYxoFOprionpxkNdS
DN7KAL6ypcmKDH6+S2M4+z2JfVU63ClYH3s4tLAcP8zJ2FQg2tNTQNOO1iQfsucW
bSSQjFCyGjrvuE2VCG0SzXu96ktW7VVBpoDO3HNRnSGHcx0H8HSMGNCRbaAXY4w3
inLHTHnqUSZ8lK6GAEf9Zq3BrXNp7PXVlbaneQF4PiBHpA0qiUbUSfLzCT7xgOyg
F9IE1E15RfiXOPaozARX8BulI2gaaZu7UgagHc6K62RnsbBcDd6ZSbQ4rJOAuvJs
Qfw83+4IB+G+3PHMoX7FVfXcNKqdbR9WmXaXQ/k2DQzMuUxTBd7DDevPd48bd9gh
VaJGEuzToxHllrXiUUd6KNgnKvExu4QXy0KpFOL3nuz8ibZckgRYFXiGw2weHBvU
rQvYIJKRN18FdNnjHEkJMyG4V3K3vxL1/AoLhpsXcroZPYp/jFaGXnPgRWKnl53F
R/XtN8SOEiseTknfMByf+6jTRwfHwzRvu7OvIKEfcr4z0DuHSlYcYY4NIpDe4VGa
F35BxDBr0q74utm84roL5RZdr6kc334c5ZNFHmp2h1S2Pi5oH0BmkG8AIYwRy1at
xeOeAd15sKbyT8P8RpDDQU9Op5ZFsNWrunamjJgiNNs/X1rZCtGwLBLEifWlI18t
eFxYNlar7wNFbkcmpAgriksxNy1PKp0sx55eIf7jnGyot46dUi3f1LMh6bJJ4Msl
GcdWAFzcxzQrCuYrBD2XnMvYik7bVsvVKcZMBpO4Ywd04Dg/+DVc4Auu/5BEuCob
08wwleRm3qFmjF0pjd9raks/UxnKmJPvItXXXMeHbJnTNN958nf3J9SCFeBctxN8
5RQiqO895n7L87AdGmeiEWgJEVO/cynR9qLGF9uQRvpH6KhlBUBJJJRlgL1S6BGl
x1aFdAz3yRNTJwTkC/WdsWVtw2awvgcBRa4ZbvalbdS1q2oAWSzfE3RSbpHQyh7P
za44MmrbVUSKWfAtVWd6Jm6VfFK31py8gpDdQ1BU3aj2am2X3HJYbwo2qeBZgdyT
au0DxOtukH8h0EElbzAF/NESlkuiONRDAB8YKaJV/QFeko4INClCD+JwV7SxWGbx
SSHq5yHMKhRN0tQlgRPmbsPMH8DfL0iuurVc0mJMlhsbCCYAvPEGTTUt5DVz0KFI
BoyssZ6zfI4WsIglGbGkGuySRw72Zenp1T+GnUTByXgSuW0oltVNXfxe6ElEDt1p
3i82TIGUqF3nBVR8gFoNwP7Fi3/oIKtHuDyWH3Ovg8jzPRQGkRwQaZJRvEfOIsHK
rBVoQ8g/L8wqs29EHCu2/0xzHO1mLLhangGWhuZYzAVuclH7SdlA0RHpFJRnlJg2
mMaXveQHsIQbr9iBkCc4zeg2dEP2l5+ZyP9s3SHpPCgDZm9Jhiz6aKkjEVAQV7Zi
RVe4urjSCnWYxmWCzo5Gb3rHJRDf9H0uhqhn+KhzHm5oeW8b/ILmXAWiMGG4V7x+
GH4XCGv2TC5v+p3Uzy9Re2x9RGVDAc3oBMTQEyPOlMIWFe8MATV2kXayYeenz22l
T8hC6fcKGt/BfJXcHPVwQvPpPWdWFSHdS2VD3J58skoAqzCCVlVZKItz+zVSvoS9
MbtfgNx/9D83+Yq9fUJYC7jpai/YIGJc2kmi8gRQx2wTGWnS9cRVj2o+Ll8LXdUb
ZLSx5+W88qhM1VCtSf7V00/SsxYe2PpM2+REElFvD3kOwVw+TP2xIVSGxNmlFV2+
TVjiloXDXxhGR2LkTUxStwVHY1UmqQThvSPLA78dRQxrEdroEjSG2k50YnbTt2XF
bojfZ3ws1xgw7Bv64MrsAg4grsun7GgM0EO9cNUoGL0ThWlFAisSgH3mGJBiikZL
P0QyrSRdXx9EmuOMBDIUFgRjdZQCJD4IcR1o+aD0yASC1WkNAubp6ExyLOdezhwU
Ud40sGzM+FxdMP0lvOmF81UCH8EB+bo36jucPcpqyWYqJZpXNrO6jL275HZUOu1N
db8M2/KhOA44UlZ/C3jIz8qKqgKmVCPfopeVGeNQk2c0UeIfGdvndmOhdSOiLMC3
x8XfCHFgh3Qa+MTxjCw8baZfqiFRvkxuzsRZQX0XLXbdeAOR7HS65bl3Wbk0fD/7
qnm40mxbF/hDUz1nIXVVLZZ1dFq6cFXzD9NDRCC9IeTSpqKbfV2BHqJmFK26uCaQ
nG5QpB92MNHyQM66XitESxhb6Rtw4i3u5xZc4H2b+dObXbVXC3Nru4lyAw3+zkZH
Wf2HfhRhtKrNvdc04PiBQUgbqNHTSd+nfKZjSPhBzn8C+oLq9iAteyLi2DVgh1y3
FwhDNs++QXt5T8HtEyLXyz/JLNdQYSTwdORDgUWO213fQU0vGYQ/RMPMHSD2+T8v
mAD6ZBG/CgfTQ1jfpkEHS80QlOjsjFbSLHmJpSyQ83VTwcNtf7TYdzwEjL6U6hVp
N4bTWaxDuSZeJId+70bNwC37wBtRKqfG5QP+IoxpY7eRr9b0LKrPdLP8R2ElVkGS
EtbkghwegpNnV96tXwLGo0anJxKBc+dgJPkyBUNfxa1vcPiZWyDubakZaFZ/Q5PR
zuuBlg9Zq+hh3VosmfI1GuacmrGZY8Oip+DcqlUe7mEROQ+IRdB3M/ZtKkM8mej8
P9+R5rRPPdmjSxgDJwA/6HP1MmmOTbpE0HvW0bT24BKilld6826nzw6ZPveEtGxn
2wgCbjBelyKCJpZDaIFUCe0k8DLkPSEwcjGzVNukV6GIpBNIacjQqx+doI+y/mHU
CsreOipTfxWeLSWpblY0uwRFVFfKiJmgAaw4FF0SATbbUrxKaZSf/iRh/OknIdwD
fx1GIHARBFqQ581TMrXEbUHsbCo9OP+5h3w0nuWqIJ+QLT1J7fYdzJ9Yrcswnsz6
ZR/HXQmKPsvmfKMmzqXUi0EE+xXMnTHCokJN5zq5hQs4qqzX+hovReq6QcMolJzr
7BgOhGCQzVDhGfL7sbPfwOVKXzt4gRn5Ns7Fb+has37Is5D4s90hKLMllk7q2tgs
IZtUSuDotOjq+TZ+tC9yS5r2wt7a6cOeLdcsOHeena3/zxKVyPSl6rX41YY1qVWa
rg7ltYn3jLWGpagMDbXFE8nAU4Nin6A7dSvVst0zgJVg8GXPzSfIgg9x9gFa0fa3
N3b9AIXu1yHWRRkmjNpULzOjxbRWIwhozFPEw2uTV3YluQLAdtoGoorkysNMn/ur
fcBgI6fA3Qxeuyt7JVDnM74MlifmuN49mwk6FIvP4eWSupr5TnsNWBExhCgmYOoO
DixOFfqQGNYMXZm0eI9ooK55De/+oqHlhOtYjTwfJRv0tiVq8sInSVCFV7CzH49o
UIKV4s7MpJm5tbbi7jKP5vPTmR53aa/izxI9zCU1vJvUX20rT5TjSD/CnY1UNUXR
/Dd1ShU3KskV45ZXQ4hMi8m/ppQj/mmED/Sg9f8rqjgLmKjV/QNf24D6gpcvwmH4
6fjvTdI2u9+hzBHyeRsYvQJV2cxdYN/s7SzlNCumSqyD47bynZWZT/UF+y/qM1cT
03DWu/SOT7NyRICqyCM577o9bcmgijfWH9SUv83llkeZoUGjttYFtnwnAc1/9Xam
TxcjuTBbDKbhCkA/i35B305iDchItRzQwkF8pLkvNcO6Ze++g44WkIxsZxBu0snM
ugok8vcJiRnpIN4YdayIyAiIYRNPt1/xyFkmgv8sMEpvyxEIZayGAdjcb6miqlV4
L8g9zPDkp5IFC8MN4jWwyf0WCjcl6i7VDfBFtI1ptg0uAa7AGE4AWlcvRou60xDZ
617R6pr/MEpwFLM0nSyMth40s/zKgXQttwD/bzBEWcE74wbhjnHm7GjyIuPLeNQJ
9tyhBFSsaLJ9pejk/272N2f0oCOko0T/n8rDiTZgbwT68ribIdF2xk0KJtb4ecI9
6vBRInHMCVwZvSQoEmLQh71jZ0JVPDpcN9DMKXvQzALmTlreUuGaoHgA+sy2NOaj
CAgbkIoK+EkM1kjpqVuZuZsOVSdb9EKv/NZHuKEMAPTPsgez54pXXH20LozfoOnv
IVDI5F6ZzYLC+gVyTOjvN9W6FdIwKvlkQX0BG0aBUjQqIu2hHEk6yRviy1DlZSe5
KYxQr7GeHUvv1G8PYLGGqGgpxGkIWU86ZKjkvFoi6YZPzAJ3afypQhbmrgWJtgJs
YL1s3bLum9804n0ObNpD0bvpoLVb6/X5BmiBbhlyBR+iEq1YeJnUxSncBdkMoioc
LkQ88PIwjft0B2f/h2OUCGPLs3go8/ojXbYeDmBob/7lNA+V1Z2ehzl2sIxH96nI
znGAEOSJLVkLOfvNbvsPEAoVZZXLKKxzZwC6Cw267nm/yQVCHPm9/7delPq09KN4
vq/WdKUjpmRRQa8935Qe01fICTZ9aFDz3zW2bgUiCu1w/FynVltU++8Zdl5bYK8x
tVKb0K1MfhYYtOwR6zzFIMTFR+ZC0jf/j5qvctcOnSYnisbZ1UJ5k2GHDFUsWbrs
dauVojd/qgKtcV/vk7Hg/ZPD5jv/KPkuddtUfFgHozVg3QRHfqPAfY0IDO4bp9yH
JH6ZEG50aDQC0XgzYBkVlEY58z6iRzO7c40dU/K/2sZ4Fm3+z6Vkp3NBX5APx4+d
tGuDikQksAT2B4JPxGL2UAM4nYtntX+kB97eEY+6aKUaGBoukCWuEIq7YFo9dDUw
PFYuzKb1f6KiAxDI1sGier67LZdCllbrz8e9ss8dvMznzaFJkdU8L5phh4fu4lJS
tR6FtpYTVpelzfAXQ5coU/9+VrglZ9VCnL+7YGld8iMaRglDSxnztq1p9zZlrNkH
wVjdKN1hJaYsE1x3s9WRpsjM6chxGJChzOa8GElOXMzwVqK0rMaAoNFIyawjKIhp
bZwkqwRntwBfU1mLLubB1h/4+EqRvCPYNQz2AaCMuoCPh7JFLD1JySLoelcwByH9
os9AOp9cyDG5QW9NyVN7P6vh9LxcOws+MKEoj67bhKoFzVBFGBLXRXR1VmwIW0yH
3ibSGY3VkWJ6yy2RXdSl0BuRvq/V2tYzcYxymJUy66bTguiEGHIFiUtuur6I1kXw
CN7VNpqo2vbMj9rTgyGtHiryB7Wl10Xqy610amgOS4W9dPh87miRR7F3nS0YxYeE
ZCjQsMm6izUDEzLQ/2rkVS420G12taACMADrNLyOgoFx9IazzRgI1m/mEwHvwCCy
w4lS3uXnaSr92HBgW2ufsn7RBXQrOQLZMQVvyD0SScNuJZzqZfEoraPJpRe6tLs1
Ah5Uh58VKwvJQqljeztpwe5GFaIoQ3Mo584vNCt4jcSC3tmkBuiuC7xN8sqm8NrK
V7xKpO83wWMq72Qlduqkw82BGx5HETzwxy87qH6s0obKVq9UIHMGSiDkThRgay/I
OZHft5fkSGxde78OcliFDC25aqSJ3S0Uc3iXUiKVEgoTJpRP1UpBnBs3aohwKxgO
PAz3rYJmBppcnBA9VhdJr3sg+fd6hA0XtTWO5ggrV4QH5nm93+eba51ibAjHavq3
eL9xpRSmU9pTRQJl+KwSg600z5uYejGfdyY+QaEXFdIluMjqxguEvCeqpLRim9ze
+P/466NTOWpd8PVzi1Vhh6kyb++plydTn6c5/0VwSAqW420/b3Ambcj6UYiaiJBh
a7DSzZY3kcxJzgCgN9pTXElfpPftTo/28qSiCM6+M+Gjsl/fyDgX2RMB4KJln4yG
+TEEMnJqT7hI5czSkB+1SJS4zpRI6Ta0+licEmwHANkmwAiuAXk9UwBscAxftWwU
lHEB8d6VBKb+06iETXg2qoLTNC5niwg37CZ2I08gLEybzDbJ904192kVwPRYHvF2
Oe159rjzLgbO74o27laHZL9dyiC5n2LHudWm6906xYyqGK1TL/bsaxJzvXyv3gbW
KjvVmQ3NufRIVp8a7tRzfYoy16tmPLcE9OyjLK/PVVPAT4U9+fMrdn3ycgAYXsZe
bEE3Fu+5N7GtgOcokTCXloOQ0DYbyH3THFV5pRkoVHYrScthdtuS8EAgsZYZIwb+
B6ci0x8p6R3ExdsRoGhl0oGmdqgukpPscq0WKHCkN8f9sFlgLNy6frK6hlPkyvCn
TUcIOuer0PNkI+UzXSTka0iU4bsT8No4/wKfhCiJgdLKZoNdU//n3vu/5dgMwyK9
k8gWcHg9Zk9kxK7hJfdaLHPjUBqIJi5VVd9bsDGUGEwNDL6HjhEzL9YEap5NHfGp
8hZN08mPlxG+T6WcBUsboed7Dmz4u7zTS5CCkB/hEjULD0yeP8UvKIOufnWB7nP0
XSK+nONjfszG8wVCGCReq3VkW1GygJtah4TM3yTxSgfdyIndHxrgoJ2BQuewFgWQ
ArlZf6SopnYL6+fh01W56brutIplkjXc72oqLDyAkEvDUt29LKmvlSJ2OETMdxCD
Yd9r/vJJjfS0dnXliyvnoTeH8RQ94FV4WVLTu/mMHw8Lo9ESlo7Om9YK27/a8jvP
CIfHLXJCCf+NFB0ShJ5Z4po8kscgqha5SIMH0LjZBFMrvk5mnm70c1Q79rNG0jFR
sFsXdbNTo52IsZzqsAOe+XXbGSOfeCRQnbyQuMRVGMqL+gxzP3SXzAi/agkuqMD+
0yn+/DvbYMECHyLNFP/aswcKBCIvAIYTEjPbIclHRJoBRQ4Q1ykqIxD79sP1FZbv
zwtP0wnGHEF7wKUVEKlIn95poVPbQrTYr3iNHE+S9wYk33AJQG+nobfB7pz+y6HC
NO0okl8JI9QNRLf1uG8sX7Ir2GWmCQ+zOlSfj1yoS1/QDpl0mowFPnEGeCs5DGyW
5P4PcF383NjtoEORi5vxGorl3Tynw/4g2bB3EMdsiqaJLxOKsdI95H6UGuYncV0f
OXT4Tm6HR0E80xPK8JVZwo6wAuRDfFmFg7VqGKq+mTm9RRiFUzga6XMY3KaCGPTH
D8nd9bSHQI/j3jYHlcmXJYGhCwQAqXXTIcAg54UBS4bi/3Z9jwl65fsFxFuRLBZf
YytcNEkoDxGj+11HIlL5YXU+laU2egE3K9vw9HWsD6r8f/xCxn/PCkowacJhxQEc
U4JxnmQJvhLhVqlx5Q5HLewA7s5x6PluNrznKSGCMrCkknlCkB9aQJXxjOnBhXuK
KKe6Y3FDQpecMwKWcmBlI1i2L2C2rldu93Gd79/qRH4TfVV30ebV4SbOzQeFfh13
eag5OSep2TEL4/mTfvLPJVsV8itEdexpIT99a4h6c6Uz9RiVyZJvF1JlNYJSunRg
isu5JIaw2htthbopQLpEhtF5ETgOOTw+uNzhwImkv/niMW9tZUt65Jx61T1olYrx
nxkeGoT4vD9mA+g/fWWhOBFsjkcTXnGZDFa+S8PlbeGo5yR8HqT6HyOEyCn1TlWm
+0sy0zaqWI3Hvay/id/qXOnhp8igrusQRLJinkrdg6pzaTUSsVGtvx4/+1HxVPhi
W6Rcn3T7d3Ajfhc3C3alc5BAz5a3RKk9LDVMuzGoJl85IIZ/8gWD3vd/uuzOElX8
k8t6M6jRqRjaB1w/l0RwwcFT81yBbVsKiG2Uj9YMtRF0lowmxFULZt6mbL8fekSK
Zcg33lbypk9dxn1RoUp5XL4Om0SETaFIQbc5MGvRaqk/igAKPOlVRXF8Tyk+bwJE
+sEF8eRCNhjJiDHRpmGLJE18Kb+1azY4J8ACsuk7u3WNZy++DY3jvBEw/4Euqrnm
XDZUJLI1shGHU+hMHQJXlmJp9h/7ByHWmb/0emfyjk9keLY7dtfsyItkLl0mKZ4T
dllAMeMeHz6+biHdXSJyJ1GkPb2BUIHAaSWwfhI985z+/YFN4jXjfptcif8vcqDy
uCuMZNY7Slki1jNazLE0mjBiAfahAX0RwmSQGv2u1hY2F6U2ymGel1CaOZOZ8NJw
sSZHgAGUD7BKS7WipeDjQoF+XBWbd+DW96TerK4PVvtdecQOgsaQlv/eNleseiXf
ruv79se26kT+47M6/tAp/aV6dFzyvG4x2/XK4Ee/A7we0okm8+yRX+BuMGGrKHil
ToNiC3TiYm2bzS75IvdmsV4KIWjKg7Ge3N2k+6sWocNWlpNzHnE+1ZW1rkscMAZP
BihJab2lTZ5nTbi8IY98ZnD4mC5sHxmsNP98+dSK2JmaTQ46ZyxfNnvKF0LWBjSl
YWrvgnUMWz8XuMYZ1YtRyQTdki09kLXvM9t2aJpSm91x9vXBZNhvVKX3/fMQTJGA
TRCvhWaOcgtiempNJzaN6rt7K4u0ml6j6k3JnHNX3LdTU97Wb1DFneaxXxcY+p8p
xq13VStBZV66ZX5OWTY3jV7l81xuiXdiq+UcOmjdAn2hoXJ+VLaADShZny1OCF+2
I8FQL36ILC3vsWn4EJzBe5LdgiKyuJyjhq2R/+JZ2FsMaLSRPT0IXHAcqIGZnzMx
QXsJ6x0aG8xn02K9/nuD3D9bkXXblIB3FnToACKhtZtATDriXZuWLaqsQZttdTwI
qA6S+BtHVn2sdCuvJFGarB62hCnsSzaFXr+5lhSXE7KVzWpJXXGkBuvJXjnn7yA1
VoTcWBt21BK4ikvbmKjAnO0Jzy9etrp3nCTORK8+g3zSiSXliS7wxh/+gnEY2TnJ
id7YsxJUA9FnRn9LKNCNUh13909HUnHTCtOsqphNI4bNs7Kq6KI9KOl/RLUDSKYP
p1NWGmHZ1Vpi8+e9MmJt9EDRuut9X7QIhopu81tQcSuNGWYuN/eXZxR5pJLVgbxZ
JIGS8KrV+K5xx/QSfT8jIdWQmhnF6G0Qo2Hqr+BAn9naF6K6GXPTBrHiJtkue0FK
/eTayBGwRh+BYkilly3HC9xhk1UCwYkZyWj9j/XdOpGcYgx49T++PNAC+xsMXJ1e
6Ub4N4/+zRMWcyjFT1SqLDl2lSzXq839jXH4e2323lQ35SP7tH+pqiA8vGzT85nm
6Z1qcJ2NAKUHeEkU+yiViMafeTnL7VZqkxvkIInBkIkqIQdgX35S+b91ZkApVy8I
HyJXBNrK2RsVuK2vlObwAWnpWe+h+NZD2ZqqEEdYbiFJgQ0kKMr/GsJ47ztK8ITw
5/wcFJoo8rKJte2mN+p7MNbDB13/DCuPjT76i9zT92U9KsWUTWrsscl2oeYuA3q3
C59/WaRrMBT2Y+5Ab0+Dv7OQ6iBdCvW2zMIFIP+3bUynkiCSg3NankT0ZWThSBVT
LoPEeCTnVDh7kkw/XG6zzaV6S6B7hxXWWDG4ixdOJNTtHitqlvzV89QGqWHCLjqQ
i7GGkAeUx6O13rss9bIUzGL1gqwLTHNKvdFtgvCABo4my4c0tVeyuvNi5FxGc0nI
PwGv+fvL0FVwJQptZpL/qHuig7LGugKnD7p4X4aMYni6EtO12DzZ1p3KWtnrVde+
HL0o+jdK4eXt61tLcSraXA5OSf7RXEWvko3jkOu7Z6sJ4lRrM28Sd37zstQtbfhs
kYP1WUbJd/YjSyQ8g2FXGtM66otSqBJJ6zBuKCsK79R4NKgxIIUo4lfOa1XpLr5a
iKGHIaS5mhvQZi4nDF+WBABatbTi4pNsSvA7Zy/ETIfnRogGTAc0gORdIVzwDFPn
r7ouaU980JCiUeRtZuL8uqnD8m88sKhGCR2NIt955iu+YgAU45WZmiDCI3Shm/7S
Lfmy+9sOjp2RpF5UJj5ivDiU9JsUvQH7uwiJJ5ojvMRSze1AlWn7eOs9UiSD4c4w
+0ILGaEzsjKR4YHJrfssnw69gFlZfu/mHO0Jo6xO5ZbTX3OdD+Tm0mqF/rgpDhZa
TAS6sjjijbTe1zVr5S6Pdb06KELLdJuI/gtR3dHxu6QJJnTFOcDLvFeAmnPham0h
1z1DpIM8zQDprqi+dGV1J88Ic1tIDmE4dnEHppiYpdbnTl7nvR1KurtqYgGP6G3t
7dX1mcQ2oV/EDp1obBI+C+cJqQcFZBP0w0vVLvkFxDZ61aHsKukTVdhG0qbg2Gkb
7yyd/+6rtE4Yni14YyxieLrWV691JOHh4vwjjO9Lqhy8VSp20hRQNISta9XWdPXm
OmzfTdyb6yOavpXgG8DSeUUOZUXTUockv8J+ZnTal1wAr2/elI0uO4LuB3qhllH9
J5hogF0Zoetz1RZXlqHcISrvDxvTEHbHRfJmsoietLTh/6UHjLPZSjlxmgJGB7cC
JxYmefxb+ATxxGCkXO8I71RboRRxcXaY6TZmCtSxDexQQGWIYoU8o5KatxP9hQ4h
uT9mbNMcwNFONowx7Oi1mxxpqrbefuCfiXZ0GfcwRiRhkWFEVegCnVeCzFY/jcd3
BzIn7cP2KeJJ8Gavgo0fRy/Pa0tpq3S2MgKNIz2H+RsWs+BasGCPsmBEDXYMjrP0
Gz8UCCdtrp92GD6p2ytPK3mNwh/3v1snkZL/q5T3Cs5dq/MSBVjqbY7QrWTl6Fi2
rD+e1aQn1RW9HTCsT3FNBDrmtzM/X+I7oot801e6FcHD9ANYVYE8XcTfyuVWJK1w
29av23QWOLpe+CFpGmGThNC1WWPRypC7EoHH0UsHzL7WwjkknoflzGsER435kj4+
u9pPUxUu/suo4wg669Zbnspb4D6NljG/tNQ1cacOVe60oAzxUBZFVawaAPOCGAjn
mk+nlnQaCyDjPtZLjy+9Qm9iP4Zm+CU8DOIS3ciU+iDFCTQdZlIIFAjgZaPFkihj
r6Xej9i0YgyxDFluMFKMMAvuQ/Cu3L8iyz4BYLU4xiU8wvxDbDRn0la+U6KA8FOB
1vzykBe0VSaCI52dW1yrwT5MACLSCTtd1kCK7MFZXossfdmDMmXTzsiGLPNCGCCs
v1uSa3kb12BUPvoXHrSVknrgvJkezORS/zHC+XvBO+kdftEI1qx+HcqlJTS/fZtT
Kgv/aoV0yioLGz1LH+WqaREdtifkQqAMluVnNE/c36MiUz8z4eQbmUmYgjSdK2Wm
5LLuxpMbbJZl3SZ+F0IS9KEN6Qda4rXKXU1OfFVun+CDJuZLh1pZmLrAg89aOSEx
LrFfpdLNFyPbzYUYZSq3uAcKiyFKZG13vMt7qGZjL0xCqd18TdruuYRBEhIf93mz
uKlgXrc3mkvlb0TeyCXA5UhqXK5i0pWgBbC0Z2VIhll3vk+/HZ28yar/+tDbokaC
CZVNVo5xCdaZ4/QWIU2/iLLdArgVw3OX4NfV0PyyQksaEMAvIzCk5t24mFtQ8qBa
cThV84taLqRLQ98rajP+p0fq2Q06bFgAMAAJLreEsY+/tXbxtMm3GK+nnDf4zX47
WyxUWNcBPgRpTK9VNrl1sPs2ZxlIXExGHTQFl+W/sMRSWFayjsQZHnztFllWtZQk
MWYFAWqi2q/tNgWwyh55mlqhNoQaggIA0Cd6YiZ4Aj20Ru+2Nfnr99dHBnh1QiK5
+oOrIE30sDpuzodO6JCZomnetGJ1VNMFO8H6rIiT2LL2xy435vRnC95okeu3Inhl
jMKBmvM+HF2Hjt5qWGsZ5arT5fPi75o2q9zDBkA8XAmgQch5RnY2sFjbbFXwkLTz
qiUk11UubMupgj+zSK/TMTuwoHSxH/xEVug9r+Ddx+QFCuX5z8Q5K6K0cpehNuxW
zxOP+z5bxw0M4Bpw8VlZpld3Pb4fYOH9LB/0NqpGIzEVjSwDTrtodsQDrD0cmC1T
e4htDeqxisOhCUrzcYiMTwl6o4PMEfxpuNgjvFjLQEGvwfbngqRXc1AvgFQZW8m2
SaZ43Yc5oSV3WM2/55u/nvNM/GHcQcp45WhK5xzvoakOfpGCLUhVDbVFkjrlEh/k
3LsYmx/EoOrvMccQUrX2kEhZyY/sloriZcna/vrW+aifWIV3vIzL80hlrzGASCyV
JrAyE0gjGfXBBuMb2xcJ+YkJmxsFrMc7h3rvl7lfqw8NN/o85zYeI6CujesgZ6am
rHtgB+Xm48jEQcUyp424mTpis/+hFWeasnNRf0RF5X1dh1sIyzPoQfkWcyX2xcxV
8B9iQkrBpxWqb7LfWESdJsBe8M2mDk3PQp3/9H5QURoEP1WIh0WELrlRE2Qi+VoO
ADcxNQCwqGnF6Q7py3UfmhhQ5yMzP29Iytkc+1X3zGMdlYCaebvREuaa16wl9e/h
36iURcVAMftgl6qLgfrW1BUUfmhbo5vUKhLjM6yDt0WP9wvu3WllSwoenS+Wo+LG
yGhWYv1enVSJJE9yiYpA3eYuOrkUMLscXuyZPf1Irk1yD1GL8seuPZT3gKq/YzBG
WArysV2SHMj6UFBJPALen7f65AN6NgfhdHuWOvKd1XXnWTGkpFE4QZcn4pRnKpp+
5QafI0sqhcB25/Ja5mjtSZ4wjIuY8GLRJErec7l2jnWtkZwvJ/rabLP75ruXJK81
roGfuNZNw2oAdhW3xZad6VhaMqea+RASuIcpI0X6zHTwxj4ovlJqGE0qYwXixubP
DfocFmhE3Uvm6QGnAKuE+m7Bz5BH83v9PbPHHMYvq1XKppeAyVp4iuZeTVqNuGUk
kvJlShAcasrZAdZFYIUctpDRS9AUHWyCkQ4wXLY4omXR9D/JGkzOgXBn1JHgqbka
t0Vko/bkR+xdO04npFk3gTNXI9/sO1Hey8r4Spg7L8SVfy1RIMQz/sri2NoTSGFj
T41979s0OiFuvtcJlKYMxgq7zYvTIi+z2bIs1+ulRahI4ag2Nk7USkVorL1RibyR
oa4iQytQNjlQYa/C7JrkjvbYODSPaw3n8OL9pseViemcFatUrlJeWVb2u3GVPmQA
X4OBIJjc2v03dHgYME4XSVOchSZEv3h4pCkBlSrcAHrS8rDv0V29jUcPFwdTDcY8
b/jUgOoToY6dyM1BdsCFdhVqtFPZXIclnzFM9nH3I5iiGmvewr6bqhGvgDwBn1oF
OvdhcSoY+ycOGSvLdEhKHzfbqHJ1AKnzidEqSnCVLte++kYOTSfWL5cYaTUe2gl5
i5ZKI19MhvsZxSyBArwKYovv7sgbU6rPkmOSco6OA7SJgYCz9nhCx5IPkJ7VEXs4
KTlMLGZMpBWIwus1zDh0AYOL7KnvaUFstkUgqv9myF8CNwWGIWssaFBz8gWZ23WL
lTTTzy15NKleg4Y4uZGoGIRT858NlhvdoR4nwQSemkn8/JTt9klqlgOwoLpI1j8E
1M9oIoqfW6dA6XV/ouJCTbv/pZdMQ+Y7ZnnNTYH8NspVYqAKreW3ayitwGYg/XID
9oRvFWV63VrhqfT2qPzyo/u5ZdIRTRJJhRWjtU+A7Mm0f8w4F7w1Lk1UYdRZHp+v
BIX2BKk+9mhsZ0f2PMhZT3TJOu2nPLTmZEMWvt9fcxk+vK++MujETDD3lEXSFdA2
f8ZJcyAiE8ExPgwwzAqiHBKPd/kGUBmxNiv89clS77VrN2JauvMGBwSY/+Gpw0jQ
Dplw0wAaMWeZjrrFO6BabqjiJDhCXtNLphXs1HrXzgLpbdIl0uU7DCpWnCrMx5PV
eRZ20ba3l1zee0uAevFSDDoy1rrCeB+IzSF7jlA0DT8INOoY/GgS3vsPeDUpaAik
Ke4SMlqoJb7nBrTYGxgFamU/l1TwXV00bJy2Cf7ZD4B76FZWmhS91WgDshQrFhaY
hWHaGRbZCW4CfesTaFjz9rcCI5SEqrtVzfB1trG53kI5zzYto+9keHSCXgRW8K/W
fQGDaMZcWoCUo+Y3tDCm8qoKsFKeZOStqPi1ewfYi4YY/1Un0gNkMvRtkuKNpa14
+7YIqu7abzxTfVHMbNYEk8/WybiaI3FUcywe3YE5CMS0ivpjchYfK/O02coNP+5V
TgtBjbgVT9X8P8ig24Objt06oaZ1JtBWkaYp06j+ULii/ZZrqu1GzrZ61bBdvPV4
jqxo07GSgC0X0K0UdtbBOdXquGgMAflpP9txUs/mu8INRfTAr6Mlym54Py7R/Iqt
7s5L26+xLYQ2DgGu/sycKJuV67jxgGoSq0u/IrUwldWn2gB+EmYWrtYN5sbFhN0N
E5naCTkTD2v2n1EJsAIZBucn89KvrXNEP0MJY/YrrzMkN4vyRi/4wB3NhXHxKL4l
20vP3INrxAeCttKEbsgdOOmuh+wYGr4wNvlfWlXugfI0ADF+iASr3FkaEAuAwfER
AhikuRxi3HnodMdBIWRT4IZrATtSV4duA7S11JeBjJf92qLW8H7WAphShSrba1w6
PiE1l/69Q5k4bOn8sFHhTDG9jfrKCUwfBaxE1zNIZB0pPFmQld6T7r/1FiNJg8kW
poo7bR5pGVutNBCj5uaLHUVBbpGSignkyRmM8XMtiivQvqJlWtTIH1QoUkUNjBEH
9/ZXd9XNvzEo3YeGe+iIPR/PgynNEupVjr+fF4RhjAQlG1jfeoaQH04FLDY4ZjUt
6b5dtDejpEOri0UXhxp+VOFz1kE7YTphpyIdEAhb6N/C91dAJqxlO6uITa7J4eVP
yafS1ETcCBf5s57pU2hnq3ZGEGhsHgCUIJmoOMSd+dAeYqT4+1m0qXaczlMTffd2
X6gYRhbD34sWwxAeNS0xSHLMjdCHca3qTnzf3oyaZV1REYH9zMljgEVvte3NdtOr
Z5VXW4v4SPo+pk1x9b8fg1IZJlm93MipQpSH4TKu5mfH+0fqFWuMK5L6KEqpZ74L
OnuPEM6rh5peb8TIoYZFSOPjAfJWZjtzKS4NRlyQ5mRiIiyWhnelJYDZPMf07R2U
rag8KkSAFWF4258R5LRVV20w2hnJ/Fy7C41+PC221VIwvfuHPW3fkuwUJX3GYFZD
2Y67XIF3YaLynClS1StGR81PZLnCdO8BeJW8I12SVjXe+QGjp/QTfeyyOujwcId1
yKzUUCwXDgkPSXob6EjvArXkU0NYNa6ad61bg1QhbNFmOFcyRrmYOQs87lcU3NmU
o8ZAMakd1yB0IiDmWubXdmNB+noU3qLsbxSWJ0TS5WT74nkXk/shpdjdWwv5gccO
56/9+PEKljX+8udpmEQrMYSLVgd7arrDHNTbz2oPgMo8+1u7bVK3h9uoB0bfKp6P
pxF+1yc5Ik7bH4BHrY0zbJ1zptj5+zN3FhS9dMnox4rcCsbjHQKmSjQhDiynWV8e
WB44peHL/BG/1y7HoM+8fzwQF9J9UDxsacVSvakRmqmFjG489Kv3vrKr5FQLl0ow
PzflRgYkas5SOHYNXvTGGAApTj45Nol8UH9xeD5yE+gzlIfOMuRpOjLcr+D/P3Za
On7TAm0VY/JlRgp7Og5wiCWhjJT4Cf0HJz1jM5f0Spgo7dfrj4xxSWDwUoiPyTyR
IS37SuPdWta/7hToSDvzfeoSonMAje7xEKlJMwQqYyHGk6fYtN1uDaeuMbKGrHi+
E8A0k4v6+XDz+8cQWMw851mmpgbAQEhTRtQNOrujwS40F5d7amVe2RpGGKjADrPI
TNowTY463/SSbHIcoW66KbURC4WJfHWkwDLHl2+8SOlXi8fPqnLw5QvPH1bVVna6
WzuSC5ZrRZCfOdaf7UPLbpjdhhgKKGSDmMA0XwURTGr1RqUU8D7R2vKM/JxlTqXT
mEq12OeB4TF5Z0Ou69AVqHGo1vs6V7sc04isvaXB/WXhLbvchUAgAqUcqsxFg+39
/NvV3CdpmCDWYXjCrbDUPrhaVe+U15Xeju9udJG+A9c6Wmu36bJVsuvL/yf4p9hN
lrEuwdm/VMsBiHgDlDajw/6D/TymMJyOrp9Wax91Mlm5tOLC38YKr6J11pZTjlDo
agwZBrZNsyZWP3WqAVPArvBy7XoUmxRly22xEMjaJslaAF5zEbfWCVV/Bv0dVo5t
xm/fXxTopFTuYdUVDGwrHwbphdMKEL9ux0b1B7teZtgfGR5GK0uxtxnrB9peUjFu
111iPwdN/0A4/U08dVQZZ+nBLb55IcKMS6ukYJZ1Zbv3eALWrrfMGEG083had21J
J54PLA8QsfQLhCSq9w2DFWCWOlL0wurAEmuCQWEXerZQwule8NuKgfOa+OPMWd0r
bQARJTcf/18KkoI1qboIsU/HH4FHbl/0uT1h4Zap35L/5dl7+dTz4EdGF/iqD1mv
R0j7ynqriFTL7vEaI6cuWEeRcFkQUprazmz2/iTr3euuU26iSNBIWXBYAZ1beqsa
hvI88BomxlO0eda2eCR2QznqQh+dlTSDVRDax464v35OYSR152rdw8DZ1PGUMAPl
omqia8MisgHwWR/g/YO6YOGZ7ufLyLCx/1QvgbtGQDdtDxYf4Oz382tw+/Bli1p6
RyRfOp6/Ew4XCcy1KMfrA8+hwDsyZ0kF7VZSxL97Fvl/x646+VXUwZJ6XOtAzVfT
9PaQSl1S95IJUl8Y8yJFfNmjqGk1cuItn41KaqCXf4JtPmyK1Hg1yUPUyfRGMXtg
LwP3SRq9GElfFZbikizahGkyL0nfy0WMn5EGJF4H+wtErMANrEyNXfNuOwqNuik2
OEnhc8+SivYowYR2v4ucM+l7/9Ql4xRJkW+eNxP9ZH5tlI9iORgct43YmS9W8nAp
ELZju+DDd0lES4X7CbNSZZ/eUFlKKkvHADA+JdPzNse1ALyHxozwLe9HRH64iYRp
mBVlyfrpoJ8uXUJqfB7BeA25m4r9E+Clq4YeHs4q/B2hoQHZqFwpFEe4oy/i5yT9
0isRnz9wrMtE84RjarQEYwfkwJMC54k212DqxXyiP7uEGZ+f24/rZXB+1bDEHyN8
huZWoqwibt0Mo6hmn8y19zTH3izNhDtOEKq0HhplkUuyakBPfRGvz15shSPc3xCL
xde8cOF3TmSoSL9HkAGQlA5kX/MGEAlwBh2dfXPMmSduCyekoMUEqunXR7lKXcQX
/yaNgOJTTTwa46TXxzvzb4RN5e5Bs/HpylZtzSkjm8d+Q8fiQD6DF9GEffUg3SaH
Pd5MvmLE+AXU78ueS07nK8MrBxW/u9acZmyAcjp+SYa/qo0SbRF9iyU4zBz4m1/P
inJg/RShokMUiFd64tKBS9fomyMqIt6uktQVD1BZumOEb+JSQNqxpryX97xQA/pw
aS5LWn48j9tLqUIFuBRotw52dspkmta0NReQXpp1yqLxx111y57ofE0/hXMCXVU4
z9XXu2GGPC0N9nnO5Fr/S8f7rPY1AVPkEKpNBGfC4ruAKO5oCpsmQrPhuIYFkpl9
ZjxF3y9LX/fa+jyuCydp8AC+2rzX0Hkdoe3ctmrDpbvzcCAsdgwwaLBi1swpZa+A
S2OFtwQ37kTPTTFf+bS3zx0Ht+Fnf2yEbuP1+2t5It6njRZo/zdjGe9sjNx53SU7
TKBGQXSZRbUqYXlJXjn3x/mplEav+o3WvhQw9btWJslhutqb6n4RlySa0rd5L9zS
bpUMomQVmBErSE7iMVjLOuZEJnzF312wf3fHXEpz+rv/VEiTAtW7+bp0u0xtw5aG
FrOz2wQxYGHe+JM8WOKJCJZsPNh4xsk8Xe9fmJabWAkaUaKT0YEIgDHpqiCE25wG
o+tQN1qCd3TbC6b9SPe0PsZXdSa9WIn/p+QAAi4KBbYh2NHGDNXM5d5TZpSi5me/
An6+pUXVRLwxQ+E8LeRJkVftjTGojwKmvgrJVcvqzRV+er7h3DVuqQXsLUNGFSP5
K0svRc+hdE6gGq6V3NAmRU98CtrLPX0vKgdlTW851HgGUxyehAOWwZIK/neoNMka
Lvdl4CSlicuoZ2kCMgJU0xZlCa4CXL0szlS+NRp4En/1LHmlWp1aVrT3zz4yIeX5
3mJK9or0b1ABJ5/lYzi6p9MGrnTFV1V5YYrGHhIJbsvBAp8Q2MaR06WlNU5pNxg+
VnnvCOjSKYEm20o9eKiNEQxpMfKB6ktaueHcSM6eSkMEytNbWmj4fxBpI57lfd+v
m2Ks3OakwBxaCk1WEOfRbwxHDB14vDYhSw6JhEKc1ihpcxlHqItAfWpt2DD7WN/s
yeUT8Y2j/ypoh9bkbfVpw06KmTn4bYTx90r19ggVtQL/vLmMf5TpAW/XNVjvcfHd
0PstfBYJaRq8USSdcdhfwxwZaE5IC/zi9rvlYRJEdlj7WA4eEELKGEMSRF2fH1T8
BG9406iE8Pvzq5mguvcDutn3vVbmArzMNTxqO5JMY+5ACWm6P9s3Kh+kktyI3P3I
3QWrsz+gIqdBF5C+JlciLpCMKQqao0QuqgYaXHk28i3GUwZnH08+JRUxvkqeNVHF
gQbWNBgEvxMlEv9pFBHCDh23nPzEKAvQvVftEjG6rTgbXcy4oOtcTNE0v0gpubAj
K9eVUsei5f+jnEJDNoTgWA+XyGTHPyAVt/zJ8UuYCyvqZhakJFEN0XNKlaFUNKow
TafvQQXG0qJ79MqbM4z8+bJ6bW4fxEhRSwhHeqzv8zvJkYHgMsOIZriOSfwqEm1P
xKjiu08B43l4VjXsimUfveEG9d2xsxM4VH5loK9r2WOqwvdZifW5j3XkDUX38Vyn
W7oJ3YZ6XDaWDYhd9qg/mIYQN/LzmjWCIQgjiojQJ3cFNk9m42bQoB5abvtcr8v0
tPZEEWb+S9TzI4GTLdqRKJBxEl7KA3klv7Xa5atbuBAEW3rEirj/1/HKYz/slXCG
TfVPuBB9IjFwt+Vfi/m6PzA6vZUtuQTpdH2piR/Oyqv9FnA6x2DjYmssr4c9zFV7
VGqmhGnj0IujUeLMjI4fTjKPgn+xY3YhctPyOUALYf4daSJWcG+QrLext+/5K8hn
aZ6+GJfk2HTcOL3EIxq+KZvt6Y9PAgxXp1eFr1yH5avPgb/sCgmthgBiouvgMD6q
h9MuQNe2I+52sRibb/zjWxiawWCEpxTnMbEpSVmKSEloV1LpyDwtBX/lwLVY62Gy
ELF4qsI+btZvr3sez3vN/8NP+cspcetlNhXX+VtX8bVGyZbUVS+sG9NYxSBgSH1d
4d8fGBOdXoAw9Y/2EbPdiS0jsaMQ6kDDPfKlxBImq2fM70Ld0z+K0fWWWsW8y3z0
WAC56ZKPQEhYtIKZBy4YOXQeKKw7LOvgHqfQ4xN05Hi0H6maerP92beuFr7u8A5x
doW8MkgOON0Swp56rG5/j5tcyaRpOJo6m38XM4JCToQxteICnh5EInO4TFWCFO9z
Rdveni7l7t8XdCo71NXtzVWQDEPSc8ZUIRn7kPkuBpn4rcxlsx0iqAKKCq0ld2MR
DsVgnB6EJTCwXYgf6HSqXDRYJr0SZKx8COyiPsWefr+l4kB0Hvdxjk2FHQuzHqws
04N1zv/ZhXlNpJX4ZBvZHU+cLtCQWG1mCJhBHaTlzMsOW3oN/I4PaG19fDRsFiyD
47bmZi3Z89wh6FocBXn8gPFlZ+dKlGuq7RD4XGpCHH2aJYGItc2/za4BTsofj91A
vRJJimf00z2zUFvJGvzvTSfexvl+gLZ3+hAnXEqqzRk5GHHhz6BfAKR0n9gmtaK6
ZMwHarKtMu36rZJMnxHOtubtjkNLmOKFEaKjPuC5WI83uPv7kLf8PPJPjyx5dhTz
mdJc24p3M+zyU8/wp0wfKVQ/Ydfj/6UMgTsGgL67pZ4IwO0PeuyxLDZgo12qrKk+
TKCt/4c7+fCCjlLwboj6o0A0ONc1LHW9UMieRQck07kLm7OW9UcE1dcEm4AMO/km
S3jO13pEQjxOA9LHgF7Y5CokX8EfS3KG+ksYZu4eS5DTSf5C1/GGCMENQsvU05o2
uKEG1A7BUZKcq1TMjNJawCTEDnhZkVzsdreNWZwiY0mHAS31k/ROO7p1QOTWSv4G
U6vjWM55FtkLHdpN0pdPpU8EXA4+8GY5BnPqhuVRaTKmwT3B/esQy5GjHlLPt8RZ
kXJptry89KFLZcPPN+JbxO9RsgmbyAVrl9NCmxSujTKOvpypzvsruAYJKg62i+j0
WkcrLalrrPSilUF8HH+oPBCJeLHydWFqsM+d8/4t0y1KfPIiINvYGZR/m8qGY588
xmGWRjsGCx2bIYyQ0zmXpQtek0RWPLGuH5XVh8OQ5NEiNde8QYJVzlrvVGwyCmbO
Xw6h2ElgyqwmWFLGa1yvIYWyZzjj87ZZiO7oR4bpZjdo3MlTUEKm5L9WXUlrtGIu
VCW6VvLCZcQ/jDXmTJxELCtIaRD7tdl31HBhTqAut87J54jWoUiS3cpAxPauYhRc
tILrvr0Z4EyQEOV9B9/zg2GgxjdMRbEsSFZpoVzoO/oHVuXIQW9ZuzioiqfpyvxE
4GyQnJYyNISlx9nZpxPAnco7ht9NoNMhCyL3Cqm2Csh0HUr3nBJdS+TofQINz9Eg
FHfBqFktKPojb+q0DrI3QJ9pfWm/T67uAcgnoKbzL7IR8FRMVQunOgllc7M80Jiv
6CXm6KLzumHVL8RQmFPmqLAX5CvzTshiJtSAHEuW9c1p3utGgWVEMlhRtErSyCPN
yHz956Yp0J0c1qciJB09OBf0rGW5r2nbsJ3xFYEcjsgqsU7dWTwsjxBAdUrdMdWe
ATxOFFgXI2b+vl9HGoVxFHHVJgjdI0TAoRIbQzQ8ZRTf2afY0peugPAHPC0sE5cP
sw8l+IswVDZYcK3c6LQ2+Hifvs8UDJQHVWd1P5/OLJsM6S8PihL5s2ngqrnSYed5
sS6fS8jsHaPCuMBLt0UV0EjbNI5RqS/0Fy02PGlkjn+Tk8lzKG3jC0ty/GSevktU
8V+Q1JdXYfvbLMCD44s/7yfsL1Gy0eDZjCpuNBtN3Mf0bgTXfM4pWe+5vtZfq8T0
eGuLom/rzaCTYrt340IgfzWV9SJlGjMgg/25AjiF7N0I1aXheU8+kSYAZ9DzB+uu
gGxjxkyiPwFxwaNKQn9kF19jr9sDeYBXPSvvF4hadwh7M6KPDctWyTSddFgXBPAT
j5PgmsTHYZk4MTcFbqD9VTw8bUDY3jZGjY1X9BQwxdngegB6ErFiacX86c+GRTvn
Jqqi70trnySW8J9mwD6NAs2LWefVq3K50uNBcB5Ki3kdQcoykUGQeOd8pI+OGpoN
xo9BGtw4++Y5O859oeYdwRb9duYJShWqX5aMBacbO+kSkDcesgbUk2CPb+hNnc1Q
Xmc37pvKmsM53xlekf4JLBqlFN7iAHslL6iL736luxtTw4DK0tIdcrTrvPdSNVDL
UO/bIVvchtFHheI950AVxomHIoClP/xPTPmbH6nZSGiO2ezcrDXhumNjr6oc85rT
SgRJT1wVYsdJ4fo8UB+CZQMtM4zDjgGb6WXm9evTsXObk2E4CKUMF/p5D298XRIl
n2zPTVuIkAl9Hg91lY0XL3UEacEEs+xE3IhKsG4+ynHwFXtrgKFRdxRw+A3ONpws
6kOUHimZ3z1k2sYyFfkzEMCa5XpwrbyXljte8XvCJ2myph8hxnxX09VH3Kk0mOay
X4rp0snrx7sMIunLU/Z/xGt6b8lSOjcTKdAHSDEXV6gekjXBwCdJv+1ax9fHdsmh
h6s3fjXkaoYdWdsVLFil+cN8ALTZqMm593NHuywPnGCLfHWkGocqSq3u85HiyXPT
S7DNfQRXlxXXSOan68jtNHmN8yqJHOEjUd41cjjxpXIl1qcK4H9BQ4/uAkjyDPZO
NvDpLfaC23ohmQb0TSfTi//un1ugILN8bqCdP5Wi7qlIpa48KJROgaIIQBqIkeFa
juJfGyY0i4ILCKKbkqf2nIrqy4f46ufFUQ9Sm8YFYmzxsD2uyJ7Bc7+jEKp0qd2I
S5rQP6m7pyBcRldsSR4yOvzK9KnVQb33QDRdaaTIyBoWtWBS3Ep5+eUqS+7xtSnP
y90tMeEqXJI3KNvVWdIVp2THZRbrbkORuiyoVFSj1hAGa6Cqbrj+FGDprWsGo44q
/3tIsT4bUQcIBkde2HZ2kWNNY4AYBXvbvWFwAZCfF/tmgqvHhjDSlKS3R+eNRmO8
Kmmu15CQuZqXubkWkt/IeIJRjMtQVsK3ua6a3NLDfch1USBxbEy18udEcnreMHdj
wSQx5kXLDoZruzF1M6aD6uOVv2nVnLB2GPut5x623cIZrQBriVuVOfTvIg8zGrj8
lNzkcB8EbIn3dEl24z8fPZnRemQ+C1bD8OJAlrmcpvciFVEwLQG6qRw8TECeDTI7
y0FxrTYdRE+DffVDOHeDw7dkOqSgZEOfjh79mvlxQCZMCbav9DmpdRvWqo/tlYkL
sF/Hfuy3RFjBqUyco3mBJ+9GFXic8uaJHDTSieSJxmYFBuIsRunu//h2I98dzk8U
iemzyLqzEu0TUXRD2ahRdLeaF72xTkcYr9M0fcCw2GcWOcUJXAC+I7tX0LaAsXaJ
hCzSNRfPA00/Q/GfYPPwNTorhnmS1TU81eryEuy5fUFyfmMm+XTa/sCaV1jsDt1o
R6BJPYyMV6bQhjFYppxW1xIT4l0FnWrWz/IcoKeVeVpvQ7WcXbJ6y971CXSBxOLd
W+HjqY1wU1fGfhXb5rEFnZcABgcyVm2oCUAs3cSagJcvnCsIDHWdUE9Q1QxdhTDm
CmT8X12CwbssUEjbspxArIVjUsbRPbPv75RZYvF6YzmjnzRWV0iKqc3tfON0fwjN
YgrJO4qM4hRmg5WAliSk36UUSIH1l5+UT4YNFR6P0cGhb7THOK0unF56pArMQuh7
FcBnLUtmK882iGNYQ9y33XmoUyGMjG2ET0ac4MZKVH5XmlEGz3LIejBJpG0BcpEO
fNZJzrX6GEtidXK3A74INifF0J44HSCe5I5sb+iI4+jaEShC4bxCnNbTXrZHG153
GYUC7a6vbWVP+wlfbm8BEd7G9ZrNCamvUXoj8/1nOSx0yOj0svt1nse6iHYDvxO2
OrrJBUMte+yidT3JIUk7APHv0Jaz55+RHpcLDGWRJlayh0KcxQ3xFPs9cQ8L/tOj
jVq0eioQ5XIcR1YsuCpCcb7XYjPvs7/98biwDoGdLo2aCGJy/4YMRscIUCGfEHrR
KvnPAt6iDA3pOsaGqNDo610UcXX6SBUEwuvP9sK5QTlyt/0ZkzuDkdFy8KjOKtf5
EI288qPxKKhVb7p49TPiuntcceRfkLlC3byMzLFFZnT/YXW/1LBcahSpu4DDv+Ow
MvPRNegp45zPknBXZn5PJKnrsIMcLSWmkTFmjUBdx2TPfetg84xg/R1rJj9DY8UJ
MBSL9gxsvXXFOe8WdScSKl4GgrCNIjmUlpJh0kTp0HSjxxeDIapVozD+MQp9TqBf
euRam4wc0MhXYcKO/rMcVB5Jr09MByr74Yekpn8aqHEu3MnBDzHykP3wqnQ+Ob+M
ikkOQM+4tIRMvqvceyHZ3ceQkdYyyDUF1b6t2pqtUcWaZWXUtRCf856JIpgJtdrk
RhwCOOIwZeVj6xo9m+hecmC7mWWsinjil8nQnz47ptTvJq8JkCpikkW7XeIbMWno
S54vzYjKx/qi5xXpuYhQf21JkOsPyjT8D/KZqovyfRn3wmd9diDb5dEwlCGoXvwj
Hbvz35sURrAfOXNQn4Cqz3CB420GYQXKrQwqfkFrAkHuCPMyQKILfIO0jDDj/9eG
Z2QIEgZnmQj+k8kRFWHGrF/wNCKALlE7+i/HMaU/Vm9jxFk/aMDX3S9L5cuwyYZx
ao1ybJvJcBB0Ro+mY8l+Sk1KK4d40IzvJ5OFIdQ4fztH8npuHejBFJcqidpVuvSv
TqOy61GZfbq34izRwWRQwkTdhNusi7NBKRKrpaEkwp8TuoLW8hmTVPbEJ4naHUG+
b8bzzIWlER/DOPF42mCoAP9CoS0Dunl4wMPqmYzqnd/ld7/UWsxwvfs6maye/f/N
ePQQvFgmz7yrUzBrttI5b2GoO03tkdJShv0agNwFgqmLwBhx5DXywGOKm33RM2cD
w0mcBrBX9G7Q4c7FNe4bXOxyzemGKjAAabKIFSRZjrCanlA5E3T8P6MZJkSHXCwn
iqKwKyIiyu1IoIB2OvTGDSftBRfAMTm1fTw5LgN07LBNAk1WjH7Y3UOtHloIdF82
han1uOiA+KRBgkL3sQmd27NmmwjxBz5ezfLUCXIEFfL/Pys0rMs0TrCLgd+9Q1CF
YcfrVCKmRhZTKQHsOjJXhlBz5E8wEKtM6Rcp/qli5nT3ULbYkRjWt9buNPxs57AT
LAm1zUrq5ZcNaItuivV3kCnNL/i5wbU6lfJoOuAHYm5nWZ0zky6N8kS9vFhRyA+W
PdjwNOI7C+09c7UO7zdGc1dwmM6G2hz37f96h0CTOsBRuhBiVCneUWo+rP94SRC9
CQ2ErJh+ahxItkqABVfDLnOF75H9fApnfC3VOCsydka2cM6xc5eXmvyN8HSGjcb2
c8HMSl4Ke6hK89SWEYslmdRAxDOYXgXMSbgCEEU6y5ygbKYkh1m7Y0YWvUN8Csdt
bJzyZtBIlZZFHv/zTIMkN7bUlzaJ0Qkzg7BIlsZMXBuyPll3A3+uKymTk/DukatB
bT0qL6XU/EyseqWjZ35dYsDmNcyopNukHxXHjc4kmzlwRZ1WX4GDkLp4Pdlwa+iQ
uHoer38aLDC2B0G+7smZMADvtdqb1YMzowOnB7qjP9hAluJXIKcqKmsz4+UjMF5/
Ti/0zVr6f1cOyruYeP1Ma2xX5vYSxxi6xQDGGsaj9FMLSp3bSL2vh/NM/r7LpZCt
u1ssBLkDpizd84hNl8p6yDpe+tGhZHzUoANNhR3muJwTnkpDVTPUYkxD3VXl4SZw
t8lm9fzUYXqusHf8AWEelL65XQth4rk9oXz+L1b+ilYIvxOB4iF0pIFa07gmjWTn
SjRpMh+s+TevErLgWcE+5//APx2gteGlQqJTg/Xv+qBdCNS0Du6Q6U4F8s0qeWv2
VTYKXo1GivSCowu9aAHGvcPufNXDGgv8lrRUhstH6KHR7b79CAZDib+1ROeUkIMw
05qJF6qvEEKGAYtBxT/jiNnM+kEJCyiNJCxSN8Uu3lSkQjDzXqzT+ZHxibt9MY6W
ml1nRTlLjAZJmtlvDngqzO+q45WiDoRbY7swC/Q24I1jcz0GqZ6GHOvAkeYZgHPK
ta5aSeIJAr/nTIcBPmS9Q3bCOqBaoxquIv4ykWxbJul//7FpnPC8PYo7IOslQYvV
9dTXb5k0guIliTvzVVIhTC2v7NUpWj1cLzbSnUtjyP72DQ3SnL1CYcQUsosf8FPq
7p4hxLEHcsBoQq5WGb4sKzfmYrAyq+Si2+GVXmh3etJt6h9y8YGxeaGI7F82o8iN
V4kOvBsvfF9wSdRl3Sqb3r8MCpqpT/3CumgrPajmpFejkjhIHnOsXNv7crzV/80p
AilIoh0kAp8oGi9WQgWWywjaDo6XHT9oyGMzqnqhSMFQ3SE7PpFSVMbRg188aWu+
rx5jmP1vxftrMMXxZ4PbCQRK79bg4maM7GA2t6C/3QKYuuaQNma+GST1ROsJSEVv
IT0YofaBAXpG3RdLm94fyQdKUzn4xT5ATiS1t81pEkhlfMR0sBZcl8nQ5QUIaYKM
nYedg5Bx8E6THcrHtoSgoLIrEeJDmXXdW0lBIvowSsbLN0Wk0EvPOTnMWY/VvGWk
vzMMOp5yqFN8hh4MNLhRw2yTiEvpQLru5PV+FYdw7QUYrJ7Tx2T0bqSbQFX/2w4J
4oBVyAzecEG84UUnrgCc9+8jsejriyDsCFXH9dM0n/CiEHDNI+JJozlGJvc1ixzM
8BaZRT1ehGZe4eVqAP2YkaXpL6I9BnSkmRFIirqgt8BFmiekMdgevk8hoYfZeA5K
KMc4wkmZrob8V1I6DneWyKttWiD7HU29hqsUcCR80/d1Gi5klPyJemW1S051YcHU
UZz7KhxBTXrP1qPYIryWzxKp/ECA7U1cujhWavqHPafUXByu4h6Ypff0alPDuz+t
P8CpukbGXHPPKx07zux8LtXeXh6GxIGEcXpPKqUx8/4wCXgyp5C6rDZp8pT9RXk5
TQeqXa6A5AbrKPHt29hM09WFndgW3nyWLuTdh6DFioWDXXLtWkhmT77l+x02B+tO
YNQV9rW+Jmiwga0RdKJW7/ydQWbv4+oIqNSIIszG+P+dJuEB0cu0gZT+x9/LwTLz
P2A4soVZVlAxZuUtFPBXjVEjIgPVz1KIwBCbCgPjsySEQE2mkOXwcT1VVtOg1TuJ
ZluoeAGSLM+ktBTOIPiAKVOOtBRBw4JibeyqlAVpRobFITLXbXYRFxUiB0zVRvMA
rw7FhyAEC6qbFkXQy6zdHDutVhIunKZzSphme3qfLGW2w4HZoj82jykmNH008/kd
KGwlFwYkQi+ocOwRgcBorJQfLAethpMluovl4XLdgnYkpvdcWgm3jRvTBhcRd+c3
k7iwOYk2gGnZw4tb0SkKeei45e2Epj0lFgW11GuWcsWAng6yniPFAQbyVD++JNVB
rKQm3GXwsw0He6Jp4MnnrkGzb9IE6TsYDzikmMrqs640D/TIpBFj0QEF10B9l1uD
s5fj1iU6FVBmeyZx/S3Xi4lw/9X2SMSfNLSbnr2nVwt0F35TbUsJjeCuCCzrEoss
mODP8+lTlUOH8uHkFs25Ls2yJHbTJwo3+lRvhzc6qdvAH72HwlUtQnHH8KksRgkP
hBGmHqsVda1TOTaJcFPLNMsh+i2BBLEbxL4JFdO5OAfWRHogyfFIHGQcCzTJJpF8
OUk/81rCDBpqxpf+C+ysjMdSFQiouExtBL/zW+mi+GPVtnO5H57kv6ls6Uze7bQd
ApaBKyFMvGBWPHvPB5gfWyC7Gua3lW5fELDQXCjZJtT8u34oqTdCaHmOu2x9RH0O
qCPu6p4kRtfn2tvJ9OMOz+BEu2q0wRUS3GAy+S3anQgorOfTOaFQKzXetvIf9wmW
VGpj6vIxAi8kNhThR1qIw17xSVJOntxom7GAgUPeEyne/WZmVLdo/TaQgwLSxoDc
LxXeWR2+xEiQOMi3LTbJubwXUBq2sXbcuPb4z3nUAyGBiX+agpHcdpHWgYF5sl0j
2a84DINq9+qVj7ghZ0hEMmhvZDcbwOAbSyQfns+mg7PIFr0RdrBA/ECRANQOv6lJ
H7UFoiGOgLrwQLbP0L3Z5ZelU/jtcY6wQajenZqepp2+UhmYSlzqlDI9azaNUkVX
Zw1OklVqWxsbsptmOjmrkpU8X2NpUd+kFemz8Xf8tgZa9lwS018Wcg/6WP7KSHBZ
6hvfC5sXvkUGZYIcYc9adfjCfHksAkB68Ql+oOn8zgXJPWen0yfGFdraaUq8pRrQ
6XEW+tPf23byb82w8AyU8ql1tRpON1CG1+35DMvGSXF5je3RwoPbVitLBOm1lLw2
vqMs+2riFTrIw3+yJcQNNMt+s6/uKAf6VTXX48W6GZ+/GdJ3KJ1TX97O9+7iMzME
zPbV3j6SEIwdPANdhfKn6Qs0kgIFvpFRJ4+dqu+C9HldQiYY2gxNzvBFPktURjom
E0HAknZ7ZCIu0NIwCgXReAQ9EO2Rf8s40PZUQ3EEbaHzrgAaPkddrG4lH+ZBW1c+
LSq2WUrgtm8l4useQH3TgHwLwU+UyzYaWd2UWdMwYsWaZxmSCyzM2rk6FiGnuMLj
j8bcqCY5sMpOMGeODkQj0jDq6VWzb7fEtA3poMdfly1HGAUCAbHDTaELNpwwpDF9
BPOZgm55mAzJsqSHsItIX90hw332cpHLUR/HLvptwZ/nk1EjC/9glPjKZNNMpPvq
iwp7J25m1SdoHrd++KLylnWqs4QcwLx8BwfxvcUWVGHXqCj+lyLOfKy2dTezm8XQ
GAdFIqL/RjB3LjVvzr7/i6opU5UUZBim8hpa9nKNGR94CJ4BHvIXSpXoqoRQeUuL
QCD2juc6zo9h8bzRu+19QhpvsvIw0hMjeMDADUUq4F44Ph/DEfpwnvJyo3IUVwk7
niwg9UYUIgHoLKPgnjo7ufkKUllGj8PsA1zqKvBCk7lrgvUnLasNQq7D8I+TL0WD
VGT4JvC64zgYFBcjctFei72d38l21SbMsWWVUIpBlAdT7b/JI9Fqc1CKRL48QoAK
fmNLVaVKRer96wuViaOgnJ0mfxY7akdlaGdn95kHfhCT7I+X1FD3lLY+tN0GGm2w
EMEw/2n5oTETnftoU9z70B0uzQkzqhkXDWMCSGuP48SRhh470Pt/c6+4PTH5q0vg
aPlE/da6e9mrgJGEVh+0blNzoZKCzO5uROtHZtnXow1+MeFcFMuZ2llRfTvaKrpm
sQCH1dL2thu6xYl97rIs/OP//RG49Bq1Ed6ygeyY4WVVI/Glw4q6MMYNiLNANLYG
QF4Rz3/V7YAbqWeQtAqEibhxNtGtbirD7l7Ritlu/VtQHFq538Ituh+bIKKGk8Oz
N/w8Fu/MhDHOMKEr42qvRi3D7hKpCi1y8277+yE6u7LMjrp58LW7LVoKaGvKYETT
X1J++2z0mRRlmPMzG3EgQ2fzGsbZwPTXHFSzLQ8jInaiNsVQv+foVuiorDD0feKY
BZJiJ/CT72daL+28s8AOEExcU6TR2Y/0W3KYYIgYn1kiEL2mlgVuWL+7CYjuUmXe
h2cL38BXaFocHWfS+mfYzhA1l5zEci/mKz8LBv77T9MjFzBk+wnGjS4+PcG/CF39
MIv8G4a5JFiGLmOto8nmQubWv5xKQX8Pfq5JSOVGUK3eWuAVE9A2fgCI2HSRfm71
Rs/4Ushvjf+BwO6dHqdzLfLAPjneyL8Nnw3nCkvAweRP1KYKQqArzQlIfYdF/Osu
C17h8WFu0zIxKceW8Uc5SXUcg5X1qdha0fwZEganAGVjdae20lYQHdbtn3Mch+Vq
mQSamNivVmFdzU5N3wdLQNIqc73EFmlU9BOQu4GbB31cAIOH+6Ylt2t1LOoK1i6b
EtxavSZHBjsiZEzOR4RkZ+ZkCN3YNQKDOGO/wVBSPsuCavHAO+DRqZJx5ByJBkiw
Qbyqar83vgwnOUCBdyW08dPa1QQ7VsvtRuhVS93sX2KIkbvemAoZmawOdb+hLPeA
ZsBW5c4NEptKSpU2mUCpWMVFLyKJL3AWbE15ctogwacYXRCxVWt3SEOMqQD6y7V6
9uKmD09GsU5MmJtdQwtdOasmumkiqBJr+K8bFRvvSAlms8G4PEtoYabs/4nD6VA/
0xehnp1aun+X5gqmDVSTl2NuGMts2Scrcq+YlcrsfjDhVFlgvsuoo8zmUG0teMWT
PVMkIj8DrSkwY56Jkt7+KyEoM7ZYMxGoTnOJd7fftymvjQaoVcLBMUy8aLyy/+5+
dJiLDAHtHlmrNOr1ruLTLkD5ec3E3m3cmQa06t62LVsPh7wVSt+jUaE4o+dhhmZO
0Ff0FvnKwUB6bN/rlJaZAlwDAZdCNiyHtFyJyHghYc2zQsWgeYkN6r8B3wZ/xN/Q
uKthg45R02Jyq37hRSKz9eeLlWsg+O4Na5vERRtflF2eeLMV3601u8ZXaf+F0Fod
Su9btvJTAXtrTHgH5ZKiooh3hqZpdbY7PdmsFjaSmEX+ZE64Q0TJ+u1Cu039JJvw
/LExAbXj2LTd2oJeIX49eL7EPmwED3nD4QZ0E0RB0oCN18YVRq+gCAJe5gDZtt3o
GjIRpY+IcOmngfNogKGvZBvGsMVlHfoK9G/QeK9DwYtsY64H2eXp+x9ooLEaS3FK
JbfIJz9ISD4N/BKqoj72RRt7JreSwSpK6B7Gm+BPhxgwCrbGXEbIkag8EiFhemqG
oHuKfclElaqscaNTL8VKeT+RWNrJkknrcuVwq5QgA9nGVFQjbDwWcL9FQyCRqAJI
cN/1utU1ZP4KL6ssQWiKCIxpxmh18ubkpyBv3Ks4MDwwYfGSh/AHJUe6b1/6td5B
+r7YwRY1qnVPC+frPW3TeYuWDnI//wpcJ/wOvqFc8gkt38Rw5gebXAlELPGoOc0j
HpbfAlsn/x8Rn7kKeK6WpF5cmCyDmXAsb2GgmDM2fovFPFlMKzztaiYFPEwamTGR
z5zTlOST2TKVOZlsRO5io5Ng2G7hHtDJWtKRtiIbPdv5TPRJ677kqNC5k6jtUxcG
Z5XYjzS6aKc4xX9jd7UDH3I3F73tNEAmcrhDCE6ZHkMgrU+0OMDcakEI0yEcVAXu
wkKsZfddv0wBd+/KLu929cPXHbsjPCtkj/nxKtUkaa6rbXGnY2vQyZY5jC4Bdpi5
Bu8tfkobPjv5DzxjRbwCAZmfhNOjFuZ79no4ztQs7yFm0XlQ+ZjocWJeywpY9JbA
xe3wsCf8x5T+7ywO9uG8Kb7NuXAbLBnTVwrprmmMmdnJN2wvYDsqxgqsMjALs91G
gH4TCZsFqF8wlWasVhL7eBWkDtrCfcjFdampRhqRHPGYh3lVClV6eiey0GHcyKzk
tq95L3MCbjHabI5KthDZMMANH6OcCiNs7gUIR1Lzjd19QrMjA9z5++LF1dLl4VFN
PF5+XpLlcyq5Mlx+0M5unxfzbEIbhYEY9QQPOTGKr9nGEcyXe3Z+IWlzwiLMkcCg
6cwusGfzIiM98XO4YoqvnT9mLobYXjOOBs3atTNbJQ5fWqUZ0xG5YR49NPlAynPS
ZfvONigZGBGGGhsEtHs4SpgoIQiSeY5BXgc2K1anK4cOYOIHih+AYtZtw7f+WZOI
Caoa55yWWqizwBkVmYk8H8lkGBt0HfEiqsuk/E5PQBMaOTFkDI2GMKJJtizgfIkw
iX+M3sEJeBumWYSn4V/jSDlNxQVtscs6Bche7u9zyHtpkOBfYzdWAAxSVIbkWArE
ecd9Bk6RtDmT7WKvXIhd+oPYOsln848OuWYV1Bi5wSHsYm19A0e+9Ythlyv9x/bl
ou2lrPuRP85d+XORKc1K9fuIdJY1HA829XzPhC1RoyNhrLI1UGRJdhFlZUA2BQJN
9v/+KyffTYZlgzUIhFEDGx5tAVuvp4VZ7zvoKSjnXxqcAWBh//V2uyUI74YcKTz6
LjvKvlMvr5agJPNc2o/22Lyn5dky4JYNEfDHDH2hiTDsszMgpamisBKuWqbsXbap
p7kW+KJxB8Xb/4TQc4bRmM87YxHToh6x97iTXDXwzEts7YPn2uYZ3JvNmeM2UjE2
D+hSy8HunAVdkSI3eOvN+1QxHvR5Jlse81maxPFIY2ivkmJbf0JO6k9fWtk2aG1b
hIhFvEqvFN86eAm/GuWnRaB1R2bbcJf4jYvdXBkTcXVSKWdeEoJ7pMrIuRMmVbzA
/fRVKAmKYqNuCsuxz+o7pdi3u1EUUmPPfLLFPistn8+lN58IpX8H6b5O9l3fP5Cc
rMTmrcE4Fq0mD1A5FVLzYqw7ex0eCaNGviZJ0AE4/FVAWoIF8cMmbce3IR88hzeS
YfljqmFajTnV6ctNAR9xHhNszjtIYhTcQtio1SVOlUYMmnhFX5Hj4tzQX4BGGds3
vVrZMVbwA+CJIW/9zKR9MFHR1HkbMCSPTsMkORClzrnU3IsyIYNRkhWB1WlyUo1g
7le+77cMKvTmO9J1X6xlUxCZupOBywgm7aWGIY6k1bjkIB6pgfRtjyE/yL+cf3YK
/XdY9ZkPO/acEoLiivsGC/WgxSwx1yAXexTxYe8Z2p0SnOA/hR+MpfBtr4lMrlwA
QMvkdFzPINyQwzMG/WqklTlNfTWC2bEc7zR0bipIU0yiipmL5YEpj6/QtjMPuiMk
bm0G1O1VxNPnwfHSM1lPi0dAP9iTgeNJFszd5J2fPE+PrDF/QhUIJVQ+iOEouSxT
5ofSepSSlYoSEwsS6N1iYdYf48pmHeYY0RKppIXFNLXoFyO7kHMoWH8KR+pgBfy5
XGBqpCXV9HaJgepVXOM9rKJfElMPew/92RQzbvq+Z4v4IQEYwGH56w4pxuOs5l47
GvXpCtBd4OOijejGKfGzztyg2SbqxLGk61RNZO3lUbwYlAJfKdPcUYAC+RPpCDJ0
RW3aGcOAq3lAwK651ECd4yMa7UR0RmKziAH5TA9Qdn0e/MWGnnenzUHLRucuEP/z
Q6E+V0ikMTx58xJaDVWT60x5yy5GAlCGbwMsEQAY5ylQwLHazwOeKRWivAiv0/Pt
q4NBi/RfrUlKpujFBsJrGy8KsyZ+kcOL9BigKoS5DDTuMRtIGfXX3+wHthVCWFtd
hXrKNacjoKnMaIoo5U82V+YC8PU9Qm4Ji4hNewoKyJzxmlpt5+p7rKz+o5EXhXcf
39N8XNgjSNFTEoG7YAqrZrp/WYjNykscmj3TmAuKyh0FXYphh6T30GyQUKIakK5D
GU8Iq2kcf14ti1DIyjzZ9fLiZZdSstHOa4JcsJ1HYOeYmnkIWuH7+L+voep+IyvF
YeTTGq2FhhgwnjmyQD1oFbIb6WZ90v+5+0bkx/chUwoq0YshWGXuytAM0doBSAgk
0wGn7XP9JdeQdwVq5JwbjLke5mcK66QvEd6QMMvp3rHG/fUYkOgqhMY+NS+Yocyh
mUvk9Fr5MPadDk/p/2Pgc83yDwYFPfaVMRQ2LPjBEe1k0O+4FjzmTozoIUgJ7JF8
HZfZb/y3HPUaRHqOgLjzF+C+9zmsh1pePr9IKS7KiPny+K8EwbJfnroyUOnOwr3z
ioG3RhO9tzSWu8mKXTy/DDfoA3TTHHLkjxab5FoFL4I2Wzxo0a6/CpFCGezh4t5i
B0UVkduoGrrmopjWcG4QWDkNu+2FMu1nS4V5sh5v2DJPVLXD4f2gmZuTIRXhvAd3
Vr2woR5dGa71x/gOeH4PLkN7xiDVnpYBayZfn1QD6Nmrx+PpHWSPkOTQ0yT3HTce
3GlrFuLee0Uqo0H4/Kjstis6O8ZKU08ZpSDMsDkULOxonE/MQ17wZal2OT85BC9J
getgV5n4/S+CWK3ts2w+UUI45B0tKK8pHoTjvr/Wh1Ph6mE6uS6sS4h0s6XoTRGT
f7GsSJWwyAEn3oYztiNKqQkVaWQyKyPne6OOF5PbTopxTvCo/WAfndsg0sw19+ob
hE6l26oSgj8TJ5z+ZhfIExh7ZvRp6FNSE8A4RaIMxtAb1BpWxQLFzxMA4n8i8XOA
Q9FXsnzpw5FR/3wUGRbk3tvXJfAcI/US6YcS3OXYYoPFjE+T59EBpnGFDp0aWe6/
E48oxK90TvE828taD53o7n2jEv3E3xyOeN7x3qsHFfMr65I6n8MG2uP/eKucYI3V
F03RtTIC95LzEaNbVRXLOK4lMUoIvcM5D4xRyKgydWTZgrlU0Vv+t8erJ/gj0Qr6
TivrxOjH3ipkzXpgAkQcpG1ybQ2RGZF8flQ9Zrl4MekNV5OiaSfP0EMrzeZ9SreO
lqRnWwzA026mCB5iTXxHE0jAhlMxP6XXVHzXUon41dglYXz15gsM4qJSOHRpRDqu
ApG2w4/VJawpERwPHIUJtph7tANlspfGecyOWQ6floxnVIDf0JlXXID2mnouD29E
MV4mAv5sMRA0kNi9L8b33EQf/NKFGIyeErg4opxZfP0xFZZoAEWF0z6j/Kj2zU9H
8u6GZ/y8OaVfLaiHO3Zgh0SauCRkdKuF4FLqPmXSqrKSf0BUKpEwvKtyQr3IySVm
lcnrpR0bDrRk8HqlezbBqmxej3OlfVV5ic5lJEo1jKZrc9TVt74GjilZJUDvrEon
GY4EGKb7SR7iixRNthjXgOW94vEjnchZLNfa8D8ssPFdUYWYevEqGTifnDejNq+p
SLW16HZVG4bz6MV0NjlLgyfsUp50hrJM5++WkRjmtP487gs0qJJvViOfLkzOUe81
eWB7hHHQCQjcBAGow9dNY/3nTihIdfcMt4M7I5hr5J/F+gJWFAeHwKIWl5sBeNZN
KdxWSZsOhXCGrs5lil+eUsoVWoj/LE7K7v1nzZnmL9H6C5C1gakIf8rTPrfyOA6e
rwst04wX+Dl/eGB6/iJatS/U8fmZvLawuJWtimYrM19+/utnHeGP5JHFEWCnOIYh
6RiCfou6aQL9j2ykSoEjwXKBJIi8WdfqmnOcoxS+FnvDhOFXqJPWzf9Yu0Oiiy10
sK4qrwvesREcsLGhErguUVrxXcgEhSXTKVdsaO8luWAD53A8D23ILbpvYa+vK3Fy
QB9NmrWhVLTStMg5svPbtm95TkkKcCkm57hOk/sj5o8J+rV5Vb97QGBDiOBZfueW
Rmj9RD53clfaoNJD1NWyqWKq8weRMRGrjR0ZiX8Hlo96Xh/dV7eRqUfzNC/gB0JW
+qKp/hlco2CwTx/2P18xKA7Pejvi7ttOoi1HdIZ1RZ3sr0eihh4djRt6mC48nsRH
9Fo3Cs2eCKxln3XYxY3hqO5MICaIU13AS8/9HFMkVVU62rmzkB+JXEfRr0QRTp6S
on/jmYdaZmy/yGpm2YwEmHQo49m97a25mSN+3MWkrLX0G2KjF/Hd11eHCismi9+v
A35NTeEoTU1IYPWVBY2K7aG1fQy7XHc2USDBJ9zHIHHxEdtHiXE5DDFGpolo7nt9
zQ/aE+nQ+gQ5euCCZ52xT9/bGyjt00JxqGm0Wy33nNkoh784xZanYKcVD2NbcuH4
JwW5gJqxuL+/RTFPGUKKo/KRY4KSL0XaYpUo2guos8BSInZfC1TNJ/cugjwQ5QBh
CEga8HwedwTRPV4cpHQSM2FgKpdcdFmBWAhWBwEfWCYMc53gQf4vLEuFOshYXSyX
HwUteIHbNOuSmPj5rosPIqQN6smuJ8bdsj1Irh0zSq51ugV3+Bs77cFRFA81zr84
EkFB3ypkotxHl/Q2UKWv5RO5t10BD32jW/+eCJgEHQDApUs2MHWF5XqkbS+OQpQi
JHYE9yk4QP+5qITRFf8omlqGf+njNHm+ojrayYfBZeFyY2VYF0fKtK44ygU6J6/H
Vpx5f9hWa96ZHYyX5KAnSYk3Vvqy6SAct1nwqYyVtABwiF5ld/KljIJvvtbRqfH1
tcPmuKR8Si4bak35PNvtYiY/dB4EOUjiLXSChFl78lstnS6PBBNatErd++u5yDwd
1puaq3zr+m9tvCI4JP5yGsZ9HAMJRPxauQZOmki4wGbUQrBMd0WQXeH7Tv0X4aVO
r2vFU/cvGi/xJw/SkUFtasXmoIBaL0iMDlZjvobSeecTV79+bbJH2gDMkjI6H3Rc
bAOMeqVSQGSwCAoXltEVOUJFaCkJ/1u+4Yqj7L6sFF7dqIH139ul3zhcMMxwKhL+
FUtRYETdLPG66kJyryIscolT1egUwQH6nt2re0VtcAj5BOSH4Ptb3OynyYZLrnWR
5K+QCqKT/RER9K+CM4h0I8Rncl3/GsKvjddrKURwP/RDeUzed4i0U0QPHW/ugtKC
3DG66deYibvtOA052NIZaFUQgnEhi7KdtUnHmMJn23Hx8n2aEG4i/0Qc9u0g5R0j
hS8tQaJpB/UPRPFnLgksDIMYhfw5zVlMi6tM9ME8up/4kMliq0jLMUNu72Ed3ceN
u/1YwPocwOQmdNbb2P5jnjpDztEHGHgsi3ZXPKzFU/menhOi/kZ06pADoqWKFk6Q
OdeDcFlqxdc8MZIxscNuXsFHbEEvznm0SEKQQ3Jt2fNBIP+C9XdPyGevTH5b2kXg
7/L9OZ8OotzIUTEF1sQZW2WoTxyZcZB69OR4Sj4Kd6NQWurXHOIol7dIvjRgJJ49
nqC6bK5bSTQ4k3pJD6+N7MaoA2RZp2ooZy0nBxNpweZtQgAXDWIhSlwr5DmKNB6P
VpOeRglD364WOYjWKm2Dg9WTb7Pgwx1kUlGcR3RpJ2pB+PpA+NYOlfpjiIKJOjzE
lUdfzTRX4ziB+yrQJwAN+UFUUnuMr68byrnmqYU3QTNnJ7r92svR9RuxbZ3ogWAq
TxeR4RrQpKEUK3gkSRmRl3TVoFNPuM4yJEs+EbrbRNOJW8M+ZyVg7RRKnSMRT0bh
mCAHT8lzrvY2ROV0uFvAe8Ilcrye/YUADYppMaW0O69ZLjYWC5I0/7nw7nb3s+da
BdF2ZwcA7CdmhCB/zRlyQWc2+WcB/LmuX6TcB/bEB3eeSiOgJBGWKN2jiBEvtibM
mg2E46EumNivVmk7mlOPQ/K0a6M/WIDwSd5tyDYWpEAYPvedT1USwvvQDz5yPExY
oP7E2s2Z8UURtcTLC57sJq1jLrXjKbluMNYSJCM8dTFcfxlMckVrkp6dtufEVtFJ
J87cV44ccmw43oKbTXiPPfUj8cKRqbw7Z1KBWk+miKnTI/2Y2Up1gGBO154EsoRE
VJzMR6uIGxMpffteXaTMoY10cMxUkFP7xjPoRMm5duj/AYNjGBwYnxee6wEjfwW0
xg6L9TxkDe9MVp7O7g3EhEMVW4tORcq25QQUKnGb3Guk0kG7N40VcNLqPfiXSOBk
kSHkOGWRpSb4eheDd47yCTKdAsLZObVxlx4FrVc2uWM0yPic5Un6+xXqUujlT2xh
gZlFB45CMa7w2gqkZATef6enDIuVve6dqn7Q2T1NjBG4wImnQQbeuKMVirjob0WT
5LU94hCZLs9qvZbG2SfrOWCWFcvohOpeafJplWSrwm4pJS3jyhvRTYp/FWqXYEKg
sKAxUous5jCCqWz62/PEge1W73ZnIaNsficeWY0AGyutSxWxbgr3dOiXcJQr6xB7
RNwWHk58R3o9/V2ZyA12uZFtvp15+c+4jdWv8VJ5F3f4DRBgJvm8xurnBbsGIHbe
hnCjsYsIH6zCIs6ogs7+IUKJ+9WCxlbHAzMFfyKiTWtIk4Q/3HVKEWCn1IUeX396
SnoJRZrtHNClQFLXM8DWeg+8PBQVQ5LT+4jbBgPPoMXIkmoj0nfNbkPV18CoynqE
SGNopsbqXtE36xsqTagbAGPywzOEqA2bFSh7iRv+VPpdHwWWagGY24mOz4QGDplR
Qp/oxH5fxbM7M0QQxaXSxhbfaQ5/AsTWC24wSMYPidpG83YTt0FSLyXYnGpaE2cF
y1MDHrhYLZoU7en6gpGljZ1cB5mbwrU9+0AwkSJkO9xuLTtvtmKL5SLTPXKfx9mh
Q0vf3DkharS0MCwrgWp1X0Ya2pJ+7i+p1S42lkqtm2Bq+vvvdUkKERY43ho7DYxa
cprmEtVeUzh4rTdsWvQj6y6Skg3kixH7j5iJ0kkwiwkAQALQMt+Dys/yXB09VLAf
xtK9FwDs14s+PUjNnrNz6DJCmGlBBUeqtx7QWjwh6+NSjGoyJ4cV/jolC6m63vJA
5O3PSIn44Q7gH78Bz3H+HdwVk7kiD/1+Z2ET2XzKPElw79NVPaOg+VhAyy6A8fSw
o+uP6/yPMl99w7+7CGNTBD7kKXqF8djC7Tvpgjrf5Pb+UAf/GuVihadltrk/UleH
8bL+ZdqCW+lsW4mA3TzXgtZTogLLM57MFIPa5njGY8hyd7oCS54SRkez2fQIor9W
MhASkA5XLdbl08xc+9d5eZw3E5eCKihQNyQ5lI//Y1q6kvdqpG1Sqsav5WKlnnsW
kUiM7itb/zEqZZKHfnFomwgBjXle/rLW1vCeEraQlc8huhgrlQfEAhVd3gyMgk3W
YoVK0wTWTBFSiWqmysHurFcAYsmA5BFMqexeaq9Em5P0IKNzXWpaYAjwPJm75CqZ
ft7KrbqkJiCkH02q7GvSoWFwuZ89cS3TV+2B9cl3oqWDuXWXbmch0c1f0sPhrL5V
v/Hfho2m2jitDCtPoQEFqatAy9PHja8GNGFsRlwsdGSfyBfgL3E17fzqxKsxQKgr
G28d2J47VNsJovQ648wFSRbNQ2KeYkCpNywoUJL5CZkZ4YYmiCphlNQjr4KrNMLH
VsXBkZ+8mKX/3V+7HUUkOV1vPbY+ZrCX/kDSGjXnc2xODfawZJPqUa+vUVSOIbrQ
kpIBqK6EX4dwphcFnE8DfSbHKYeyDUQaTq6jK8L6NMwh5+A14iA7sOL3WucpuTwU
rKEsGpuOuD8KS7sZztNUg5cP9OClAZX+H/KGFSQBd9VC1DRCA1gDcADtaF8QIJKb
B+SCZKhbxTYXIH+ynfcMgLezVFmHWrE/d8SM2UGYZwTAHNILE+uvdfC5YcLKcRgk
VtGjlqs/az3sfdRp9EGpGo3cd2bClq/RSiFjyZa9FqLYKyfXNwOu/CFYFuVCVGtJ
psVt/SWY1ZC4TvtZbriTVyYZQfwxXA19EqW9u7+03cSMSLlPdyZJ88WxmWmO+dWQ
a3HzjABP3WMmlqZCkBqZ00KUcKao/lL1ZdqLBwH3dCx2TaPg2fry5EAGnzAF3NFh
clpEK9gWdv64mGrAo8XYfQ18FpqvM12RQoobvTsQq4Qw5ipo/IqE3Y8UUk7EOIQD
3iTidk9ezvlrct8cVcLYRJm/F0TriUuyY+GmwbhspAGT7wKIJvLGNJEFpsJkIGud
lavmE0pE+F80Jz23r0DZI0GdO9Y5zLQjr1lFGu+UoEjp/sQIWSjdv9jKrIOsNb1A
v2m32eNlPggAfJMYtmUXsI744pVggkg1ZpNZstqOJfM5aJ+GRwfBcUJ/F7hvNvq9
szRjCE7XBY7h5nZZdtxx0Y6tuttHV4IA20BH1e6wOLHpCdRawzpLqiZzwoTxiqv0
QPMu3spQEiSRPW9MR+flRTkt9ogy7Pmb3bGBSGR0PI5fMHXkNXFCceRP88RREHeR
tHxpIFbEX72pQHVO0/EmI0ZmPCnJE1AaZs4TNkNXKK/HV9oD8wphoFQJ+8ug326S
hQnkk8CXY8MtLdHdgFsIILYpFY3XoQ8V9n04RL8D7gVK2QeqJBl8bHMRwd/Jt6sC
igVm6d54a/vP9Fso91FBK/3RQNpyy2TR/XT5lAXws2Y56WLAtQGtojrkzl2HKkdu
FHDi+tu5BQAEedlmZO+AnlG8ctEhqYkZVFX/zY82snJqhbLaFO3YJHmiJnsOBvwx
XqIY2FUTrNuHl23ldjNQTIROzELn8sgtwoKEHEsaiMpIKwCJUzMQqPgVlYVEelCm
1gIs6SeOnv9jSDUWFDDK00LosF9Y4MIXZOm5dp97mX3/5EjawXEmjuR0bzhBDmcX
NqWO9MYDASf77bMRJJ3e19DCz7eEnDtQrd6DmXbaH3DR0+EUxGvpk9GdNSrRcahl
3SNgBQNO3/xJ2fa2tF31sLRA2OXYPug4mg9q5K0ZAGYQYokHWc5mo+BPud0GIRNS
bpSgEkOoic2Oc1yO8IwMFC0NFik67JlG6qVpx9UzCvX7+aChcy8BW/2urIGk7sGS
UChMcT/9Ba0d1nk442mdQgEDOtJcGgMOy+BF3MNVsFS3nfDqZl9OXrW9Ez0liLkp
+LDzVbS/C2kW57KMgY2HE2L49UoJhme0uZ1DGqZYRfuZKdFulGDziZ3q126geu96
qBuANlj01ulqYqDL0S7z07NdXOJqvR41eqKEMIczYW6NnBkwa1E4uoIYnXNde6x8
uycIwKoH5PDEbTt+FXh+gvZLIZCbUs3hWn4HgcORHUANyQFPfX9g9wG5sdyEEb1w
0KmyI6yQ9MvAJPkT0YISre9EREw3/E/9NLBCEzCqOFMr/AZD1xVDUA38zthoQLjj
i/7EEyfp/OMwMn4CfPJEQ9B6X7O5M9KFEgW8rZdwhuLAWZkz3VobU9i4GgzZExIP
U4uJ0BvylalTq1mVpENPMyzyUNoWihtNgJcZs+rohIzOQQP/32S5Jo71xlj+Q1gF
KaRQkcYsKkUeJBg/RXxMzHsPrnR2TUuEUvaIRvB+ZQkbuW2vz8KQu1xkgZ8CwGU3
eEjzN+VOv4HA8ooAnrNEt5nmQFFsMNysjwBWNTRAma/PRupV955Us5alVM0rfdv7
1mnmQunUaWVUo0zGm+GoCw06lm54dCAjcPnkO0glECqGxUT8hRCCsvKeKzPtkq8f
4jtGu99jPO6Q9ZubH7nzYi/fdQUetZWMBMwFwAaHXg5vadC0NxQozSViOhgmISaM
0d95dNLoQ5fX4kRICc2crcsYGGlrHMXv1aYarZwRzfP8aaJgwjaQEMDcI3bEClV2
M7Vy+fH+q2Khw+pJkEI+GIFMQqLuwCuDGv3uxe2aQpGHBaqHztbwcWddH5Q0I9qR
WwYPPtAPORkHsf6eJi+AkRV+6UOqOzIdtmFKxV5uoK4WyGNSxqlwruvsJzdgSZwW
xgqnNJTSNbvENe6lvzMKemCyxrh1VAniDjS/WS6MvKk70BFSpw0NnUgRSpNT0yQW
UuBqVBfTiwz6BqcjgoS+JJbJN1jri1NcGMvjaUewXwCn5iSxFrKM54oFn//ynoSw
s6bEutgQFfeueqdWPA3BasyH/1tIRQpAq10IBI5cJ9vBmbXI5zqtkhycWpFgmVzp
Cin+PuxVCy6u9NJHs0UEYaFJFI7q0lhPgRmOj7GlKFTfGPYXTf0hgTzk2XqBwWW0
hkG1yhga/w3eNnnHCvBeqCLwzerJl0oYBvjvW4Wb7LiOn5dApMIeRN5HahtP2nUf
CbN1ca+P4eIWi4Jz5OKxQXYqKvm9MK5MJQKyTDqvKMVHzdA9nwA3Sqe4k91FhxES
K3iM+Ut3B5g/KHmAiBo8ORbcTQmiLwB4DAC4dpljvhHbamTpEeHa7cTiTDkTSUdJ
giKcy/fhGFQ/ez+Gg62M4EgKKzFBzj5wgEjSXUI2gZ6xXI4iAgtDChsdMx87vh3g
Es+J8POE9IepAaGLYNqy2/YAUEs0rsypN+aRLq4pr3ZmIrq1t2GKBlcidcLPPj9i
HEVF6cNf0BismT7FSI4VE+VJZa5tU0kq/bK05v2LHezmiV1sVEXAWbmrGDhWr/HU
3uOcZ4+ePQHRD/eXUhpdl13RHawetKprR0HiF2OYOayTeJjDLKqjvf4mGyRO96gb
bXlnGQZuJj58aSz05p59YB/FTADnMkGzBkGLyDDzxGcr814kYTwxT4zYqDwzoT9V
rAAsJ91Lq/0qFWLDduRI5Npq5GxeRbaEkci+k82pBxThH1xx5oUKLtQfmtXgGpRR
XKerqq59h/LDaRfFFdIQK2bewMzjIl+RmImmrGU50qqtI/xMc1SLO7RXSVJi46t4
vw0gqElg4n7/zdb5viEBUuzdYSWpk6Oq5W5X7KETr3CNiE3w4lAjJNIJ1fex/Nra
95VXMnF+C1LLkZZqpLlA1WsqRLQi89nKNJ5yjp+iOe9DQCy97A3VpSS0O7NI6M4s
HQjK39HBDGUWQRMUnKhDJeeAN/guBozSOc0N7aY6FvMEKJ4IYoWteV5njfIQy4yq
7N/E9gZ9MivPQ7r1ZLVtmPDrlmH7PBCEerGcv3eujw/idZ5NS45lacJlFyewl9tA
F2ZFQ+N7BpTpW/WV0SpgfVlwyW2+P3gUcHnKTivkGyfJ/tSqZGdvdcFFR/mYGrkF
1KwDajUi/pTm4r1pnyIySxgZrSM0IgDJMQM+8XfBRPPmaoNUUqcglqf9+qYl6Sgx
CQH1eO/SxxHnxHEJqWl32SSAoAEt8/Vf+MGklY8DTi0J4LeCheDtirSu0IkIC4W7
ZHX555HVdzSeZYIRZDorjxvwyGYbIUOKS7v9BTI7t6r/tqUYWjhfwJPRRFecmGZY
XL9uEEtzi5qWC8z1WUE045fHx1nnEFt1OoQ6t3teGfa2pnC22dJnyx6uI9QJReBy
jtANLVA8HzVzBX5oekP7iZN6bMO7bOIXVNQQrKsRZvf6a+Hhh9MZp99B28+BJuJg
tWmtoW86OaEuM/STYxu/k+HUKUpwPYwyvF2VeFvxFdtbQzml/1q9xV1kARLwz/Zf
3Z+ncJMCNi102r8akk3JJrQ2Dq6/pnH+tV5buJQ5P8aTiS1kw1x/jR2n3W12acS5
d/jtOrQXiE7K9n7rbakrRVlBtRJdrQ3+bPae7n9tSPgGQS2ANMezr3qmXqXiBwEA
F93IlW7hrJXPNHiUq+NZqMOmnJWJ1J9Eacjm5I3+G9nnmr6b7R1UlhC86H7XQJFp
ueMucqYPIup87kEmdOHuQ1oS67BPN//Vfiu+UgFP3//KoNrb5NYps+RycTtft1vG
OUnAZVFshBP5WlFGTaboENXV4vK+O0q3ZyYzvKCJvcNgUOCWGleDhdy1IFQJ+7OD
PvquaCvUXzT61SCoSRPDqnwo/Opp9+Z1758TCdMEpVD3i+jKiq8hRWSsabhNfM5d
v0mDmwaeORxD9ybL9/Bc62ktsgwxRDOmWohixISdt+vQ6WpwDZ1OS9cTxn7qQvLK
drkRcsaFaLO14GRyZspOo46+28q7aM354iv0dylwbMEZLqS+3J3Ur2yeSAr6oaCA
KnPA4cu/v24WkC7Sz8sfAc5ApsKuj2WAIV6dNWrxMShYOUSHwcxkKERtoRb4EYQs
kv+nuY5GiRCcdhxFNXuCwHjX4BwEbYNJZFPBL6PlcbtebMKrTqFN0g3MTz1Zr2Re
X+dAFyqgrJ0th6P039ZIzwSrB1zU3LnSXQ2JGq6SC9tMoz90EW1LktN579M8VBb6
lNbTWiz+tDZg3ic6GBkkj40CdnRajrK4fvkP8uJ8MZ9C7IraEVnRXhT2J0ogZ80f
tCHdzWU0C6bBzZndxNOUX+yoWhVfl0nQ3Q9MgF6UIy/2rfNrCgWb6NMHzgPSiOSx
o7AJY0R2F9TtpzJ2KJhCFCMjP4uNxbMNbw4ELWb+N+IbLWEel8kbWeJbTTftmwrM
T1O0heqdhXoaqoGxEiZJ4Gv0EVjhVFQtytEdxsE8RDQoW18tjgi9cN9HnXbOL0Cm
PwVeey3NT/cwwrwhvag2FbsiIn4xNsB+BkzwhWdwgmkDGYD0ogYwf1DNf9vjUsn0
asg1X+q0AzGmjXtyKcByFCjyOaBthQ+azOhQBb3CHqSxx0Q4HItpW5ZxJN01UFIl
Vax+Q5/JgXi6B7C3VkCkrsbUJRLXgAzkOd90+V1wxAqhQOC/4xbCIsNzJbx+Sqxa
kUFN5mBeoQRc/mWFVEiJ5t1ND7OayCeALVXelcfN3PtVwoPUH7+qU6ffZz0ZIdxn
k6530jjV4SWF0i0JbV4JdmJPsBRmb13aDJXp8znw1sB/lfrUPXu4Zamygv8vf01b
+y6cLZSPKKhdolwD10DxTqEv3krRCXu+dWPMhtHbi9IPs5tLsaesBNslxvLJoLOV
8cU9U6JmQOnbUQgtLx8IBs8w4JcMT4T9/Et7iP3C0t9CzLQkb5tlqZap7VjpgtnN
bmAkfrOT+PMrxblp6QrLQyUwEkwVt+CS2kYE3t7v6vIq9CMwqZrG11gym6i877/B
MqzpHzHMLjiH25jNfTNF/L/qAEpgm5B+ivFWkC2OhG9k/4zFU3O3lxWOpGRDueMk
SviIxO91Xia7TYSbkyXhDa/28jXm8CQHEBUAlu7oA7ZiDB2SdaZUrdFALUe5WHQS
32fZdfZ6cr+FK4gXslapfdKBCqDtfSKsVYw63dUy6hbebUthsxBoe7n960hxTgH3
u2C094LaOk1LRN+6bzI1D+3KxOoBNWTWRPDAtl9E5X4wMj12AjQ2qOhPTdYNjKD4
3HIwBkcUp9aFpZE0yTJiz6L7tKBbICp/cEb33KJP3DLZ8cre9vTsuvqZ7yw8l4yQ
cfPWZnQuCLWfFqZKpcRBBNZQoqd5X7PTkywcCNBMPXnddCzHCANx5g3+UzfbzfQl
VwNUw3yDPFdT4L6YVwStxFgu1fd/b6S2xheKclWjNqFPsYVoWdD9Wnn/JzbbkMnB
rVDl0dFs7ISvHeOvLulCrXEWn4IRA2uKs3V8w1/3s5QezvlGvAWFOWc/++w8i+wM
iVQ67JaHCnlnkovlk3PqX4Evh1vK+uSm4XzCesNzGSQyT9IoSaHyKJpBL+0ts21l
p5VSMaxlojpRXBq7yJBoUxW7eN9bYV/4sMxNYqZFctNP3qi0rQ2hoFZK0Gim7Lut
gfCVvbj6FUg1j9jyXC0PlXMgFaD1UaXs5kHhsVXa1T72i5ghS+f+IARlfgBfB6dR
gd3k1BmQntlnwAUhXH3RL27go66vnZtMd/tA9mvvjilu7dlPotEJ8SKD2QkGxmoQ
1HM6wv/g5W4EX/GAKtk8L8p8tdA77cQfzBGAfYEoOqwhM+rcW0CL6hw6YLRgBw7O
OpY1OP9TGGV/LsNXajDmctVfOkyugvidgMFW0oMP4Cnt7RiKuFJPE4MpyTyNPu4n
VjP9PXRHtgSoAPuR8IbjZoKsq1ov2dOWQmMKUu6shHeT1gLEo2oLVtjWWYMcSzWE
Pa9ykrNAU3rhu9cXQXhbYMYOGuLdbCCepOHlo04XR2h8ArNTOLarShfjkZmRILxi
AkE4F0EjSEZEuwHfbONfbm5IMFDJn0XGXxYZJ3O/d5mmfJtkuWOApnAhQdDowJeI
/FETELVhfG1FoY2Wpw/hp91utejF1NPxW/RLnYr2ZFgtWX9DlFPeQPhH/dL1REYx
q64CwpoDUvFe2q4xv1O+FL9JJ1wS/z9cZbyKE7k+dSM6Dbh2gDNSGx5sWhuHr13S
wEJm8oHjwJBz5sC3suAfMqc4QUbPhEcMWjAyGx1ihMhGISxKUoihciaJV/eMc+5o
QU3QZSYgsvrMWfIJ8hG9PZ8G2k3zyrac9QBlgRoSGwklt4O5HXfeJemDw+3yVzj6
3MwgHT9IR14bMe/8YhNJT37pKXBlGG3Y4YNJhdV1hjD9XCJRad59R+osWhyLwyrC
zgHCUSDm1EBoeXE/BNAvCfNhA3tT/wZTzGfhskRhpEMvryO8gi5SvH9dxvoxpeQA
8I+PFhCka841UFjWaGdJHTlD0+6ZGfFtwIiO/odNtFnVwYQoMaZd3ggRxaF7Fw8A
ULXISaCuw84xtVYtpa6I33EciRStfXfOxTabMDLslz9l6LHVTk0efh14t2Ybul5p
dOcIkZXiGI1e0jkYZ5sdTItkD8CTfi13WMT4itEoQnVkrZ0IJTtKHonEW/i2wjf9
rHaRYh464L3hobjdvMKQSimMUQzO2m9gJf7n+4/aZI+dYQftkC95otPy2ZvEBCS9
kv+tgoDwT6qvClbTpl9skvEIo3s1aDiXMx2hc+z3FnTqQMDkBXE07EBpmlZWWCHz
QBdBrirwRzpmI5nGaxD/YM1i+PEpyBXGo8nJxkLNfgYkfyRNa5F4DYo8FWQnSdwE
+56Y08kxEzl2SIwNYJWz6iuucJ0Hy8Adaeg3mSJVQZ1T2Ef99SViyZ9gXAMVPxLl
s3yWvxcRGY1ks51jeGBtDsHEpuS4HDZdAGOyNEv7mupxlsraGnQsLOsITrUhq94A
aw0j7fSLt+z3lmq7j7oJcymNDDym+cQ+VoITz/yVzaTX4FlOZl1up6NFuNCSD1HK
/WipFR7gTjdueKK7iq3uh0aBbeTWwK6XG9vyIJRu8B4PrGO08B/YgzD2zqOkUOFL
q07c93NrHVGcosRjvHy6YuesnzXof/pdwTagMKw4rfX4kRd4w8TXROFGbl5Z+8Pd
78+kfc8dTWBDfswPHdN70CBBTvVEWJKS//zVGK8s/R4XDfx/7R/xENIwQZBQoZes
PS20M+rHZI1iQARq3AozbM2pVaneraaXbZHw9xPKKO5B2382oGbOaY01mxt6o5E6
xKqHWOfwev//qil0gSyNx8RprREwrOTAoCCvqwuHV7+hvmPKjhgOJDpV5FtKz25/
PCNklrkEA5oOhas/O/kicues3ES+XsSYKSKGhmowFfoJu1mDaDqHxV5quAyNwbqE
0tCuasQU5ttPyZMMJstP2JZAr2Xv/J3YoozxYwywSRGvDqNDj9SUJZbjnPpeC1VM
GIRBdzfGwCQPoNxOgJ0MKbvfjzrtcRc4XOF1B4DKN0wPXeoShCeLck3VlnuS5wsj
hWlV/Ys5AgJMF69w5q9q7Cb82eErSvWEvipvMppkVyLwLFmmIPXE8GQbs612jZTj
94LFAwztlOE65ZE74/wRz+RAihgeLvxgtvl/0ptX64k6XM9Pltts9CtAg2Red640
3A4BcZOCgyYV9cGKgEeJDIV908nOzWomrAlC7QwpiEteCLIAKykL1Fs8tUhz+KDq
67qAu4vYzih2r/AfNf846Je7sFY6yiB5CoAwEWczBoha47Td0RlRg6ynpXXyrHwY
/S+Ez3nJ4BD8sMHF1TMcrcAYJXMUCZvgynBIAF199HZ91f3k/XbWhPgllAeInp2T
mjSs7AfyTOgW6v3/KTnDOFxvqhJMEm+E1+1wPn28OjWHvOAPhECaevKeL6v5PPNp
jQ3hLz0Mq4c5dMr31gdFDA91DQAaVu8JnwLAIFIEtOlLnGPA03cqSUZ25sZrfdXB
86tROc8vqQB2h9EUl0kYtwaOENHDjL1wLGIdkkdk6T5H1U1QmskHRYNMx4+Zuesl
tGFFUBzEHcIJjaIn7FMuiFvYNlYNZKC22V39xwh3rhgLLlmSpnh2SUe8udCAapXx
zXbAMqoCdj8Z/62VLUINlN0Pe+zt9Q8RjElJPL4quaj+Wjf2+pW2JVojGOsDDN9Z
O3GpQssS/R9suq/DHogHMe1bh6UW7k0c4vwA7Rm3UZwde7E3NwdwPpOjddoT2Jf/
sb1SRIAsrGEcf0RfPVEGiaaYIXOwjW9caZt5bf1eEVl1ivJa/oplBWudpsFztxNk
k4fxmHMcSuVcVKoU8N2AIFaCwf2Za6aj03g6e+f1CH3cPH65AjwhSZ4ciY4LU2y1
O3a/m/x5ZPpqqqm9FF1i+3SBcotwYdivhr3lJdB4RnjcnqhBTRkv8ZRj1nR5+SOq
AVBVnILfrSvVor8ohXAyavHpl3/JE6loLIz7DMq0SoQ2cp8J7NOHYdnUwbGMx2WF
HbpghREWm0HBiJscKMv1w+An8M217vIq+trEJiENzIsSSp8i0k9r8Npw1FBRYgwN
xPm9ki5rAFY3BxHWLDI+Pna7CbNgZEZnfbdO/tAVldgC7FiBdkkVQ7AFVRpJj7BN
aqMsRE3rx47lK9SGBjdIU4MCbLlKKZTfCuTf/WjmMHWIPR5aYPOVk+ftu1OjIhQv
F5lC5ztMXREPgt2kaXr9cysNfYcsIOAviJTiFrNAhrvrwu3pjg1uWVPX67uSYS7x
tYziY4HzsVJl9d1pSlJv+PZXG/PAxgu5fRpug5eY+ajEchx2cI6a5zGyKxEfiZkI
YRnQDiR5dJ7gttbdomtoBmdW8XNVjVVhPum4bjK7Inb0PHcCbkkpwFHgFgZsDr77
VYGd9gnBFOTtXEAtKUSkpcZgTMPYiIgM2BZK5cDE2wquAoPvUFIzB9i3w+5oMuI0
KB+9iWiMXaQmpVtVuaHRScnHbIYsaoZE9KzeeVtNJ/rV2BGCJ1gzwSdlWGM5ABRM
2g6kGhXLpsP8fhZU5tIhgt4XmKp16zv1YajUdYZSGFJdVyAnF9pS9uWFZeG/lnm9
LBBqKcJzbMvREVVY/o6NykMnC1AehxqJnU6iz8jSRQ46WuCmbL7izaycbOOShbbz
JgGwG88K8y4fg9sUoNgrfoVnTTpnXbi3XGMIs56uCxQryBhYwH6sAatEDksKxo96
kRT3GBxp8PsqXcJbAL/QdoBuPZms4eYgY34z58mISkaFyppQW3By4AZIQX0UQdni
pB8SwYNCITNLdsrZyOAj1jyuoM2e7bGMBZYSttrncouwfsM4SZPvG0SZO4c2CIVX
EQ2tE+wuPnCMzrHczI/1B6O5n3ieHb2JyaEKzIwm9hA1n3LAg7N3TLu9Hbc9u73j
3wW7S+zFjwYvSmNJvd+n+L29rJA2bYZx49s93alcU4OvBABtBuO+jupW9OE43OS6
LOUHr0Vgo/bOMi1/1x4ms2Ly8+M8DNrkPJdOMpLtBgMv36lgSBO8dVnFAR6uCqOV
H220YmDWJMermQfS0h3kfdCZpmZf40m/FZBGwkjGLIauCeI7/NXoxryYG1DZ/k+Q
lHbiWckDspwC/yaevdnLofbTjsx+3TEkIRUf3YC/oFDBJjDrjQhrbx5irBc05E4I
aPe6u9DHnASWuXT541i3qC0RaKi6SX84oJQ9e5nYb44K79YexjrUI1d1VnmO/rnm
a9g+N2itJMrpAPabCvyx8rq7N24DPEAnnnLoP4EH/OD/jNre0HYOeprX5QfuZjv2
cGrI520Nv6NsNp/SqDeNcYyIk7qmqv0FRcM7/unn5glcwSbMMi3fBgNUKpu8sA27
6mTaHNVaNU7XUG0sek4giPfvC49aV39+y6wB0IS8+qqg1KvQtUyqyaO2YFCTDWKI
VQ+7kAf10SQm9Yck01LKEQSPLiLQFJZaiHGF2/dWDFdc3GBJftor62nugNO80YeB
CpjmmN0SKPZsrpR9aqSF8AF4FkgXSJeF1Q2RN5QB8LZu/o7bn+J8hA2K/qQUagM/
t1xLwC6cceA1JkSAI62HC3mqf1i6a/eEl8UvO1CZsAorojZfVCy738XIxntyEHLD
GVDHqrf0kL8WkYP++NVetrd+cZxj71pX58U11z4G09H9Mtwdg5VfkJQdhplTlepL
98OL7m6PjMNXmc9s1fxpWqkaGf8aOK2o+gNU9or69SpzFtVl4lgD7ZPfxD4VdHJN
z5qpiRG8qgVbxcBs9FLNojTFQcw54W6licmOCI20bq3SWtXiBAhiOB4OiJMhqt3C
GoGa+L8vvlzYTmSsnu4kIFdc67UTZ1nPLCc9Ce/pe505MG58nAhkvYd4mKvZSWuE
G7iLJIsvlJomTeHsbhKHgLiGWR9ldEisqll332sWylc9l7EtIsNuHk8T+zAjjgxs
WPKFQrIbSy83WnsgTrGCwTw0SPBqI4P/CYFDWhAQFUt7vgEnM51EVpbRX8lOwNOA
Jh43UoFBSK1/DG8hGFb4m9OWFJCrMjU4fE5T1WXDOosElXvsH0q0q+SNnGiG3sSY
2ukWTIQGen3BlzODPbngAcO3TXRfMPVVZ0aXYfxo4Z7wICMuNcJBu3OiMD+ONXxE
YSn/W8XVQ4Qjd8PL4hYZOFWf4y1fLv/Q178uanIdtpLMfJZ+67m+jDblYwbiM9sm
rDBEraJLB+Bd5E+VGwQAWa3nO3qeRR3vSBiWSNrSngsQD4rzuIkXxpqJWs0v06T4
JRk86NgNuTqozW2nGSlo/9sN+UnAgta1kkSJ9NQT6Ovx9JF7cFoEyTo8qBmcBVJQ
lTFRPa1MPRzeRMRCzjvS+W7WtPhZlvQJMakObsg+pa9TFO5Iv26AHfXA8/28vX0H
UHjEc+2tBwWMsNJdvKjGNBnU33gJZuokpSZTMjZx6ZxvoHycKeBhyi1yYAuitvVz
lLlqMwxj5V9zfY08mglYSJ0cRLHG497Ns1aFR5voa8G5upPPhAgDcAWl086qXDyZ
BS1jw1fthK81kPNiZlGudfrj8UanJKNqlWRI05gHxg5MlLO2yE533UZuFyeefxP0
cdbgI+GJVtEZhEUn1ctRKy/yFBIWMK2tAf+q+N5iTVtSdXdG2x+LzlfhtDybZLAD
EiXuTmWE2kY6UyjgUnRzkH59PVorlZGb1FXm9EzR51kNcUMKo8Nu/DSq3eamyQBm
nwYFmg0+arXKILEGL+Bug+50zgJw+V+1YFphgC+cfWDBAqQlwnsBoLvkEGYGT+Xk
ztcMzztfP/b7i5CuHr1a2nzDQZp0NKjq+g1g6T732Gy1+1ly1Gsq04q//h6AIPu0
YEWwbjezxw/FU1YnL/NTwqEJVM2nJLR083DkXC4suiFir4HN5lhrxHwejOX5qNeb
um8bH+Oaxvd2aS/eRw5bluOa4xAc3FseBZDcacRFa8rRAhnH7q40jqCM0s3l3Sw3
v077bGPQB99acdn60sdHmngEwDMbZiHSeRJqEWZv52YNkmzh7Y9eWxSwwqBQveXf
wKZ1blKkX1gPOMUrnizZTvP9AP363omWQu2+GyVD13gqFgazFnr88jlzwd8Maxlt
VVRXcYZ0sINWB9OwE7X4RndpXqXLMrjr42IUujPwSEuBrS5Hvu19ZD+2p1eGrD8b
Q+swgsxatEnjJzaocnpRuugmnhnUd5DN7zKgx8PnIiftT+e4zRWeluK+8Jv4MeWJ
MrKuCvc3xRKC7wFogPxUfuZ1AlLYP98wxJPO3906uOkx3Ji/fc4Klf1JdKGKR1G+
3rr8nzJpJB5VNC5MaZTNLn2qiucpKfpXWoQqRLbOS4JXbQ8iK8DoImKjIeCnp/kw
lzOfIWAC5VLC944rBK3zGgCG1zuqBwxtxQYBWaG078NwWtCm/aEbMPMkfULueaYA
A3dM7TaBWLONkU5DXINnMb6Ak7xg4e35ie97YE2VdHC54+pKkLi+UUA5rElnGHEH
13G4Xd7w+gE5ejGvsbhSpEDe7EF6/xS36OjDuSyeIHfERRPNJeRRejB7p2MKEfC8
PeRqYCibjKRZuMTBzTMZEm4z+dDuVqUrA34KM6l73GEcn4OIZFtNVrBBZK4lYJzu
lB23Ocua/SvxOky5/G5Z1ZdeKNTgdl+vhfUyCYlNT5YHGl7oNQPig0JJ2yrRHQqY
4b8MPynTWHXMi0YexuJ1uzsdKUbNbmeWBVwhxNGxVBLUIVsIUzFOaaOV2heYJaC+
sNaj9hz6NnffM/UM+vSkuCCVTLze1rHsI27eO3kTIC/MuGF4j6Tg3rhm9EgNQzN3
+q9FvW6Cy58MXqeEu2b8fRH1N37r+BN5zbNGxHy/GIemUS6P7QqnmTL+yEQYJY+R
/aSxXFVr4jD9hReNsZiQ+xSZXn/vJAt0FX6tMv9742erzQGV6F1UrmGSiheCYxNr
xaDSRh5kaqDQQxy+ie+p+vl/aC7x8tksD0AkLS1dhr631jLb0M9rJ2L7PABkryyF
cj/g7+PDTV+VgP/EiWeV99fOyg5Hek6Mdnurg4BdB3AvJcSTuP9ueqY49PPvFwFN
S9k+9acFxSbk52K+z66uIztyMpRfIKtxXidHYIKQKXZcbNd+2SeFI5dmyjXKpUa+
0bNzhCVukjNK94j5L3NQRuXfyv9wmpPP4I2DDb6X+gHLBIgXcCCdKlNtV5R8s40I
jcJ6p3L8fa2hv0pu6A0R4KFWjWLZhrFgfVIKH/5z1OnEAw8EsVE6vemjN+RobNr8
X3F0B4yUaWFZqhNQJ2Xn7FDgl+wraWwSeeixvUtcbg0GO3nhmN8jhY3k19yWZGVe
Qoemb6ApzG3RihvYlLFSV6sg+ugzImj4bFgyxWByddub93QD6CDFebZsKZr7F87K
SBaFOYjjUGhNUjGOUtqYllE65v1L2U7bN9gPFZ2H6KVX/2zAaYa1RnxwT+8DoshS
DWNHlf1cGLJ0uMbv+RTPYla/8Qg7+FdUcq2bvsbC2KhbAzBLLy0Ja/LKTvJ5v3XW
/hcweaw46O1xKhONRwq1S9q+a3an/kcCVvTsmD0mSrqNWNUSavy3pyPO3khLK10B
/PG8w2rhuN6tRW2eUaEBNWLwvhksNuVBUSzVXRcCBQsQavsvFEVQDWs1kW4aMQNQ
Jtd8mRAN0j+Q8c0nNnLfby3X9ZL6Zp2R/aA1pKSH0aLWXqK5JRi+24PDmRT/KcZn
51nox9iMzKRswBeDEysvu8MfXKjGStgFu+jwJ6v4Gj4UYqNqRsQTU0PSVo5kqnwa
mP9kM0Rv/nwslj9CxvdeL2dNqIfYPXCANJJV/Q5p2TZjq8ECqSSbHe+hdyr+zVaD
ETbaI6byl1PphVaZmVopujYj8wYrasx2g5FRxgYcx6NG7rUwkNCZfNxS3Ipgdpc9
lYeIOmNAJoTzfHUi2p1QHi1vhM0VA50fIiF3HMu0i3/zboTu8+1C/gId+zrnWOdC
nwL1kJPJbFdoA9Mk5fxwXMVso2b0sOf1hkBRSBHEYRWObFAokORcLbNQhlML3yOx
T4dlq/LBjXKa4DBWK5P8kQ+Uc+kq02+o1ddI64lA1XGZ4MaasI8rc5vZwarLA8QG
i5HOrQfrYrJexnwY7H4QtSG2KC77J9UTZIwlUuf5214R+v2gSxVjRXHm0dvOpqDQ
gT1qrLtAbOSspEGrIKVWRWjMzyzk0d7c6DdxSe73FYpSPqsvZ99dH0/Z5UWul3Fk
E7+17bKHtGWcQh9HIBwGBHYFANfZLJXtSYxNKVmHaj6zU1HzsrRykkXU+Fs9nja/
CzzxMov2ZNNq/LtPLaKE8bGj9v8iNNwv5BrQKZZi5QTBGNNYbPe84Oy+ZYTaExJh
fUFCgCf9T7hAhJb8ioS3CLZ4gfaBbW+xRTEeMLrdVQPc2o619zDcq3WnpDeHESJ1
IP9dkAoalbTLEtjodQjeedFjGmbIjnkzv/8XIFjgmTZfb9OpPpzWMCcd5ZNZ1U3v
pAIO+pHEsy1rNGPGZUD8qy20jcuc3Row/NNMgz7ib5vl2O0o14byWX/w2sipXBJp
Y5PoyKn/mamCgZhD2e+3icC06mIqIzgWHX6BtL3N1NG99jrEkU7lt/L54PadXx2p
g3jmUa/If46il/AxmfnxQingvGDe8hOdSyoJuuOzM3Qn4+MRSWq9ELVEqVc95y88
s+c+eKdkL9E3SoGqRrarM3eoLP7qbbzLaICUrS1u5AK1kNH/Tgupy/3Ufs8Mjjfb
IcXJALHS/cBWK8BeTAwui6M2vIXBgxMg7vd5gAdR95L3FMB4xJRBC6g/EeSY8LFb
87Iw94sNMjxbXTpTpFNkzap2AUBRGZST1gS/UCehBbqjcrQap5c8I8ux2HVNhMDm
AZQFOGfOEZnl4D8J2QMaT57HvUmH1h9QebrWNhnzVxF1m60eEFVSCfDQ/H+GsQv9
1gnYmz3vYDPzNZRzYQPl3dln6n6xugE9aMgCS0FxN703S9HYzzrjkjlUZFHTZSN+
z1oepmCNV1GSKa23tB6QZk06h2qeaIZWChHc87QGmjl/unTnUPBSGqiLJu1cw9Xo
RH+z6RUyAgxM8iDWFk5Cjr2Ra5Wc3n/fX53FgUoHjb8dnradhKKlsycl8MzDe9wQ
yTNJD9JLgAgGwt+CB9WIjaBEmn8odKVszR4eQBQv6w0UJHAEguZHdMKOyYitdz9d
FiIE1K7CGvF8GTrz12C+3JBfV1vbaAcji42yqkA5KcQvN6pAkWqlZV8tlhlNFrUW
X6PG16l1ZdfQBAHDLSqGOXEFagT7rIEeBmiODaFBXpOcK7H4zhWLeF8+iNsb2lH6
OXExC2KPei2WoH/lxtraM0oSLphBDBVjfDIInpczFSuoRa0QP7F9r6VatgpX+qw8
noB64neTTkB6vzy/41Il5VRGJFgrau06xpUV/C4IH4+vbwsXZuP0EbTf2dMXvS/I
9V+u7o+XkGpcon+6Yoy+dpZrp210E77R9aT63EnnkPaAyynUW0D9t1QHIdnGkWJf
ISCZnXBUWKpAGbmQ5NK6mZXgRnRMz1s+pZLGIFeM1jEyxU27/pbmDISs+ODDh9Vl
5PtcLxSteu+//9Z+ushDGfKhUCiWhYwYySSsmTXiNNRIfrt9qzHZUwhNhaIwwHgE
Tv9jj0kMKRH7CeAAL3uEL2WT+jRK28fYMZxNQSv0PDNouti/gYnhjWTPuMuwm7F/
P94y8BSPLx8mrJHC2QHLyXuUmHqd7hfGez54gxNrHcLM14xGRqZrNoDPsKsaKuGq
gCp+58/2sYE46YY7qsWPsbPbTb6u79Fgz90S+UjFyDCukDLwrG9zU2czkwKXyFAf
FE8NJdRUVIUjFHYsmTvX0v0GOPZAbP1mJK2kovRJvl2ri8Pt8g95Z3GiCxFB/OHw
+3RMAwU6QSaS37vdQIZwH3lvlR4xe4a1qhNexh3X1DNI1hE6b0E7fwwwfpDqY0UK
OzDlwTIdNqC7jYZ5Ejfnne4HUVXfyFWI8Nd0194Q8TkpNO8XVyBDNmMDqlNHoJwL
wb2zJHI/jGwLV1JbnCUknL85003h6RuBdPSSxz/F3/Zl1070iv+sQYbI+Kuui1XW
eL/S/RdmzBFZPOXgKTJAH5TH0zSV0kX3jC3fFZWboaRHTYH6xfAKKY/MupTpR1Ls
/pCvMFlDUk2ULesnhZz/jO83qAv64QyP5Y035fdvHHyGIpfnZf4GRL+k0fmjpLLp
9Y9/VY0CPn1vEZI8Y50x8xyuoUtGn6dbKZLwTjsME6x+ozQEhBR0hx1+XH4y5a70
S/LnYBR4H167hutx+fLww4tsYofUbNjS13uCMWLLkZd5rpHodQSxoCQPzhqZOyke
4mPPLFLNdosK4qA8mafGG1shGfRPEBKfi+8Q63BZkz4Den148Ca0V9VYMoygHbE5
Rusq3Be7id+qOB0oCxHexw36rF+wN4iCGtSoJGJSROYJ7VPULahaoq4215IfJMrf
VeA3YALAX+WI+mFTGZONWsKcim2xJ8n/NduboxxxWxLENhKls31YTvDfbzNzNeo4
nzp1myd8sCnmHRTq/Uk4nwLck7hgs2zXwy3NSdVDrqZQEMWKtbYPciElWHoG02lU
/EjMxoRWjWRqwK/fSt6GGYMECNIbECihaWQ4ySNpre5Y4OsGlr35SkmcuMkRKSkN
fMWLRLK8LYnhT6lGP9kXMUto0EiYCgAXTPtKNRCdrf3o1I43DB9S0VE4zwFyGHnD
2DD8yMDu5KV8mU8eaekWvg1PTOlT/xQrlqYUyRnerruFEuo2cFlWGt2sfLK9qW1z
s9JIpkuwabAljdWz2tWN+aAeh3Y8BPdILRvN2GQUHn8Y3WLpU+rbYK8dZ3mwowvw
zHG6I6GWNI7QXbcDr6Feq7u3HMVrS4c9FFC7fYgUHB8z/W3Xnl5N8NUYJ6bsZjUo
N2jNkCvhCmBzuZ3EA3L6va5ZSUSUZ7Ekj6gs9QzmL8vHtVrYZhwjiM/N1e9elugo
lrR2Ip2gMJLYOau2SUQkDumJLPuTg+5S8SuKUNZ5M5vUnaAJD9iLIl3AHoMX9ip2
ewxZC4GeFrc7CigGo/3iK5O4wFsDLzmqgKLzv+kb5hspRyOMHr+ePtoI9i/rO7DM
/NKBgMcMbOXEh0gwUaCrNncHo4tPHar9vkrgaY+1L3l5hmRzsX18LERZFynTiCJV
DUwtfAfox7Mzs09w1TaZzZ47rrSqArDJncFa9pXHTH/l10vpwrZWMDssnkBifNZH
/JX7gFHBRE1TChxnbW05DO7U7XB2vXZmOx4w2soNSq/TTkBKLMfPKiF4aXimt+Rv
6wUIiexO0ZOepmfq76EJfNem61yLiC0I3Rmd9V8cTqkXtebc1/5bYJ1gUH7XST43
sWh0cUyNGHCeXc7+rt0KpgBbauMhKT9kR4G3c1E9mGGHAW9uCJoaa1+e3GuGN6H2
6XNjWOwkySCVA+GxG02dhtdJ0h/jB+1Ed7J6NEaN91f1BB0Zlg1p18XPAsYMH/JL
NtW6NskjdF/ailAfeOCRxLIYN/juvvviqR4oVNfZdO9iX+P49Xl707nDM5YHYl9J
WOfFbIZRmBEYR3b+PsSexCOmNfC5yH2DabBPa/jbGHvCxbf/4zXpS3XiKKaBYQKG
XmoFj84k4SdhDDHlMLEzA1hxOQDXxndCUQQoJbD4Fih9aGfVXgatfje9hE7GemRY
IhNcZjqh9Ur1GHcM58yDH/dITy3A4zaaqnMRv7gBnjXeWsu6XC1F0DOhJN8Qg4+s
x404Dl2KgbjiChvdWTJY8lizJKi0K6HmxB0XsGtBcLfYOjppBqMRYBSNtR8uA0kU
iUd68pHFV8Gf2oK1DwXotjpItUvREqhkbu/fxJC49fCJIsf53bcINPkFBhcIAjbL
BQRzlVT7TU2ZqRFNX/+/mjrmJvUgkwTV20NkJ3Me+2WIUQq3FcojhTBL8RHogAoN
awFEl8VpOk0yYQGmbSfTFk4BMN21iqgGlDjO4kWBiyLcm/v53QVKsT56zNUPDhzH
XgashFj7fQvwBbUaV4oRrHMyCk1SVlTjRQF2BCt4BjBqNKPtiIoTCeFei9Q9JvS0
95vUlpxs6kdPZToa5Sjyk10rAm/FXWw1bzlMPNc1K2FWfxweY3gLqKK8NdqN/r4i
jseOqHXfOpf1VuUsud0ptk8vC6yHXP3/XeG0XV9ykdhPEJtyGtTbj7fIXV8Idrhi
6sx/L8gsUHZF7viI5S/QG8ronqnYr06kiy/mHw/SnHc9vPEFYp3HHwa2uXLMjTKq
zknp8eUIDUGxQmVWlbdC4WVfLA0WgOcqUHmb77753yTkZJLkEHgs23fSnTCcIQ7x
drIkz/sY4q4mWgBLOZil1O4mQ4dhnOmq28LxVx0LrSiOyo4+rsvfbiv7j0U1C3Z3
Vnmsaz0Or0W7TEawYN63QD0jH8eJQ2kGeYesiK6iHLWlhvCD3BtbwUEDWAKBcsv5
I+3sCQYO5ltFFF5uPdZb5tAM3jrHYPJ54j8JcM/DLgcwd5och3gADG6eepM50Rr3
WVG4dYH+2M2VwDQrIGHCoJ3ve1IxVKbxgZn2Jr92iNvS1hklJd1NWLSufgy7ai0B
rkJdB08DjE97yv+8q77hyJRhIYOGAyT8yHBKbSB7xDQahwnINBUlDKaSCxmOf82C
c1Y3nMTfsbuPYPJ6hqHbuSqjjX+LeRl4VPk/z0ZI1UMf6xMhIwHNJI/naS0zsivE
ULoG2TIMQh0vRJRLIk7ZRL58jZbKJexSMfTqLoV5RrtBB13u8rEZ0kQvb3SkWJ29
OzzF1/RqdfG4I+eVq/BvTO6tHhogZS4fLt7FkDBBg5hkEfHbBnqAsEeGthq6ih0C
vXanH0O0PbedJz9SFmGaNtHFrsbBcR9ruyvQOrrXN6b3i1n8b3iFTmrRGkWkn3nh
VeW3rY+APgwtu0IWPlbs1FgXGXyzYYWLuusROPLBdslidzHGM93w9/iwKP7G3EOn
mFXgChQ2tD3sxnREP77J4zxa9mvylie33zOyS9c7vFbPoN/btnG2Lb2LYNBp6iIE
PR64V13UDyjTcTGJ8XrMZLAbqz6X8KiMHLA9T4iOd/anKRWZNiwXmS1ZURzKjFGq
X8UgE0VW4avpiaxGWubxWDYAj+y3VhyZMGE0O9wboSaEyi+ssyRIAXa1d2YSA+4J
a8wOsq0SAtV4M0Oby0g7qHoRBN1u1VEia5pC9AvIdozIEZIlSsMlkpx4dkqKg1t9
FePahKrvCd8h8JnCLnv88DNMOXV2d48U+/1fwtCTWR7BTrICfH9pBHZR+1MJMlfh
jgEhvNkbD3mze8Nr1VQ6gyhlKudhQnOB8uZ5sGmItlzTPSWKshhNv+1hyl+PaqWi
PPZsKYiIk/TIYKjgKVGuSVqZ0t5Ip82+wztlvSv8jVUhYqlNUuZCOcBPyIrgJnmJ
McDKnLZQrSTYRnjJJjthrdseKS1pIhTtFE88Komu70cDR/K42Afkb78WqIv2lLoO
SDHZf6l57WdjzfiHo8ltRMRI16tg7bXQjplRepopu914XR9bWBQgtAByBT44Fvue
EM7uKFrWj2J/Zc1U+trOoIzk4nylHFTwOHQoBLTSAR7jfaX5gXbSXL67hmzALqRi
JBEIb4sZCZ1dPHvwhyhan3y9xJBe9iTAGUDu3KS3IPR9uDlCYqVkaWbqhtN5YCI/
Ix59ZzE1LL11UUYnISUNe+DkmD2b3fw4Id5cXwNsbZcwIzfrs6KzGjNk6BTq0EmR
Ta5IkRT96iYvAI93+KTrS+p+8Unc+j1UynyMqDNvT4umPCM8z3mP6ezhajVCOFb6
YrouHGFXO4GFppSF9oRqjEz24eJy4xeyzXpHfiH89EraME0LqhitRwvdfF6/qoxP
CnOy6YCA/ksXzRVrjVc7frUsgGv0LnEL3D5OVYrVEtos/0OatWYB3QA3HsKFkgSY
1qySbhPtQ2MeWWkBPZGkVkTEQfF5s4vr3JhU7nrabeXEZfeMZ+dNkeGJg9duGktf
uoLgVKE73gaElnzoHdYgPN0nZy1cgOTn4sb/YMUd8cVHikQGLwHhVor7KgAFxEj4
PhwmU1zbt6yjBHrTidBb80FDKyMh9oeOy8WfuprHNRw0NPI86hU2lXC3/vDBtPTR
P/iylX6WoE33WNlAwZYZ2lQT2cb9zGGPCIoMUFhS6dTOA80AqloUN/rOwAdXo6oj
ZfoYZxyV5l7KVlCKpydnXGn98vGbzVILqnxOalw/QqSt1KWe6/JSXHHdEkuXwQbH
A6qqHCH5c2sn6KMKAvzjbxaciteSIj5xhUGxEg8Af0sST4Kw5B5O9luYh29oFCUh
cVG/PJugIF3CnSdu0NIQptWIkER8le3xeie4Q0+uRbSVAcWfF2witjiL7KNCgkId
hLkixX4Ya45Ybm7A0zQ5hR48v6HqdohCkR9KYBGidXpc8Ef2OBYDGI0989ouryJ2
TzgesbelNJBHJDM1M64JdYTJD5d2XW+giQ/OtJklavdytZvoxJLdstJjRm4mSXds
dRHT/X0KQHj8WnTKJPm7xlTA47R/l3sQRHbbdQKIXn08ISwfMSLJfODDc228gThe
3N4BKbT8tHYGq7th9WnEo6eZRKSftDKczNwDI1aiml+oKz2W89Pqky8fo9w7KrOY
jwrtv58xEKCX2Fl/I7MYeSo97uUdIr28V2XtidjA60wfsIeyjB4XrcBtjYSvvehF
FeSNWjPwVjENc/vfsYRFy5yL05W7rnNIcpp+ttbAvnS5NK9p5JoGYwPkQGLYloLs
YBl30tly5hz1DnVa4MmnoQBlVzVUvGGlVwgqdm2QbeqoYMHjaWd1GQRqzpeXvuWW
gi824qcnK61H+XXO7JcXOQiKJx4QD2yD/gCwVokCJH7Kf57HiQZ5ztav4akUXpP/
UYpMoV+MN7YvxOrlj7Zh7kWbhDetLwSpbEwK3W7pGjRQIwFeyqnrAmkGmyW1pgll
FH5tkj3J6bSAXlegEMKHOW1nwBAj5lPCDvO3g+OIN70/XK8xOFC1DU2OtDAuaMJr
cMPMHW1Pmmp3ktrokWZPe0Taynh4QKAVWhhRyUL7jCXxWCKaHfko7/A+rP+ifJMj
tFdKDmb3iPFGXMP648C4/MA35K3Y36CYKvGkbg22fotPCoXrF3lBrPSGAxG6pz2u
9hqa9uztkPe7ekd+N8BxLWULtM0e9pYOJm1u8X6v3DSe5OU7R8MuKOsXKFUrrjLp
69FikwFUdPEXzHA+4jFmTutflyMzU6y6sz88VSfCwGg/y41cE/OGXvXynmf/8Edh
cruiJlXnOlLj1Hu4jnEMZVbhIgJJB3zMuIaO1A0rrMD5nHomDJtcBdAk4tUVyrG/
TzuNf10gUHBoq5RlQCzaiMSMDYIMaWCvk79e8ZFWx4x5Q7+E+k3doWgqYBhxqgpn
LkcR2qghN0Jqvy+yN7MlMnV1OuiTH5YKB69JN2LqpblfJ6W9J2qIld0V7kc1hJwP
CDY/Vtzm+jOkL9aT7Jx+pHUXLzDPLmDv8wkjzSjFLEzXN6uHQWPQaC/N3gWeQ/k8
zBBFZ1qvO6xj6rP6e+MFO9vJrmvwKVnr4Sl/2xAAYHmnCQDyLQDZGjck1G4urJ7s
BBhZI0YcwNa7U0bT9gW4bvcu2MoghYCXCI13BqdV/0hGOxSJWqWicKKta5qiZVIM
JDlG+15Pvt6V2b/3QD3wO1GAno6fSkX8AGQ0Bj9MmK0HwHBKUH9yopnSEYvpYfIl
CUMEsD4B9EuH100dpHpOFgThWMBveIIpSGT3I8i3ioThbqS4CpR3R7Yp7n/j15Zi
De8fLePvncbhHbNS35GwJscsltlTGIr+8tf6hVU8QOSaGZZrPsDJyX6zA18YcgjU
1LwLiO4NzSWEREaM430XEz5rMqxXuGdd4FTUm48N2bXZz8/d/xuwfHyR3pe4CxZu
ffP1b/lkzWOesj0/qRZOm7dLz8dv34JxaFm76hHa198VDfml1vCdWrhbJULJwgk3
4wYn+g4d78GQQr0yrFFGfNxr+0mOfFRsi8Jwe7hqu8PQ2mQJY/exn62IXOT1gD0Y
31M8fe6CfiEVNllo5j/eoWGyp5tCtMSYg5Gzgzf3ItPqVW4pZNmy5hoGSRj1kxCL
TY6Q+G4np//sNnenCJ//QaEkiAEDsLuN8kewNJMKc3JouF/ikvF1jvYEP8JydD6O
VuyAn6/9SPR0NF49M2B34Wi7iaZaqfGVjb27SNS3N8dxu/YR+x27Fr7V2GVPtw5f
0TMXnJRFZ/Lat5UIXmq65S9T7sUbNPr1LMVYfAo3uIqU91CuWEFPnp1nwpyUI3Sl
6GpKdywy3ZKo8Cx0Pu9s69o5wPQeEciBL9o/h2acfd9L8lCd5bYeoBFHgXN185V+
Ql0gz12KClRW7+hfc5IHyGMeD1DDQa6UdJIXwDUbGvfNU4bHeLyXIxEyqlSOzGuB
yrYdnulErvxeGoKo1BPcUQw7F/B6cFKw4Bi0Sqm6JkusWf+6YBccdelahaSAVxv6
bJnQiSpWouQ+42rWJzDi+y8TYs/icdBLpJ2jldTFbhvFSYlTGInjTWv2wsSiHSsX
W7Oj59Md5UaVDC8RrHWfRWUlPaHZDFAQJMJ+3IaYYczvPScpeRTQDOuA2ooOKh9y
k1qruuM37o3yrmiq1dSvGqX7QqM9Ict+hhifYj1ZfSUJK+1z+GDUqGXWnxL5u077
Mk2kOarypS7SM8ImpEZcdfKeuyal6FDrNpHtH+3kZlhx92QiK5msFoPAhw9tZn8r
/psGRXMER+sk6geAG9hjEJK4bTNtfVwAhlVmVFezGOIDbvp/Mt1VNsjT8/KF2DzD
5mYCCdskzZUUhmxUPPOKd8WaUrin3NwSYtK82zQKaAKnqnwppBB4UciswsEnzFsS
1fCzfXENjqwKSwUcd86Ok/msp1SSZlAyKeUxy3anwYlfrIt4cai0vFKE6EV44yKZ
vKiDnOHM6+40tmz6okMDxJv69PJuprdaujyv/5tWIduB4di0S60531N9zqg4/C/p
f6ll+SvsT0r0huBu5C7jB+xb7aCkW7NPAoeiTxGnOLVm/suDP9wqFSCWwnrB9zkD
xlMZi4cE6z+T+zeUV11Qug9FaRKJ7Ll7m5rXNnyDReD4c9fylZQtPkeJoOi1A3LW
JMoYb+mWngffTwAIMznossuBjiONOZcOYl4JvTejEQLAzGRUYKUE9Loa3Qpk52+a
ov9m0ysDmB2odWDsez7xRwfRrdRkGusz6ztcpYI2QOgyAJDg73Cw99PWU8XO760e
1v2gWWHARoevV246Xk2Qjmp1jLYYAMBcBgwId2iFfIMqGQ01UoHJnAIQVQ59rseO
jG56NDvb9dlm+vtfppWLq6JwDwYGg5LuHQgJ/tfS2Rn/+h5MUjT88N4xVRlLIhSw
FBUZI1BDfSC0JtCSWRGsPXVURdOL76xxMnyiOyKWMOXXY3MRJFVoH63j9PamBJX1
n/uOVx+wfK49jzJIaU4tdflKbtrCdvssInHk78krhl9uUb6vAF8XHUAmYB/P3IUX
yixpB4apsx8J2q++0xN1GiBFjha2JLdzdw7Q2DlwnQqgA7pIarw8i7QKTGRWYo7p
TvMCCnoNexO55dvIxWz2N02zS+yaBM8cKf/obtrP0ssnOB/cF83C32HxQrgNRqNa
KM/qtpp58QOyfBtntjAlDnjqjZDioJe9SLM1Wo7g/dUUVUQkkRxf6jVbihTJj1IZ
plZbvRLyJy93/zPhnkZZUvVh2TmP7NrHxkvioptxO9zR/Vxs8w2XouWiowpXQWDQ
Ve6izhM0ELEnSlDSvfnl1GHUnPXczoTgP0eaRkoRnRveL0Ed/h9aYe+y3ssftUpr
8lJ5fHcFc69CmkmcA8XAxWib8j4e43mXnZn/LFq4Rte3b5WICD2tSEJcfPkN2oeF
UfJabvZpdLNIAU5EmEAN59ImomKOG7oiHPr+B2KK4cONTKnlF5IxsIc5pukLDAWI
Um2jH8ym7rmlsej2mdgUSi8NGK+Hfby1atrvggOpGE5lnlwCIU29qfIGoK1xvZSt
cwc461X+l0VG1zkI5CmvtfsYsJsey8o0Jbv+LpaCgTU4T+RalA6p00hOHwb2b7Ty
E68a92wab3B1GIliLi1Dy4ksnq0B61LwP2i6ADxBGbBEOdF5UeXQSUcM6uSJhm7d
a/RveT6He7gHecznZiJVhWtJ2hMtDLqvb3hzwpvmx3CnSXVOoTq4bfpQ1s2CsXT3
RA+DruFAEOHJalCy3c6zZ2KjKzgHLfzV/0/SydZ0FDNk04FwdHlsW3z/FXDaRlqK
zHCGUnQD6vRfE2Ppro5l4WOdOeH30NQGexHvrObb+gdfoJsBlW22ssc28fYMxcEl
a8HIcFBkeHKjzYaudinXtdvhHeMBjAojOSQx9wYjCY/3krf+7a5wB1FigtZI5v+d
55ElVoNShJZeP0QteE4pwmUwtVu9lnb7OTXPWeqm/VwfSE3F2k4pLcOoBVzJoKR7
okJiaQ/HoKdsKw0lFFy6A+MfJxibuMcgK9hH/ntAshSDw6CcCxmF2ZSvr1pLu+XI
8Dmqe5t9Ykm7idKkSApDbi7Bxe+kDycSnciMTcjssekttfZpxrQ1vZQM0Xg0cKWs
L+2P1MovRf+1y2LZlzW6LI7+cpJDMgrytfmlrRNy+2kXtZiYy5WLnxadIOk2XgMW
hKt8p8oDdMMR1f0J7qs6G/lbgHh8+4nfxNdbOcAVsv9yl2lsLb3YUmFnvI5K9T7Z
jtOHolkNIuuwXVLq1CVs+YohnfJ4VKtE69sm2fxoiE+jsA4bjqCxwEpEolHRVIJl
ixsDd1OIWLrAlnZXSIMh2XCR1OCLpjjNVu3nHwFgzwzzQGMg3CI/2rMeqjTMvGCH
Tfoy6Sk721INNyhYodQIz/jC45VRoHXX5LWyyR6aoETp9g6fuPADoEU8Q0G5u5JD
/L6BrBkk31QC5JHofvP8ytI3FlEmwK8YjMTIRpC0SguNcamXMfg6o3k20crU7GD9
CULGme/8vYYqcjxMDpV6lwnpcpUQAxt9sTaxZMXA6QLasjntaYBxQKLRogmwwVsw
DwsDZK/il5V8ES0EBi3OCxhZp0mfS2vdKtRkA1iplnaI5LDd6GQwv5mu9ncHinXF
cA0FjyRQiIFcnQxkhZHAdI7BHUQY4DGPJbktSbk0Ej3xiIp6mwsyySnJ0I0Ylhzx
sIaFW+OZ02gTrpfJQeii9rIaFp8z+NGT7JOFHZQYG8cZ7O/nHmfO4SlvK34XK3zY
A3RoLfET6ScTfwTopD5V//mqpya1uwKVslBWuex/Uykgq2pSLFzCPrhw43HXULzi
xtdvx9q5HbJzNzSPiRWSM/ueeexIm419w4DWUoa5vsJuH7y0PGKStE1M5RNYdR1n
jp06Z5wzfQzsNLC7r26QhVvw2h0QybQWszyePstbuAiD3RzaLozFwDQMs9LjMWEK
BcerOQnBJNrz7DpaN7QucXfK8FyPvt0U6oZTflJ/d2kiyNHjunSwx+v+51dokkoJ
3lQyHr/UYipXlI6pC1UepHeb0stTsq+VJq6ujEvClhyLkrhEhmbtkpYY3/MkNE+F
jGIi0+nReJqTGjrsaJZqn4gdvlpayfKVxodHu3/4F0fIyBqWwkpUeiqrEEUp3Keb
MDkPojFncg5l5QSF9+LsGiI2PTZP68kNxSAP5V0q3cQAi2AR+OF/qVZpQQmtf8af
6wS8YCR2/drxZIngiOqt4G+0mmiZ4fsXOgOcOHoy9XEpqh8XGumvL+IerqT+42GQ
ygEytPX2HHxnxhUSjcUF31klsu6iNojLaLyn0kiVQamPGDugQtCpmHXGQ6xclGsg
Wztfh0/I+g4ZPfBCHZ02mZizsc2Ni42bB08h8Anz0RConM6y0m/lM7luHCaqlg+s
jflFb8iknF4qwG/deXuVMbq5KmOQnR7MNtLJFA3vGl3TJCO0dc1QMOy6XuxE7F5R
929FuywL8JLYkDFtDxh0BKOg3sOkGiPU5G+OECva4gBOsKAg1+vL5jzCpl3IK2GJ
4+EAUVoe4ojG3jLEO9EA30tSLtjZbPnjC2cveXLwjiRlWpE6GVsaM08bUuSu+CAB
CKjaz6PMCH1+kW0952N7wuEOWwy4q9C0Vuh+ka6OfNc1cuCifYYbBcqPQ8I5fzbk
Cha7aWS3YsYd1R2tSwZky1pvgH4hldLf2tsSaZxNDonxIeHLepf/jlCcZj7SxwHN
mzWhJdY2JOim9Quj7KgOdRMR628xPNrHfTQqv5U6vfM5wKAlTXm2Iv32ASeSXz6a
n9QtvYwmpVHQOqe3r1VxD8BBj1JPClNHZoxIxaDxKDFkPhMEnyZX4vQ8h1aphgg5
TjtkD/9vRvTXKITcZImhKEx7o3LM4fTc9deSslL/XuZR4aN/Qsq9ZhmGYXlqwb5J
PVhJXaY7QkgYdEPKIsRPJMQO8upt8CBF0ojHB7+GicsIsz2+r8+OCnj1vjU6vfht
vHOMt+vaCbYJiEoWqIodbjBXdYhb04SwE9mHjk5Q1A40c1GyMxJqHH1cWiL2u1V1
wkvpr+eIZ9J0GTQd2APzCT4ATw6oRb01nBVPJ4uNAxErpcObIUgG7duVixQZympI
EuE6Rr4ngLOY2n4FNXG/n1SMLYKmFGM0IRYkremSHif53og4jf1sF00N8HZKujN2
3ihHDWV7zygad+G+qdO+j2INI5Il5JU4AfTieGS6hj+p1ivfvsGr1f6JWbctdG/x
pNOzljVtJB8H9vwLxoTcV4ExspbsrWUjoKCuYqBHcMYQVwyxzVob0NHMWOzlx6Ap
edz+tJ6wAeF/22t6QnJsF1h+RoFKup5tiqJcqI+xOZvUR3I0I9yh7gTGLJ+PQqea
AyXoJNMamSgQM6pNL58Z5VhV5ZeAoKpcnYYAICiMX7dazsnrDWMtPllInz9d3cFE
OpAjfVGGnsAeHuNUVxmADyKzEHBHPPgOosE0Sygz/7uvAaBOs2BQv7Q6zDwQWCJ1
qPcrvcBL6acDPf3LUm3Y+sD+QBHIIUTToW+Ww/Jemp5xJZPv88SyBZaRhtgkd8Lb
YKChCrl2n7GuKiDkm+Pft5d1fupp81wiPBd6NqqqBibEepQRiLB7NerQMPTB/OsK
yY0otutKUPIHi+vq4FQZSseFG9ZFshWerYN806D6SVMuFifg66cCLqM1B0Vpy/Ci
SDvlK70pYZcyPMeS03hPGRaHqd3qHbdnd+LaJf6RQlmAWnsD1rE3+neyT7yTeozj
4uTscQXlb+tqj52cLNRBHI+VNynuVl/fr+c/L+iInfycey4q5Glhz6nLXZL28Sz1
PDgE0rhmNAMnWlIp3+95NSSjDzUEQUauPrlboln588Uk/UsDmwvJLMuw7S3OVfOw
fqDLfVoz5xuSJQuv/tHWFJtdc2Z6D0/thKlqG+JX6FXfdTGtzWDfAxUtG1Uz899J
B/1lVIfOojYWsz4dK1cLDgOnCa3p2Vtv939eXALq61vozPUbs9lJjyFMn26sbXZ0
stvSvRApqd2zBaVFuxmfIiWLadO4sr2gRtSqQcqmNr/dcIjeiJWpAgNC/Du9rOWy
VVBO3IE6a0nNy3w7BeSR6x6/R3gtB1Ve2xxQwibEK+awWBM0h8NMdElzo5tJbock
SBHcs5N7dmi71Oe2Y9ntES3CVeGYTWdCVlf+kpaZApQA/Y15BELC2K/wBHxYr7JZ
n8Od0b08/hm3KDp8bA2nYXw8xtW076RAfHzWOUh/2E0EXliKDgHnDpyXX2ONYSey
9mBfv3OY375UxuruqEXcr9MNWdnaKYc3ew8SvA4HbqaWybjZgbrS+p6jdUnsbU4I
R3QDtb4g4u5UJvmCFSv0b0zDKPjXq/ihjb3zTjP6T+hA3GpynLI06B/XlgE2aS5m
6iTDZfewLIQ3WgAmxbX9VbWh9KnbswA7I/8oJCCthCz3l5uhHUA15n3faGMVafW5
KQ0qCR/IeK+5y5Ihz3BnLp0LpjDEGNLuDazBFW9f2+rb/dsRUVyPbC+lTDAd6EKi
GW10l2ZrvPJ7bDDBtpah25EuHutJD7aH0qlzzhc7WxvL8ufPWR3xeNeWcI5n3zVV
+yB3Xmt/hjd8hQMD/f4i87zO841JinOXXC3AYwnz6C36WqeQAe+gx2iDha7uU781
2FktSmmRkxbkk5f3dkHN/1UDFVlg8MAnb6ackuYMlEQguzAG9I53D02rA4TtMEPh
9B3kDNLBo44zCz2NItBLafCGqwOG9fohuN03P7GubJFOeOtZJtDuCjVPRGqRbHaL
kU7wdiUsdiulWzitcu9wC9/s1ba3/uOfxU38ChsNcX6WzcSC0CDD8HCpK+28AXbk
4dY1M42mwESaTkorpU1ymIv5oL9nMRaIHLXpegb+79dL/Zwl4gs1VRXUaW7MVjlx
scNL6j1i56tW9GL8aRKyrWJQTf395idtbEZqCOei+9OAI1VxxKYFBne+GBfrFAac
qN8M8njow9KJn/qbAC9Wdns/Rl3IAVkZVo/zSE0vaJeypY7TarTU4MHeH/ABItdI
ihXDxSZWR1FyLbPZ7xLrTPPexnla/NgUJdiRe3l53OjkfzQgW+0DCivKkTRl77Uq
hWruuqcNojByJ7jnFLWR57tePJeKpSgCXq+p/8az0snAlIg3u4MPCoE5kXdRzHHe
bNLfzgKC2cAePLLrlVMsS4QrzytP3DAY0eDjX5FvZcKH1ElG94yvJgZU0BuiGuiU
3RtHxYvEwPoljZZR26vuOk/7TfPrZrTT81WSZW+pNnVSPqzWeNVVYEozfgQp3kGn
+iZgRhFhPK7uOJYUsoILBgxJ9bxwe8GlHDVNU/LJlikawDd0F91m7BPCey9jncpW
bIWNfvl2nbSQkbz1Q2K9RqL1EquQy21SRXaCo/o0GWKUvgwNLCxP0dEFHFsDxfYq
NsJpbICXfeBw8W+Zy7KZ+uGZvl2HGHT+RxM2e8uUthzjUzKCMF0RSCB7BMFd6iUM
vzmxf4ZJjWh3D673/tLnMgcGPCcOiCF6cYAbffkBaaFkBQQ0EkvWZ3cJPAioEYJ9
qTrhLkpC+doeJWCLYjDyXGyN+wXgCWEJssQj+Of016WA/fdXI6zt5ucwkoHdvf3N
1gkGwlZfnsSQMJ1leiTgJYL85gJYayxb3scIATGAfsUV8rvy2bDgzDrfcD0SYNZM
8qAmruoojEFt6I+d65PYPrc7v59jeesI57cXMq4yq2b43R9uE8fn2gTWYBVYNTl0
i7qbOVwpiaBqJJhGRZsDjR/M6KTKerfmvy8czIpwlQOvrsIi5ByH0c7nUt7rGYNV
Il2M2soHpKBIimf3ta9hq1XTH53eOmX6Hzl7Cvqsfa/5DE9eW8AJYcErpbuMmpO6
IiYBiX/iYMGa+KercVj/XcTOWf0smzHC4BMNd1oLJJz2aPznWnOdlGtOI6+jcmq/
kYh4hJxSxjaN9tYthwx6s2ibmdRDju18BhntiaTOtD7Edf0RF1dR7Pj23Cfsmr5k
QSjTWHeWJcSW6rrVK5nG7HKzceUtvAF6y+TdP76mKvlQAev4nDhbpcW6f75q609K
/KgHn/AzYwnFOWHUPxeHZnQ9+LNfjKnt7rSYD9x6QTpSKu7YUWSTom8tL87dGGJr
/tWNBvSs1nW23ahswK7DNafpr3q27FNVgLCouc4rHmMBcpIfzV4l8bI6dzG6BxVs
mqK5oJm5woZNNmFfJ51sp3UtUyZTa+HNAb/2rd1TFbr12URbfy6YE9KJKw5emtyR
5ZEyePQMdpxZmJGZtEA3rsYEWQIGkxxGM87vJDOt8r2yYizSSNBcqI9DSnm06tno
UOwfEs+ZNo9P6/zswLTEoRkI0RAZBowAC74/5lNsbfq0ZElEKhsbpcVL+ueDpaFX
9R+O4vBtI6qFG7j8IktFbFWk0kuXWI9wTMpXPR82/q9WUSVYg50tbxzVp8OAGxTA
2V4sdwN8OI7Vez7ThcWAuN9mNOaJd/kq7xQ9JqqK4XTaItJ9glC7Oik/2d+zBlzQ
Ag8kqeDXoS5u5QWXzOOB4V03TH+oA2j38E7gYWJCJkaJFEr1NJEJJwhegl69ereN
4ivk/kGDcR9CRGS4kHXYOVFjulaW4A2vSaAgfTn/9oxhIw89EMye3CctjQ3+NLXp
aHnaV7YLQZjstE2mv2j4PUnwsKkir6tPJ7rGJgOAmDDeB+B/uENyrPTzQ4gheAPi
Ve92PDbVHXXNIeuWHUBv2mmH5vHdOqU11m5CYtzAsOkB6uLN7C3LSvavYLUSOGQS
hhDYvWPWB9TLUCuNgTWFVPOBRpALi6c1OXSqZQcXyqXwSeyb3HnKR6AIGyJ2IZx1
A0fP6CN2pRa/NU9iqDRMxxs7CW7qsREK9zxSPyMU+BcPIe+1e+1c5QfjEsSh9o1Z
EUtS0UHCH61w1JRaf8wkkEdfaYyMbAyBEaBv+gS7/U1xKfjGKbZTezgMeb/AB3iL
SdF8x3bQJ+4JWwJirdfptbzJsl5O3a5baKEcXBVKmxR4V0FbjWy98WySVZV89mUZ
+UiVee9ivOg+w4gk9i/2JLg6/MJ3bHbtd2mClNN56ae/DkTHbLSHUXiS8xJe9RY7
o5vQ4iLqctjeY5AkgLI6b/Hd67KFOi3Jh5XRx4fLWh/ye/WrPEq3+uwqEjExqKeH
C/sRJanhTTwIJ0Pu6IFt8v9efUXEVYXZa4x6PUcEv8dDPsANChVV2IDk8N6Mpdpn
ociR6BwBJE7re98tPJA552h+3f1OSUFNUd7U8SIX5SgKB6Ng+K4R757wPLdNYljs
auDw9RKDboIvTjZdGGGbYbDxk+d+faEwjeNGk/N6CPWV4n7cNZ8OoZBGN2Ti/i89
AVtNfvSUGGX3MFpcAjvBVmyL1ldrVRImruSZNilZTsuCYf9kPqHuskgL+8DRs7SS
APM0eOqwvWjIH2R3J+kf1K/KsedRcIDmdLZkoZur2bSiEGjO0axuW00eqVpS3E1U
lSExBbyPNNHHYE8kQMzKcRUaSSDGiKP8Fror4ibTGiKPJkEUnhKMp/4x1cncWkRg
5z1WC5zK3GC7LHEmKKHFZurCkhBmS7xanhTLEAX+2dOAlJ+z0DoBb4NDQRcDeBgA
3eUU5gvSSRv5nznMmJEntBuKk2KVYOSiU7tkgMbZIMB3yyej6i8AoBHrycKZCrkx
lWCEbOVL4tO1Q/TqRahvW3biaZPvTBkGMmC3IHZu3sqZZzIthJXEMEGUU67kFpz3
6rUdT+OQ4KWmr74P2DhU3+Z8RQCwbLz48ivI9DRMemkYyDKIE/lP36PEyOynhp2A
6grWoKz6rQcwT+4FtedXqUssXdiiVgeu3lDuL9Qca5yMIt4XzrvDnfn8UqpseBit
8kycxGOB36aQ+fMVOalxSIBV+bi/kPjObno2ro0nBTUds9bKsTxT/sjG0dJ8v6mo
V7hRtys1QXjojPnJwUbRNyL9AC+1b6NDLzqor0NmXRVI7wL6W7N7FdbwpMNXKAg/
U5Q1fvx7CvUf4jT27CZMai3smAL3iecQ1k5MydC0zot4kkaMgah/dkk0ss37tEzP
JJEyUuu0l0A4jLre86GLMlYGEYY0IqHbpsqiB3etIvkQR+ZvauZDGFhXkDCIVEIW
rka2s/7R3HGM9ESwBqV1RwB8F1rH6ZhxzBXHr9P+bgJz9FyX9+3lWkpyMD6GLEVf
6qj/UmMERDJkS13IRw7d8K/1r7cRDEUEzpYhY0+o8pOpU635nhpzr0DxSh6IEu/o
QNSqdKJnx6UskQh37NRdHHPkCDnpkFyNg0OJlnv6N70UfNtsfvzH3Z5OIc94HWe5
WG0prEnn4Dd/fByIZP4fOO79WgtpuptJwPQpwAAR0FSJPgLPZLSu2PBF9wBJxic3
Yp7eparvkLdyB+WssIHFbNP5yWoxUF03psbArkbqmCCTPAtnw1LsWtS4aXFiTqhL
Qd9seVlKEfppV1Pck60BDJFmhVRJfVgFf2eHU5jt1Ec25weSuu3qJycFLHebHh5M
Iw/QYWmyqXlqImLK+i5FyUcEBDjhsXxywhAIm5k1R95hU9ZVo9xwqWuTL9lVIcAw
11tFAdnMHKHvEAvoxOr52whc+yqdxYnLVJP1eW9A1uRKDQzFWCjKuOzfZIlTDi4A
ZEd9uzfBSy7GKbgBHOlTiZ1G0woLW7R9Q/nD5dxPIDbLsZ6RWkHglb7v0SWeCslK
zF42ZPqJvkDpHypqZi7XweXXINwRV0ujLeBcPTZIydQ1y86+4GdXgqEtL0EHGY2o
AM0xE/QR8Vc6xSTREJGtsp4jZUqQihpXLuVuokqwt8EygdSyYAMhQJ+IrMSX+wYn
71mQ9Zy2UCpHth+zenQjFdFSVKImLoZkzTTdYPc4Gwl3zVjpYuB3AvEyoWnu6rKR
Yx9p9wz/wdzrOIQBU7RizUZErLIGLkcearQIL4+5201lqHXSc8jHkc8Iv9FTQlCl
p4VXiMrCNom6h5smmPEWMo5gIt9DO0Z3k07R1P7UELRIv75e4q2kuNQg4dVXonOl
H5JnDYssWjlNQdqFyTtNELd0/HGLJI07PQ3hcU8G4kcpcO7MWoRFR/cLkKM5e0ve
MTVDTSDZXL+0EaWoifpX24XI9u/aEpVmX8Fsyv2EMYiWUfDsFhRu4rKqaDtsqJbN
cwbnj8T8yDB6HAp7neBRn9h2vaVDmd+v4xxoywLNzru+jfiG34+CsL3Q3TckS2Rw
52Xzpbh/EhFgsL/uQYgfWt6UuSzRusFX86EmDAifEFfnJSYUc5+apseoC1+L9aZ0
Dsh9EU7FsE61QReqZETTpYJ749xIY83YCHKXIEgGC7OpYOzfuBVkcHEJ/On3F7ZD
C6l0batGAZvb8MMgEvBbYV3Lbs6HKtlDPIBjrOS9zwE9kUsf5vQNjRchJkdgfG7R
HsF7acwq4OdcOZPhv3Hz2Q4WHmlk51acJff3f/VFwnHLqGc1Us6fRRN8dzLAMXDI
C5BQxunOLSfgBKNvFFwAumWx4J/DOGLxNxieMeBGqswyXMaM+jKBxDzScqQeiPiG
Yq5G4Gal3F8hHXt1iTbILtmlc4eylREGeA6+AMLXBJvngwAXEqNJAxnVnkuStvFH
OjPv3lW7IQSxP4TGz4T0NTG3bD+HVhxmaOc4+w+gkmwp7lWCqCNfLsW5YQfugSc3
kXsvuHK+FyUhrh+hw4HJWUC360DaDniXYoWi4omKq38wxDwDr97JvcLaooqMSmyh
JpvmFA9nkT/saJSM8+IaYTFt3Q9Wv1z+IdhC3OsC1jX8QxIszTrNe4moluflli5t
ZshRwJ8fiEc25tp/ukJ+eKzFBh5S0KtdnqM1Up/CkVaXoKfix6s4al3fBi5crQGC
Rgsi98Xd0RAMTn8PLcE+yhFOu1XQKMJxq87ucv9R5CovDsMY4E27dfFZ7SyLFrfs
vU9QSh+cp/2KFNY4hbv9ukpR6rraQuKrmMG39PqyWbRuzGIDg55PWGdkW6IWMBwr
TIKPUz5cN9Rq1rRv2w85vo0BrZgom//dhAe+/EyFG0m4lydFw2aQ9jyDH/LmDeoH
+N7A5yn4+yAQ/Qf0IKTKo+zfFn4aslvzsrvH7pQOOucLa8ms9MpDig5rfnhfjQLx
6pOvp9ruTe/Qru73up9soStxPtUQdbskQYxMeLG20fPZmwDHvSUbOuqlVBEe55j0
HA0YGqht10y0UPWRRq0PlrvFv0/L18H5+kwzbQTz6g87kFEA68IRvP/qrszQiyvF
Z2ommsrh2zB9IiMbaxXbCR44eleUIPV+z6G+5FA69cxKKFgjqzF1IwL9HDJp4vCA
/IYtjWfJUVU58Qe5Li7KLEbulEdMqSyD4EfEe1wocAz45rXg0FKB+7JwBp3afOk0
72hB7IbUN1mtw3afZwQC9ZhYMX/DApMOVptEtY/MlK/KyCRvXvI5ojg9+KYm6hf9
2scr5hH4tvyc2ytwim2av/WrfboTyME3dnLBcggGh7j6RnzflgrRtHMR52lt60xQ
RSnfkopIP4HYE53EDg56YTOsyMhden6Iik065Sv68zT1WKK3KR8P9YufGoYypeHH
SE9S9mExJdMw0KBO2Q4emt9qJG1zFHg7oMxzmDGejTfeyjkeZPxNjK0IZRJj8bv0
NfpOQ4oPVCG4iZFEq+18lQLa5ADrmOPL5xU+9vLLww94WUb5Ck+JNA5eyKTfP4QV
SVSNEQhvITdLTIoMn9PrAKtT+lMw86Ite46LEpeggn0cwE7gi7F3VIFRXTd/fMBg
FPMFGjn7NuOJ0GxovYU40ImbzqTQHgfQInsoGhbnb09C014FulUVieG0bXUX9vWg
U1VKBrV0ToEIoNvueha2Dwnon+ZkHcOTqgqQngHtAyfXJozpzt3mlrSzm5ivviKq
/Ku60DLGVhYoXC/QSgO4Z6sXCVa9Phxu5Lp3fhCzM3gR13llJkAx8aYxlaqVET65
TCzk+raV7JYeJhQIhpP97P54nomwgwE21p3sqpD8y/j8OwI7ilmnnJQgDsH8E4rJ
xVFZbTIsIjOK6rxRnPbisGDbjhSJ7DpRAfhN/K4HiS6F5Zuer0KtnF7uV2eSFoe9
JGbb9IVkEL2Xzat12tca2qZJ5tjm+YTs900P4F023AKMJB+SDRAp5fRGNZjxIgNH
U0U/WL7M7JmINkoo2td/vS5xh52TPVBXiGfVwv9+m4ECc3zp8SPdIpjbIs8ElPg/
MGoK6a1cRNX18Z4ZcHy+VVCIqcHaUjXuidz6rYm0iBit7lzNWlSOJ3cunLuZTX6j
PFKFIQMl2OtP4utYZhM3SqINUT/1LOqXNLgTpBk8hmyIAMnHTaxgfryQZ/Kr4D/b
Oc8MiJuNvfRGmiEnkxyz15LzWkrnY0yXv4BuOOSc9JCEPo0AxdtWI/HbRU9JkGe+
Z5xRDyjgBpkMzOHvQN0Nh+fA/6Pk3j8EjY0ECSkwzZfah61+a6pnTUCsnc8riwx/
Cgw/65WaU0rOEhBvJNq1+LRdCJjUUB9dSYtCQ32nsEXxuwk5IFbv+wNeLxa2d5MB
I3lIO6XaMJzXoSC0Qje581N2bmvOA2RY/s+HUTY1xL8+1G/pqWfSc6g8gTZplroE
PPeb6L1AFcFTQiJOfR9fN7n8s6byl7zkbxL8gkQjWdIGK+RNO/NP65pKg8zPu9ZA
icfp8bXzogCrt5D2WevJm14LTq/ASZOW3+i3s+l2cSADlDKUciKr3JNURmMulvFs
Frn6/i6jpkg3GBsaR9Kdh8XDihcY6YTUa/bRIuOJu3u6ToJ4l83S0cMot6dhnuR6
gEruqoJJHtjIl7UsDByGMEz9orTQHMlI87OhBo4zJIaQKVPz3B7hvUVmcPFn+YSX
12iKFv3BGd7QfVPMEHuAsEZM0jjVnJJzB7buiS/9Z9621EAKipAm0uPmwk9EkriY
UKlPRqvQB4P6ZhsjPlQqeaFD6mG9f4jq3kH5GX/KkMau5UlNaRrVSIRMHtQC6dUc
rPDNzQCHTj87+63+EkdGUWMj7slZwsKfE1R527r/GYhpUVSYSoZagBnRDhS0ECtG
qpXqvLM6ipXnAFX6X8H8Mpie3aADxf5Yy4iFBSLdRoZOrUpxejb18anGM8M6UQbN
0jqGq1Bn1WdKlBx67lsYNXebf6YjxyUAHLYv2wvxe8+vlfcgOgBUv9fLppZcOnyj
CduyI2ox5Tq/3Uiag/AX/aCGbZGYOSqvwYSzu6wbhg2TOUFM8nkewmImet4m/m6/
+cjVlzNMDcE5Gm6qr8m23qcKhaY33+OdNgZ6dPJe7OymXbM3G+X1toGMCnqR7ZIW
TLRqvSDeTeOSjegHxz7Yc3Hxkc6X1Lrba3enIEHVhDk2GTGqpoQ//otSw8PJMvJh
Mc5y/jKXCCwUFP1mTtDJd2w9/Wtv/kr8hP+dMfprNgGLG9uIK8oq12hrmuMDvGB1
3kjZJON3puej9ESL+B0SryK6wcZ7BwyQ2z3R1zKlybgjc7G6PXhU8y5KY+ENxoCA
ObcV5NxPf1f7HWNwemYrirhhTXYTwJ+l9JJVxN2h/LRr26wEGDgCh1W67aRFGpFD
EXZVIYAwal21DxDDo6I1K5HTpbKqgeF8IAjKvYmjUbZJAHHfd7R2vQRO45c47zbQ
QsDpmOPy3nKul1dNJUR5VbiJQc1BeAWprP6BFjRP6XVrZ/tW/Zh8LP39mmaJJI8t
4qba+f/eErTP1c1CmymjHlnmhoYWlk4k/wWPwFed6psAouJQG//HIHLhFl33Jgsy
ZHAdfAgjQICB3vtd5b0nlV0nh34dGcY2AQHJB9Dqoy1DB8l7+i0a7rBtB8XYqHkh
iI+uf+fgta5VXXzPhsIpAoycOt9sFAqxeWH5sJJA6+9zo8fYD/fw1BKxjgfXKLLo
yUPPpqSiDvoxkW6FdwC6+TmXenTAwx5gg4ek3ljuyrZk+nKPXxTsO2aDtoj9FVwW
q5HDzAndhBelTkhQA0cjssbodLmDBz7dhRI5VRxqYhMPwXEbbdhIQNy17pFSl5gd
CJm+VKSMUD2P7cg18PC+In35UsAZG4fwbMLxuD9hpPs9Ym/O68JJ4nHQDgyFX4Fn
JnHe375IIexLxFtp3r7BC+eon34WExqiIk5VwXZ4tf6u6VKKBCun+2tIMfE4oLrw
Lu1C0EzclTYUmFleZ07aL/wHsr5PU2EeJtoayKtNC/y4OpUIlYSGGjlnCHfAAXxR
HZTjh99edQmWxQq7UIOYE171utmhNNxS+IbmLXUyKam5d38UyvpzCoa3iZc4W+JB
e0SmWVtPg517f97avmC60vu2GS8WR7DbYm3uNMkf1VdbeJorbIlfxmZ7JkFAHCaI
Ff47w5rGTHMWlvywvgHlkNu5ZhULB5e+RGqa2QXhNXsNNMEp2Yf19+/RG+PqUWD+
bMmlOSvZunmPonio5jJEP6XpYsMa9DZrjD0UBU5ucU2GOO0QkGqHeLXXgJWJJnYq
66JVdWI11qK4u/giB7vFTNYeR2gI/r0IJRTDl5CTxOKUUFyZ6ZyPkgHglPXmGJyK
/FnZuHaUcCj2DML5xgg/rk/OM+FQO9nlZECKcxK8YV2UK1gGC+lzWLM/MNrdtkVE
cLT6riBK2pKBfYyhnNnc6MJb1yYZlZT2+z0sPqJGaGO6EnTkoibMIte+Qnxj45bE
1iywYoEBsvMz6U9rQubZlATr6bu3U+4YQl4DSjSqU3JuyrxMbSWqaTW1UqNjeveO
Wg8u8ORSTZYHZq7jqGYwDl7aZijnbn1pYzd5PwwqTx1/In408ADtu0A+NVcHGZzx
67Pr47zjqJ6cUDC7+NzMLIkqsbX3BNeN8jgUdW1TXR/AEcOryF/RnTZDOeDEcBhJ
LiSs4YV0R84Y3Em2aRFbT210RersIhKECFjhCkbrrPoTQkZes0xe9B7Xb++faVqa
oaKuiyYSH3qjOA5z/a4Xpwa/vYt63Gh82nvpqR6S9c7qh+ebFksRfpyDlgYTLwJq
7kjD2OpGfQFA6lm9IAWPpJUhAUJNKVtg7YshGrpaDxCRWzIV+963Wj5YD/b465qi
+kKGUcfcxmeopC+Mu7Ud8liyUfMNRX0/+0s1roEqHy/awLvEIguYdYA9R9tiED+K
6QdSSK6hMrmPGaYooRHNfKe1OfdueR6FBohaaVlqdB8egIyI30ROjcBti5Zf/ITq
UvLSZmwZNOkCpEBZx5/yv8lJb3VTl3um40TEA9YRN1rrRPrABjmxrI6xWDjWnITI
tyc/bW9JwTobA7E95vu06zJ5mC3/RNh6M13YB+4xj7XdZgbYZHiPHX9wCdwe2Ekc
+Zb1q+O0QJnke86SWnsYsz2fRt3ZEtnAZxDWvmD+/P90lWDP8tme6/ZCEl7kgq+Z
rVxnijEkd0I0+jIQRUJjIOOBzj/Ch67nRjVLx6ZTcKyPu3qThmcX3+aijGcbLO1b
UlXq2YTOO7mQW3mhvSt6nI9El5Cc2KICsTgnB98uiG+YomxqpL8sP/+hDL9/+ajf
fV5cnhq8F+mqFlEOzDh1iIBOErT+C3uKLJV+9iGqGFyf1Asa00Y6jVa51/2Cmxrw
EGtKd0Azw+/k8wTNVr1axd74l8FjXQdYbbOCqmo4Z66pA++DYlJUFmA4Umtc8Ul0
OX1tEZi5/pkkOdEg4AMe0Kdn1upnMBuRVRzKe2WMP/sIcFKVRTVp2SY8SGDy9B8i
4HG0ntCYMbFP88CYXt7ovdXIaGQHczXyNN8SRSBzTLKGI4I4UEkG6IQjPinHvugG
2oXbxWJPFksewmA9j2oKkD3cty7Au0OqAqPOB7SKnVG1j8QqGLFjVY+HSljLwF0S
EzzPj9nPMs/qjQXsgXy/G8OAVQdPStHxZ69OWDjWmvBHIzh5pEbcPZrZemCw3bDM
5UqbQcQfpLC1vsLMBfck+EPovhzGr62kzCDTvol3eZkSSnVLJYd64qilTkwN+ND3
D0x0Ow1NOIX3hVKd5RZqRQ8D6wNAX3miBOYoXODgaGbzS9Qq4yyYTI8STFKlDVop
csuurXiOSGwivqEFE0E3ZoAHbXuA4bqq8hKWA/wipm2pj+gV5Lj4R5U7GQR3vMCv
y4FMRrgBVpobLf+ezrUJiiRc0T/4kmOdvxMXxPt2kAkT+Xovv33oCioWZVD4swUN
L+5hweHRFzCYKHZFP/VRyKdCBslcrzP8RAXIoLZMH7J9ufMpYlwsOKSUoh6bfN4P
lY7M1Qkkuhx+ziaIDkG/7u/3frB2tobUSH31tBzus9tH5N3+B2Q8i60aV0qAr07o
ZzGcliJ54Qx93oIaqfSvwGUkSxccy7rBrjLYIUVEzKl00k/ET0r1t8eWm4oFGo2x
DdHhfyTx0lFrhHxHDSdo/U1SI/1svTJGQ5YDjZL0mopncRw+5OlqgWT/Q/Pjo+BO
zFyHe75pGDt+eVRLDZpYdy0482yiWYiK5DIey3Ekdjk/33pItdwZvabxSH8u7Lsi
A9bn12eb7E8MhR7Fi60inHUeAvzEF5mDbws6vrRuAp+Ceqy08nCPfFb+AtpuKjfF
m5PJ/50OOQEVL3GkaxU3G/mr8+eIgQswPsSXZIGXj5jasvv0n+F8gR7T1drN6T1l
DNfVtxsDF2FQkLF1jxK2VJd6ELl0GmaudcoKGi94tbGUi5ZcDNHb4OjCEBDbeiuQ
RLNKUk9pRHkBHrTrAHHeKyDuQQXd6EgBe7dL912R6IbzwWIReVHtKmMCp9W74v3p
BIBV+PvY2B8mXIJeYBmlA6FMTyenVLI4RCfoscLJhKdE9OoMZjrXo+NbXN/vsZea
3upjSbFmerIUWeNKUPGFWzOAMcGpXTLru8cR215vFCJGtpu4Wl7KZrC10VB4d6g9
RxWJkx3yba3/qb7WZADj7O3zslUP+n69bbV75zF8eEwGq4q8H++2JTqfctfl0UXW
2mP9Tl9L9Z1LYmsCyrrG551DThMrtVLI+opkF/wiuG/qtmFanVD6MTgqb8Zoxosa
93U76qYqp8FUXhzptFUlw6ND0EkDt9QQshLWjsgfH9y4YszTTqFBg6qSlsph3fbH
MzLoJH9hD+CXg0Z35I8V8wxPia5P7Xt7qptOPeQjggltHdzu71L3FUgnom/nPh92
R1zkV/eihkv/v2l+yqgqL8IuFPBujMM0sCbmeqcRQ2jci43McS5vF6Qd+yq6Ai2O
Tb8wEmL3fYfqbceIfcUNt+cYzjHJ0F9RM2stiiemN2wJdSl/qilFQOaqt8BjH2Tw
+towguflnfIJANqIZ1QYDfbu1pfT9cYawbpNCClQESrIlARPIIz+TW7ACR5fZ1y+
YruSAIkdxqY6UhXW2qTPIPCrpVbPptRngRAlqoQ0nLp87NPP/fr9QEIAfqpLz3Un
X02QtFc15r6/QK08tpKLGVxYiDE32VtdCsST+UNZKg470VhRccAs7yugPdfpezBZ
qnu1xXJhkTHBjD+e/se7PVdnpwpXycSDWxbndkic0iqwNKCnX1in/DrypHkM+Op1
OeVWpzibh31y+TYS9qnc8CraiTo+4o5gs0LOkCfnej4jruv8AQ7Oj6IyD+BAAGl6
WtU9WZQDHAiL5M9KdERSUHUgjfW5u07XtamPfWtu22Z7ikVl7unE0b2zAjfeXwVR
01N8PPxLp03Y4Fl2yKFnXfSZm8zib25l+NEXVIuQWWp8dL6a8cVF7wYiH40kYy8M
LI6jSmdbGFTWdeHpBWvDr1ZTIG1Yjoy7IlH2zBzfH78xrECFZPU737YAeNuJjGx6
0kmbKi4M8YLJVStbT25wihGo0U4rRCCUKuQv4rQxlJYIfvZr4RCQ+W2zgjsbT2PS
WKnaaMb7sWXvvQA+uO5i13q01UpczpcRlDI9owNS+9uuEFP258fOKh/qyAZ0pWKe
BmD2ZS9/QRemxjOOQ50o1JMlq4NvEqWkIl79F/vUBJNGNQFueaTWF/BMIq8rJS7s
MtWeOGx6joSmuM2hWZWM7HPEcIf7Jv2eyPzThcxxy+or8Ms64duq2v6IO4SIJ+H9
jlc5ry7719N0AdviTro8xXPlwWYFQmCZUOJzl2PB3hiUNJLAn6T34yQG/TCur80h
mV2mPMLxTQtjYcYQ7ofEloYb02dvlo6TTf+D047AxJ9m0hMnsKXORQGUhilv+8iP
XahhpbYRzVs2Jex7YHUecNFpSqcx0tInh/crQNfuAAe94OQCaaW+X31GYzJELuXq
9+z9omYYlaGAzb67TTzLwRnItWPCMvVmbvFWiMJVpGRq966SbAt/X6dJEvdKr+Q2
8Zh+0nTINOHiY5Fm1/Bdoi2hSGcBiMw7gMDwANPWELKwXExBYg3MHLvuaifo4uSQ
RmB5mTWWsdgGdlGHgNCa6XTXHIfn4neJ0s8kbM4H2T0tjN07/da4eWG35yICu8V3
Za4AL3ap+MocLnVFgPALBuUEeT2ThHRKNLuxtNKz8wm6UrfdSivTjv9DEeSkT38g
bYS1hGgXCV8bh6sXpIKjzetdhAdgGHA4XP5fctkczpwdBno4qe3NIzf+q6aRfIiK
vSZy7TPYrb2HPUKzBKa4IZeDz+XjcBKju7PPKfbvsFbocpN/boQTDXpET7iObOXn
QSGGQfnXW3WQgWd+3ZABSENaVTitMgUS2SztJ+cZh0HJDPuskxMCzk/qFu/+PXpR
q9toLUhj/lZ920cnk8v226lw+Aese8Cf1apDIgAWM4iqU5/oJwQRZ0ksRLJoqVzS
qYEuxF5h6Z25c6m6aerpBt27aWcHS4Meo+FyvMJQho+nRwzzKr5FECyyclX32V0n
0sinca0VOltYOLIO73jSE7Z1n3oRcYdsKRddzq8/zwdSQAwkFZkfpj2r9S1Do5DP
+qyIjelhiHPTUC63Qy9uJNLu62n31DtHH8Os7W6zFxfgNmGG9r1eoOJAfYbIGzQr
2r1/chqnIBtNBanMgTJUvw+AEhTQgT2r9hUy56+myEQTr/rfPyk4tWjSi8Mq/IBv
MkriBJcjkfC01P0LgEaPvjz4ThJuc/WHmhFIlQ8ELLf+CsRkFe96xo8Lsvhm5H2y
EV4UXqm3fma9gjUnTJJ4P3COJqc8D8nfBPeKu9hG1DCT5JSwG37KaVG/WI9vbZjL
HzmMJKnkXHS30Fzj3wgP+x52U12Fq+3TNvHIn1iK+M6WYUnaD4weG8VAs6sPVnWE
LIS/age+k1nRC704Syec6ya4xfy6PGm+IuIR8aTYglsmp4x7ey+LP+HBiyt8Dzjx
HhrlZlFtexaTpEvk7pPIkP7gg63uNd8KW3DZ2iUydfKtkg+oAByMmsAu9QoQeG3f
h55KtvDy1k9i8QCHwz6cul4yI0oLKyUgJJVYtzy/mNClhLuao8iLPmjagmZ2zhMK
+5QenZ7cUR6SqIqVNIQ335ugsG56SUFFWvxn40eSWfRWz+PPu+CMlXB2TyeRgq9X
ohg8KTV9sj0kUzRUsBF3VB/mjy3piQFggeN4nYOHJ58VebvhYBnzbAshnbQrAOol
75zQK2CiBMu2gFbHyL1Vg67Tj3DrW1RdSma57CgOwjtn+ImRTKqA3zL4tVw2aWBy
NWHP0GGssIQUYcpXffcQI2Zm+0IVfdu232xPRFur9WuToehi+BC2X4ZylnEyI5Va
olNyJAP/iC5vdxwkSdhEb8kbw0u/o3LySM6anvdZrrcO8tJ7j3OpUuJC+XQARLaO
Auj1IvIE4+OCw/ll+TUanXVf1aWX3kwEWvgQN8OB7WzExUy+AaVA6LigIZwvDJp6
/9JEHaC2izTo+uNcRZWsASWQYMg0kZg7mqZN7qQ4PlCqHmYDB1C1Ae6rH9LZhaw6
mVN/XQANevpti4vpAsHG1F14yfIg+0dKZyKVF/F8NvrZDd2AzMzIWyEWVk7UybzV
uFr/+vsfTo3SXry5UJgUMDhx77DMYkJqrTKlYHVgTQC28YgAB1olPJ0/n6+YtPeJ
BkvVx4yWKNWijJ6eRqqB4PsMRs65Urm3l+0YkxLLanGniyH66qVZ1nZiDsdaSxJp
fqkehAwRkdqE5QWcwRDTUk3XPBH3rwLakOFStYr4nKCHj6Tq+6gxW14fla4RAYx6
J0cQjIVJ8ksKh3d4Q/68XtKIAV1A3kNezhNszCpzro4GrjM9qdpsHojggKa1HlVo
114SKM0n9y1TQ9RUXuqlREz/MtUqBXBhgJvmSPdFfuB3s9GpBamUpqIyR9F1WLQp
pyO0rn+xrjhn+hwlpJwgJhpVw6+8yw7GAkMqCiPLgd+4Dv+9OlQlCEVyL9jcKSjb
UD0l05UDEu2OiSV7MoprOgnUouxgOypFPUAPFnpYYMP1onYO/lM9aB60cw+G5wN3
B2cBL8IUZM2Eal8asN6aZ6417K+zniNsBA/FVW/yQL8MQ2/Vewwqnk23ZRg/dweh
Zg+drgYzSB4KlQsa98W6q+DmqjElBpn59m16ef9Q6l+KA/ql2a9Xyun2hgcTS9s2
X4n/l7FBNsSNz0TzuYJDNt0z6KXZuVKFnLyLhnfK6FICr/yPEKrJmSsmOYSV18+F
PEcXFiGRJdctTDMBCTfm/toXxgKVtZUjeEUMqfqpjOerPMIKL+0imWJWiwRUzvoA
939vsapBjfOlJKKZAZTOGe4xZJN6fmozTbToxpLHvq03I2cIM3X0nb1cKzvSnY76
me9A5K0c0zXeWZUK2rConzcEu/xT3C2n+DyFlkKoDJ7DqyLHI/MRPn6y7DqkfvwC
C2n/ZcMWDhHhZvGjhvKqgetRw8hbKqt2TPJN3FcwTYsaCDPAk1Iyq7QU6oa0OFJv
tOLDAY85tzLLBh9cg5sNDXzPRW9uh1pe1MzUtBdWUoKS5HvN86hi643AT/t8nWyN
saSY/v+HGbLoR6q3URtHQc8XnzDXTMlZ/voOoZw6Z88LEwCQzHi1kgLvWxWSIasM
z5+9HkefRL86NEyTJruiufJQKY8IphI58GkeCcnv6WDLc+L5eU/0T77iUOgxTKJB
qD2uoxZBk9DVz3GRvy9ZHaEVcBP+vEP6jD9cbFiesQHRkHV58Hqr2/UlZzbf6Vka
f86wxT4JR0caROh10aDXtS9hbzNZwuoJ+YAFtgPapw+sekRclvc6ysyfBQ7ZKQJ9
JJ0bcv7Z1kZ4mhKZJKjARKq/7EtYU9FFOdP17f6IvtcEiMt2hiN0GsXID5/RKN9c
4wkvh0/AX6+yAMTvKddZ30pd4EDogZQMDry5b5inw6AzdOhOYHG0Fl9UOOusZPDH
gr6T8qXxqt8bzbSfywFnrmtZpkKKDjSb0pL4AmQGsKXKJShv0sbTyaZ+p6qFDXLV
SrJvxC4YFKU7r87Eta2ZGAM68S7p7KHJa97iZlGVFxbsHWkM3pj9zgJlXufVp7yV
Nv46r7vV1hBacCXrRMp8R1ldE9roJNz+hYd6fqLU90cRrbEUoxMic173QiEsECMr
/7XyTxUQMjzmtYdMJ35HeMW/GTBDuZ4Se/kRV9bKSuleyNUmMTimrg4N/6cehmaW
a2Hyyh8lxEmQlox57X/r1vJZMWwiWlM7Npr3fft3kmoc8zwKSQ/zm/xiEr/64jtP
YAFH+nt4kLHQ0mbl5NEaNz87//NX6X0/AHZjMap3csNfW2yzwSTpPo9mHEaezgWU
Q8qyUFoKuFFnf2W6jLxyJ50rlTL5/hZwFYNplIrq7XQFLI8Q0MlJ/cYJLAgI35np
pXdOGTKcReDyX33JEjy/EG0S8MRhn9RDzjNT/aQg0xWVcrqgSf8mxT7FKkufzYYw
ZF7f+b8pDjrYWPZFKz0SHXNg5bqVN58vwx0pg9Vj2gvp+b/pI4d4FmWETLx0t/dC
MQF7uXIaSBlw92bEnSb+b0pQ8Kc7kZuaCWXOobfyl1LM/mRvdBrDLeqNk3AbSrMK
C9KJisnGQYhNCTow4BBO65lX6X6eJPINUXFB3On+qJpa3MN2PmHq4olrxzRHbumo
+HFwtzZgJK1Hp2xfupmcBLskCiH8MoYdg3TEZXf0vruzFDT9JnyHoqC8rfiY/9+N
9DSgGrdkR7S9o4m0OTGBu0J2zR6PZUvaseWdWVirpcrzc2SDADJ+eRzUGjaITSMw
EQZzfNnChHqsOyBL/V1B8H62EI6QfenDMY4oT1E8/CTTEtqindLIxGb0MgB3Zo+q
+TQrLESyfaW22ftRQwTqOtiU2sVL/sfji+RFR68QQWVUEPYbr9i1JeBd4yYaIlVh
h2COzpNW0/K/kjtdqQ1cmwTiHRIZgdokEtdTD6VR88ac+hnxKfmZi4T+B/WQPn+Y
l5v2gl1CJdl65AYf2Gw46BGvsh0sG+SsDG4fmluDOo9jBoyWGjqbD7+XkZzjvz8w
hSCUF31KxMuDr2iGN1ntqEmTZNY3S0exxzQTkpMHTxTsFCsOPzWgenpT3xg2kqmo
1/ufrMgocY14UNFQvUYNaKQV2JOc64Qp2eQN6xDVGkSy2jfcPS6pSxyydMtCnqHO
gcyQus7RQYZVwE3zpZ4aumXwSPnCks3jEa1phhrJPnAvq0D6F1GQ6bCnwCL75v3/
n3weCCEOGgcg3tFgY+1zch1AW4PoBvr2FeqWQiPI8wI/yXwVfdejsi8YGh2t3v6p
ooV1DLtL1fn5yGlqGWxQGRIJdS0/R8ZzVGyxTFk+uR56hG1LcSbHnZNa6O63v0ch
uAelvlkxK8gjHeAhegVprTg7loIN0ju48ghjCxPBW9pfTdlMTZ06N++U4yYQ9LEk
BHDTAJnGW+rpG5bINnlzywj2gYk6oqCyzWTKbaotf4QkplhiupJz72H6aYosQ4SA
SCCUj5tzwc/D2PSdDMZFs+IRoCROS+SOn0ec6QMKSyMJRenwHeE0ovOvRf458ONe
VVLvc19ux0RgdQXX9z5d2wW794yQdJLr1xuVkReHXm398rt1iRfKJVlPKFsigwzs
lkhzeNS/doAAUZm1vBumUooXp8HbrINYj5tNVfXm0W4D+PHMR5lJ5Sqht8iEGaUD
55YIlhIzwbbTU2RqOvpZcAWsd7j1fxLSci1I+Fo2ktX852yW9BInaKX/D+wHkhK+
dSuuHPtJRSV2ZWIU5HQKGFsLGO0dHi7k5ryqGz85Ie1DlV3LXpPox9kn66UrlZjm
v34bRTDNhw3DALtR9tonVRPuOO63kuUmf+JhRYNgaNClEV6X8PD5sWjTfHAYZeZh
m8jdoG4aJE7RlRE4YXzZ0RYmODPyK+HkvUNME8E5CBcEKL4wufGMhSUq8hJ38c5Q
wNsYttDjpZ0gPxDv/QZEtF5+H4x7yQNn7vWlM6fCJl8Vowe411ro7nXDIvwuwsWE
6xrCD4TyT4g0DwJH95/bwGb5jL/h/y61YSvQGaYlaDDFDwXCTj1SQ5ResVM/0mrh
axlh7OtwF4om19eoZXZqOfEM7ofLMbb1FwvtR6kqPF+efM1I5Zagp9caEMKbVM1g
ZaEfz+/ENHeiNoOHwziU7pUJmMABgVZeYllVSXQIA9tFwvzZrC7p5RaizkD2dYNe
T6tGUcL7Qp9WUxF4cTlgEhdwWzK4gQSibOOTuEFxj1/n7wHzxUkuOoI6SDmJNlqs
voADAHoUJKSjxFOVNm6KvvprhFCbip5Jus6UnG39IjaHGJ7MuXOt6ULYpT/rx2s5
aOtJqXUSAr9HeqNEeThc0kWb6oKZuE9nspPnF+kP9uLI8d6DHVLb3Ho6PsYJa12b
qcc+MuN8E8nNkHOOoTWhoounfBqswd3DpgqBcuJzseVpXO18ivtUARJ9NK0dxJRJ
EBl8k2MBU0qxs+vgCvDo53FwQxIaTkzjcwrIswr99bU9eZ3J7ZqjsTlXyoqrcPxt
9xFcT0+CP25MjoJ4bqfVZBtx1Up/KUfkYeL17SCxvQVhzT1vFjUM0wfxgc7fPU4s
6ByTpUKhCDv2MufnrRRdeqOOu5suJ5nSQ7NTNgAjTkuyyVMO5EAh+69dZosKcwk2
O6LR1m/paJNJ6FIHqA+1AE8GvGeP5olrCAlXbDC535G6iC6gxnEnVVuJTPZ18Uro
91o49G88tNb47AqtA+tPgDO3wcFSFg0EkEsmWrY4lHUHrn7HFOx3IcPxgdtk3fOx
FKuwHPQqjJbVlnlukYBCoVA/iN+LZceoOXj6Zb1VQe+B1AwJJiwcJDERniAu3871
C+jOsdVAc40K2RTCXqg38OybBXwcCtQGeZ3k7ob5xv+MByHuHaKqroWAqW5fEHbh
25SLlg4MS3WZLQCO914WnhvZl5NTtkDfBljDXB+qGEsYQLwvCIAyejB7qHkP5g7g
LrLEFPMqyboWl84Tzp7Me1Cus1BMbF75FLfLZSpRqV1PRaMkBmCNLS/UeCB/sHLn
sz/4ppnUUBua49ETdQF6wQCZeZ3V7bpNZ8rC8L+CswhS5eA9Gtm6EYRT7qjJ7SqF
KeGuliYUV9WFl9Hk1Le7oKGNvSsX+EqAltNF31hMSCc2/w/DHrY+PLDrB2ecrFPD
YzcoauzAIIalWxwKEOEeOBkzNbHK+uP8x07TFAstAkyEo2EmYufgfKwni8fgpDPw
dIOuQ2CZEXjV7efOBrKi61xu6mp/qWl9sP1JgK8j/zKy8cjD9lVxf8aD4XdVipvc
OC7tkVoqGKa0j2MFqAb/E9dMf//qlSH0vcF1jyOOiy5qaPg+gz9kS+zQkkjqv9pR
UjKhzV53acFupiM+HMwXCxKbYZ3w3/k+cHmZ7vr/hrdxqhLPeQRRw80166n2OSAm
WrMIwKeQXXAmI1XFns2QdbGoS78YxCQ4kFvu9Ip3LqocdfDZIyAJWYI24aI2ptns
6BriYEXNOjlgy11hCR3ZLuOJ4yNkC2LB8v+Hwi44T7OATpQV2kfpiqkUpU+GLmzU
NsFNcemD64GUQjFug41CAzasxJB2w8eNKkBqYN7b8nCrqA8QmZy4a1R6m4pztaXJ
UsvhScklowPSZHOSJWob+vocAtgzsfao87jSPDiuiOISBallpySSh9YYWpOrXG7+
r5oiUrEml9Qq/NkL/BqYF7wo5mDdcwaRqkoRXdvDML9BlWuEABxFg0B4biMO4Sz6
jyz2z/mpTn7MCz/GpyolV3L2G63v9vnWhOwGCtMLhRSZ1EFJa+vP+rlczYxOIB4Y
JjMIB9VejtrU+AQbKjFBRTDEmcJzQq1acKS4/4+WWEfCqJFqIgcdq/vas9mO3IqC
eihT8D1fhkHGrv9oIZ9YSIfCIB8ZgptO2b4KOzHJfIcJW6q2tvXsV5+aFwICoN9Z
gSphSOIUVQ2hQ2bJ+p3OHSlVhjQcfk+FZmAPB7k7eeNYsq/yr6yJt13S0lC7eTj4
NHDTl45VsTT1BBLEEEr7tsd23ecNH/pirlQPC4wFX95eGz+ZySwLcEUEFRDQraQX
vg3xo/PeWPwoQFYgc6muE61/b1kbCJ/okv39oM5jIHfh9di8d2hrlXqqhKnVycPi
sFkP1fEHA00tfpKJRwqPdAFRzKlGhDW+2sdx1W8+8aCQwmf2Nbsw5crfT0fuM0Zd
qtMbYsH3n9UrdXrRPSnjmXcZTZ4mmDGW9uparqmL5x2ZkSBHZbFus1Kv1zPuvxZU
+oV7fhujHJlsfu1ilV5BChGTXN4RaLQ7xjyT3d/LvZpOlPk1NTyJozCakp4BlKqi
J6nARHmnVeDMuIVAUriUErM6ptOM1KE1Qkudb4EMvSKOXG3rldFYqSvM/MHPzy1x
fgOQHskLHyhFg5JuVzRHeG5aWEW9irakTJ03VJyR5xqH2qPVW0lLA7veBuPJlKCr
I5zBV1u1RJzXV+NJeWAJpfwPsW3RN9q5M/Eob1hzyCibgdOYqNK8vW4mO2vV9PA3
G55iour0qY/ziXC6rBodCj78OejqL14tIvZ3QveyiiXub/LcbNHfrfteo+j+apWU
5EzTn7mwDD8a4vfy/DTrhNyVlUvWq/3A793bo4fcN0AIVIHdN1ZKfSJZ70mvQb7g
VppdnPmGMfpnGN/+mAJHTuJ2wG5TBlyhUCKQ7u4OiGWpOdhngdddh4s99Vz0Kowm
GOk+3EGy/EZkVKpZ0qYIbXKBYW9rdzbhRk6qiuxDwGoznH+Jc9A8H3pJ5U9IoO5n
MbdmWmLJ9lIL3H6Sql7AST8cjt2lcKu3nVkrc6BqVEPkyN5hHDUF7YzfcoQLWTis
y7Oi8k0Ghg3sgE/7IXhQe9EATLk0dJjMBprtbEWjVh1O7n9QrsrxPTlqPejG7m4a
d4r9T5XOvGnBfuhiS7SLFcNkVTLJzDL4f//k6jXTNaXFww7cbrpyCbTMmEdHCog/
5hgMOvRkbYU1Y1TQzkXEHp5+Mj2q4/kucFm4+0U6u0xwJKJv/2gp/SbT+CXTrfy2
ll+UDWNJ0ZoDBxsgV8SaTbj1HWJ3TOc32+mBK+x8cTEfuqCqcCfp0ec6bIjQ+xSq
TKtx98n3A+qDRM7qsBaxGE4Q4CH1Ia65nQspW9DWHTKSiThA11vMRkDPfr53vZgO
ulkoT9en0og2haBtcX996zHkpOynW6ZvNfFentK6SI+77tsY0Ed5xW+IJPWOtNDG
MQxggCb2iSl713JtOkqqqziDrRxCi/yfUB8J0LZaKMvVWn4pZg8vzSqgK9P1AeEc
zJn9gBFyWFVDNogrmx5sU7PNzRyaU/ycgygPMv6Kzicsl6zucPaRolciGrKnc4Wz
8JU/z1HhOrDXPIYUb0BkbjEPx4z/loN3oUs2IYCIwy4m8xbJNE5Prr2qCwAcJSpz
wiLnX/QmhtslLoC0v2gh3hKAXCezIAQ/bZEgSTXjIxkHBHkHxljpRO2SRDpNEVl2
EIJtdfZxylCjpte3+MFy1K/j1MZ98RN4x5Qv02Dl00g/R9WGYyWCx7mwA5R678OK
72jh5BSO+Ub/XxMAiJ8z7McrarAHdQUc4VUdSOOqOIzCNCFQ4XO1qbgkaAaBatUF
IJI/rCCSLLRiFfs1TilLCUGt+NG2gAlVnklhzb2nBXfHnQCZ962mauWn2TEk8ybN
Bfb7i0y3SOPGYduzqvoDEhMpBURqq9vzLaxkxE9tLieyLVuSOmRAyUVqBQdt8qjz
kPskdXkyKM22wiwUqe07sNkoOFZAK5tZqcofBC8MdfVQU9IEQCAjvTwuG7JEdfGB
3Dq2m4+f68qZf6C8Jyz1xrReYdh0Jpt4L3VBn9selU3UTXcHyr5znvOB3PVb3uRu
m14s8T21Wvtdr2vMMLETxpWtIJm0nGhZaHMAmDvKB0MC6hvxMUR3LYwJUr9gOob9
cVNfoIYBbRYo5mKpEj7b/SvnqmwudUHkjycwWmcuWy34OmH50O4/RCCLqLd7t6ix
mRdYPyQPP3ttA1qHdyKzPG31lrjCETNIflWGdS8CeE5ykyXTsLy44QGeyaNlQB/d
EuPHj4KqiV3Af7gJCYLkosGN1B1cPiNoty5507FgbmpgIYrMtN/11KrMsMvD9CTp
mmTNCbOLsxv+D8U6XNbMTa2EtRClchvjaBGQAVAfJoIp/fHYtMBrH2a8QG83rxjU
74EjcV05fqWhrCYZ8/W+fRqK2jjFFeYbUWbFlM/UB1EuZ7A+WrsyCQUqZBuduK+o
NmdbfMJwnx5IE6M+oJcCpIeuS9Jw9+7Ys93pEVYI8m90/XMpNJPDUAD8EWm7I0QJ
wjFoFGlslDsCUynDb60sY0rJ0tsnoS4F4z0/KcG5uin3bLpr9O+5bAe3vVtIElmU
4xIg1DdPvqMfvTMrrPUfySbmaK6QCCzGCTyTItjRd0fUyOxkD85ctPCIV1TVoAm+
YK6njoBXUJiL5N5yXRnp/6tQXJiJnSmg3O5o+2Qejl+F2PxFlbrCkcLbUv/y+xTJ
d4XTZu5eohqywNx43qWZQ8PJB73mP+dbvdCi4Pdikpaz9WI0LhsWpbS1iFKG8rqZ
wxekHNNcN8tBxB8uMvuHEq4ElZitNhi/jWsC9csT8WHYWupJslsyAGXFCDw1gfJf
sA3nwJ0obf4LKQAZcaR71DS1IUo20Ky6Zw3syHSwG8+UN8CAz2jkgnZeokEiRLii
Id4nllR7J4Bi54w0mPwGuWUTt1JB5kLiO4iF1AUsfD0LxvmXC3JMKsQAUSwVoQYK
KIsic6xW47bUI9KW1yJOMgvDFjLWquv7iXAP/OGRUgItKmn2sqKew84g6XW9CZDz
TdBEXT3XDBIWxIuuiq0h6ygTP/rbGGAv8QJqJ+eUInUr4aB2mDFiDeSQbEuFdK/i
2zjU+js/fI9JF6PMdZ1rWZhW3AMLK7EH+INadbUpSMRUY7eNk8FjSMSaMw1/qRpO
DB6kJl3VKZ/nHTEK3405LQOZSJglE78L6VQV6+/hkzgXZYCVgdfW95ttVFN+m7tL
/UUsaceMGBU2EwZ5GPAef6tHh35GYzdme03GOMi6MuJu272/LfNeLPNFWzik8VTT
kyqbxxWKF9d6VYYR5CbM0V36cQjiQYq/5CCkZ0N4suop9VJxnSNSBKw1lYaNHOyg
s3GpMOH+q2FqwbQhuKE+jb8kUSm3Km+DyDoV3h/xKkcTtKzgvmgfTUuh3ZmrM1RR
M0BIlxGmzJ1c+EKmIjJO9RolcmvsaqhdRGpi/wINWQ4XJFrVrbe1LFyTsKzvBctZ
UjrfSA9v1rO7kjUwpS7npMhse8c8FMx/43ZYwzQbuq4MTbv4U6pVXhRHVTcy0Zl4
Aq0pZSQ1Xi35zSHrPBr4e9EoNJ4+SEsi8fJOJSkUvS/YbXf94X9d5bjq5k2Frp1a
cPaIC4aRkWMorempLf4pNqybX41MnafxwXuXnGasZJdaIEnVXwQvdyRBkStFlLVG
8a2S7bHcuHOwauL4+nc1x26DlwtxWtIlrhynxtSsPfXBEH/IqtmjdgfVF7SrIwR2
i1F8ggSJXYwPubNrWuIKTaQZJ8izjhO0ai582Y4byNGYNwl/KGpw0c2p5gkNuB6R
Rq4IJciYH6b+U/TuPpGACMGlQP2DPXAUfDg/nn1GsUwmGUuEkawvAnVAINKDCFka
5A0QIi2qqkV58VT7OLX1lbAzEd2lChqVQ0YjqGY/C+ydpBbcKobShuvuHFKVD+JS
gZttFKmwoo0sVe+PLKPHalZjf3fCEOHpM03v59doEcFuQVY1FefiKW0A3Enb2RTn
rfI+FHuIZe0SjYOy6e4GqT0qmmnXHLv1Vrfk3/cJEbdpZlLdYmbeLqLJgjtqOWpz
1uKsJZ3zBOByk5kmkYobCwOL5/IIT+gY+wUG50CATZWibIi57KgGKuB5oZt4wnMa
H+25J9TjpxflU7Z0bQqzrKT2nfODDXMl2VyC3PiPe7ErNs5QRVRVwaRy/FrMV6X5
WEUPMEjnDRWqbdTQJHIHkeMmUTWaFaWrubA267DQ5ZRE/hr+Jm1OHwL0kPNf52Xd
VkdZ45BojdG904lNtDDCMcLlnbcQ091/zJKaYhKXL0NmLSRc8uHiAKMKEnxBNA2B
O4kHdZTczXS9iiTpYLFFUr/qfVrxsNhVMMTqpEK3EEbIPAF/tKDFprEaRbQ132FX
nv+QBALqL1Z0e2CmOVPHYFRbM24VkMpSYiEoMPs5zy6DL72IpNDWoyNmy4zIBgcL
yvZa5Tc2FA4/pfZ+nEvcbf0IWRjnaoBQcyI+IlN1q8z+MpYGIFv7GCdZAV+FPl/d
vO598bBaqZdXWajws7DCSlng/EL4FpKGRA7uNko90GlZtRMnb0jz0UWdSjVyTWDy
q06lROZgSeIE/E2B30Q6ifGw06GPrgqgmH+Us5AlHUfUbSt3UTphQXYhLn81DNgY
NHu8W2WjTSZPrIdr/dPOYghQpYFY5PBGSVM5Gm+Z0w0U0e4DVedV6tJTjwbqVKBJ
DCv7VhGu2iRPbRT2EFbSEhlwWc3frLqjdLKrSivO/Db7OfTAu9O0ZyLny/rsbVyp
ocUMKX4jLo0SKOmnejkgyZj665M11sctHWKamK+Q2DLkFhA7FwUWUpCIyXN7+xIt
riCDo+zJZFC8zvaMAHEpqTv+LMiynIY9DYJB/OlInQ4dQ90DnDj2SqZjzk8AlmiG
FW33p68WJuyxFPW2Ie4mj+hYB7UhtI5cihCqVwMC4CQnDcC//Tm9kRduf/FwO4C1
wRVubazOsqwCJx4oIuSF1Eu2amj5ImE5ZWGFj1f2AiIsSV7Ar8qX2UsKQB5ttqn0
q2KKUJO8fHCr0Wl/dVjTUFpr0mAff1ONtTwbaOuHomVf4kRSL1PHlj89qDF0apet
z6rknSoteuMPayri0XbEYaMNIKd4FZuSjHy+SSg9Op7hp9aYfZRmqiILJ9Gxr8bL
IF3kdtvSpbixh/e6Jari0+sp81zYQtHaby8/N/nnG5dqEoF97HlDrLDF25+xutf/
UbYODfKERIWOECZmRFr9Is16+i0V9El2LXcJ1kO2UtTxgZbJyVxAa69mtlXqXnSc
vsoHFnGuizBRlyN/osWZqIpPMLAvyDbKH+LRvMdV2sg7RAfW5t7BfqUCKeEKINnh
8O3hj5D4Gtcv3ZhJyv3AaJaTYlc0dM0QI071ic+v5zXveQKdWsLlApz0MrD6ehLX
fb/2Z9M7iM07zSShataaemuTtd2L3cI+Ht75CS1KalMxKocQZo1eKS/2OhM10qs3
VFNTPZrneNRAfXwUYsq3MtGURnfkKeseFjNHWrwr3stHVegSlgxJnuSXf+sg/xBb
2X4lNN5RtQ65zlTqJ6BJ2NcaRjwii7df+jZd7P64P7ApXBqzDbQTunoDSNDWhNve
v8SLWxu+6sM/sRoBI1sAiC+jx6oLi6Iw6Pa9W513iAkf60ARn3Otp9UD+bpG2UK9
NfkWSNE6S+227N1ZKgt5T/urUtUSkCIrbFcQDuEAi0eDC8R2XdS5ocDA4R0Z8XWb
YvkPDchkMQx/EjK6v9pjbKDKHIraBD0j0QjxmP9RbywSGZHrku/C3PxuAEs3gwcR
w/2GtGqsxNuaKj6kMmEze7gS3JtMQ9T+QWJm/S3teJQgYbVw3gf+N8Ric5iaxXfR
9G54jqqXJfsGiSp5/o1aNooyOkeRgBQ6Vc9qtq6BasbN9p2Y7u8z1xduexSqlWsc
YqHH6fduUpNOsoG/H7X5umyRCyaipqpjog4UPRUEWvJ+9zio5xjQ3Tpkhm2IQHJ1
xVxAuOBdgCHx7+597Rj/hgtkfRBYkwz6Tnw2ywcYKAlBcjJb56Q89FOVu8Hb1SdE
ROnIkCJ6dQ9KtsUEEXcZXGSVLpej5ArcCsKSW+hMjOk7yH1wUrkF+vQ5SCyXG1oP
7bfMZcvxm5mimkB9POJ/U+YWY87xtRKpm1MEEE7LnGdzvGHj/eQMUYK0ZDt87XNM
UhvuBYD/U/arVKRAXQFayPngRIiKXn02D2R5nwFgb2YAbODWJu2v0siyv7j7ikVU
Gc/f/QP5vzHHL1qvCy+j+b7f3GPxzl/o5FpodgeoI2qGf4VVTJ44Y8Q7+tEsGIiu
M4wAItB+zws/Q/DFq64895r+IUpy9nb8S9q4zWnw3WAvdPxY787jDZ5lG1wAx4db
yf1B540m5go5I/tpJPNNefWBN0EBloe6xT7DsQo2i/nzwJqFCWm3XCK71qMFHm7p
w7ToWSF/nJCiJUIDzxnQImRzDQsDcWrwrz5zONtCKeATUbvxtW1I9Y8apdR6gRzL
4f9HxTJaUmboLTBxcsgfM4I/pWBdQFF1gerzBhDDPTs5pBJMDXJpOPWvBi5RPaeq
NLhkOIESshScbLAafhKrxjhu8x5naIvYhV7LmN4HOhCU/ZqGEEg+UiEqBgM0BoB0
NmZ0Nsw3fdEH5vNoxrfTIQXqzNBip2aTNu49qKeAYDEFFl5iSCjiexw3JH+QL2vk
a+pvDidWes0gDgOhmhk8PIAVP+e4BB4zSVngNSCJbNkgZQF2E3GCsL8QVYVTe8S4
nbZ7kFIR501rUy7inGUt0AwanBjotK3wZFfSGXR3zy/IWoDKBk4grH84EZOyXpb2
p1I69GdqocMHv0+PeDcB+fUgW4khds274RdeDC91KqXtC7r2MKR7uw+exUlmxFF0
xNk4m5bauh4kCRjkgD0H+oTCTTfBu0O+7qbh33NWTWfAdzb6PakyKrwZO7va/gNk
qYCdx+ih5hmnJ3XJZx5SqppkOsd6M17wvJrwfMi0N28n9kFBva1u2VEvhdiD4lB4
EhJVLaW1PBKJPPuVQ3EPZvivhaqkkncHSVfs7TLgEdpraVlnu11X610ixP+IAjTQ
z4Pd+1WbibPzJTdwu05oKWUGE/yZA37hmPz85drnKatqrpItp9vNI28aaRk3o0jW
M5ZDuxdYYqI0QGmtak06LoJzLKpLwCe/Hk52pjWXsodwkiJRI+8qDBgjdbiCYDpU
aERrB4mErGMR3SOx57JXVVIpWnw/GZ3W0/pc6hx2UKon5TNHGARvJn3csI64Xzqs
qQ2gibILsjTaMjA+sKApdWHoqK7DQ+aFDu9BTNzaRZ98owkPXdmz2e4M3YWI7f+Q
ie67NzP8hSbTtg9pxDewUtRYBZPLDkead2QwIBK8O2XfrP9vWwGZmgU9WjmEAp5y
HVepEg94k1Mqfv84rSTP1zfUdtYlj4eO03FhHEBE6a0mqhGTo3wklc3zXWYwyzH8
IpSZYKjbd7dMXcbKjS5I9IYkESXZ9RiFO1lUH6L7+6dUHtnq0vd5pvAQAJAaFQ6F
NY1bew8HfYsaLlpURYFHm5d8Ez4nKUYumIoZTa983NQWA0vraO0iT4UZy18UaNAu
QQOhNte7fpVOj7ZuZqQf9tsJdRs8af/t34fxAJ7gFfWZrjoTnW/Pi7wXm5GkMn+o
wFSgDuSRn0afy+GHflkscVcm1RurGvuu2oX+bo4IkNJz54IBq2P4JB+5f/NbwGR7
aJ7GVgvQmdgNrMC3WI4WFrvHQC8Bjksg/9ocgbZz9+YASPQhyQ8vEf5P8kRfn2wE
Sic5Mi/I90Rd2rgyKTPZ2luoeAGfquHLOjaWM+M0HM4dB+hF6AkPxz0ZU/wjly7w
XSxVmsiXO6+by663d9jEHwBOkYjWTmfErt1mcWDn7Y0Jdq0gowZkeoi/3GnDMPSQ
QH9cWGl+nFytwVI8YxpHlet95Pr5kJIsXEUIeMDfRH0ZwjbLpEDf28RPgPpvXcx6
wqxdYATaozHErJWbBt3EbVWLBhaNNhTJaBB/pw8PVOrRKOWGlRZvmhU+tt4A7YCd
TwJGE7A20RBU18BDAlhT1twgmiidid5RCh4h0SpRSAdxTuaUHje817mXCtU3ghdO
vtxusNpUgssONY/lfERWQxTHmydmBG3JZ4BcJz/DyOXnUqs/DAjhpRXwSkqztOSo
VYoYscP3Mm1IxVPBDYOcgBqBGOgBegOeMVjeeo4FD0R0WBuvx2hvp/QS7Ywd3+D4
UIBS1rXl/U5r3xss1qa8fhOh5bVirMSz3q8rAZmip/y3XSWztmTYXnC1Mczy84Xz
IDHFBMMixUTvbqHI1SSUQUu8QpuWf7YZIuxtCTNLHmGGc01mgR3zEIumjmoq1k7v
UHd4F5ewERQJafg9vvqaL+6hGFmHVrcOzQFwPRLk1SEUxWmMEXSjtRTX4wiWXF0d
OmQOos9GRe82slmHdITI9RXuGtqh9jj6/mI0BbICMiDlb1qkcYQQBjdD2ghUNt4D
SSmxriqLHjxOVElTXO35utgXm1RH5CxGCfY+hS4QeD1zle7P4oNV0BsPwe3JOSUY
hPty8eZqHFRLS6lHa8yuoGda5Lomh/tWOK9V/zayXXyo1pImCWG3ijxzFB2PTpIU
zYoM1RqC8WGTQGflD2BoWojqtZPGU2l/6/MmbVRJyu7+EFdXOYumuuMPz59v+ybU
cmn4pMIhICPwGxD3gDjo5ZsCKITn/GPo/D3LOZWt9G8qvG91CDrt2ryzW5dGQgAu
J3RqvTHXExNvvulFoYwkflQ4aU+XW9qnizosuZCBg2YBrWvHSz76rmViDLLGorkl
7WsIxlqyvpsk49mg4zYGNTEgC8a7xKKGReDdZslGlCHEuhM6svtn1k16IEOq3vEA
/rcnewXjZqIMJn5jTaIEMTQZC8eHQVwRDIP2SE74D14w0xeeH1iDTU29XPvF3oWK
XxoUcfdo+Hc2216gtnIPPfz+SRfqbCiKP8p++edzTyrst80g09KrDGDDWuxJY6Zh
1EmFR8YBPozqzIO0FLltIzdD85Gf1pQl4w8EwggMLPegU41aDv/2OHGXJy77uvLP
hJDXqBvSaqOHBySB2yOAoZu5KhUn4AOM9dUHumJZsYFPR+EiBn3qv9C0HP1I8N9V
9yqBPVAF0nsg8bKpakDB9cTCJGrdfxHYxMCJtiqEYiVC6RBRhZpmohBK2MjB647D
8btuQ6l+1yWX2y9mBk/sQcpPZdYL7g8WbD5nKGpa1r+7xMe8KJa+sudgl1FLAqT6
2rFxoaBXxum4vchuFpShwdp8CrIu+RdmNZgxdeESxQpqa42yNXVRM9jVzS47I9Gw
R3Z7o44zkhXsbVE2Te/RydPUTCOriID5mP7yhcMMV47MAWmwwGHOUyteZo3k1eGt
xN+V0cUiVE1L1lsqKGLukNkGsXO5uBctnpJ17SXgHchdvzAHmLhsLzWygGgRMlVA
lQl3upiGPVp+CEJhiGiqyPr6GmMg+wGJLExpS3eDafZ346Y8FygGROwouTYi3YLh
y/1yfnK+BehXxkQbhxQFWY1KMtC+1cenHb4OYd0ShndZgeDKqqZw/IiJCIoC53D9
qHD7P873CzwfWzhRwgZIgvrjSdQGdScnEnb4LRHH5PHk2pc0/f1x6jYRkDo5jR5E
XbUm0zSaUWzCELCTGLcWEACET+b/kuzJHn89DRqZJXnz27MQj+KJRbMnC2eeJruf
FawrSr4S+1wEHPO/p3EBLPHyMU400h3Bjg+nrqGulI0ypmff6GhifbrCeCWUbufe
J3jsA1F6BbwGqPLaSdL7ll6ubvufhMzvlAReyLO9FUwwvctVkCTWCSqRljN3Lmq/
Au5tPpAMKw3FxAC3nTWoXveu5cIqN2X+cY2wifhTlCcO0OF4B21BoNLAagPMDqhR
2aST7JyrWOxnc1RGAI2CD3rGGccR13c7CfE/z59leZQYyu08guy8ZFsN3mVoOOcb
ol0Bm43Xre8ZKTQu8Mgbe8JIKGhzj0dWhqG+HLCazmpRQIa8i+3oZdumECJeSiTV
FEJNNJ9I+BWIv/J3OSPofH8pL1igCang4uiZ+IzGn98oWXPfrhYzsW89EPPJLQpI
TAPu/MR056DFnzF4isW7K7QaL4faipufwYHY9Ncbieh2PujAt2ws0srLTukn6H0h
FT+JO5+yTAyP/bKqxis+vDUYwbC5XEZNaZEFQige9p3+KV/1DnCMUoZ4pdNUWAah
W47JL+ELsk4E8HjnECSwiXqs5u1c2LTcaEY05QXtIOnYLqHb3v1RhtKCkYlvr6/5
j5P9T6gNIrpaEth954JFUtboeJGxnuQGMTvKjO/8GakgPpSL9yjIdPjQ66snL+mW
DkKQJNO6RRN8WqMMvOeYHkb5WSqyWQSSezMTz6Pd7aqJsMxaP6TG3WRiJYyFzkiS
GuqErqK2dNrzneHKfDkUbqBYvjTko0TdtHkrARkZREzk9iQtyulhMY5WNFDwiRuZ
OJwpU4utmycz4m0rCUkc/BVNOkxtcdW+CLZnaFSjeCGFD2sM7lh3eRclhKiNAg9Z
s8MPFb5Wy62w/tO3FelWPfKbefiZfXc7sYt8SMxUuYLkthkVPoNusghZqYCH0A4m
VoXUvbY+z/QjKfBsd8Mbn20+ex7iKXKgrX2va/qOacoD/E0JbvU9R7WN61VHUXKt
hBqHYPeE4OX0BSYdjxgxGJUy1chxVKsoy8FEc+qsyS10Q4QG23PgcXgSQON08EYD
VaDeDjCOlxzLAuPSesgTFxbyBb4nRG2D0AD8mOoRmdI/r1kFN/EV/yiFGfugewyA
zhcckZht4vuK1k4HBoyHeBSL596oECF/ieNH9C13EB/t9H5Fsx1EygsqsmxbOsWQ
/2jaTd/6OSHEWDkR/fM/BoxuOjTt6FIhccPXS1VYSveexcpD8A7McsPEzKthSrqn
pMZcp3CJD+KRrJrrlbPbjtm9XpEy4a6tPbQ/Yv1QhiBBS+To61lUqRDyoGoDU2g4
Kc/z+WsBr/u37vG9dd2PuFfvEZy5btCHFeSZf96DEVA5XY9yEKkcJVH8FFlGLzzU
m+1/691nGxIb0H1n7TiuS6m8LLRZ4Iso6uAj3cl2Wh9uDH3LtXFQVSesh93kvurO
zwGF4XiFqqFGwi4OUd8/s7ZER6S7Uab06JbeN/t0t0KnB2xbtWqLRZHSpTz9dspf
IvGb1u0YRyVVUvzYscGOAbwE2TkGhkCkcZvapVQjX5OY6WXySNPiP6wFsLUHcN4C
SrnrLurZ35qJqRwkl3neLUERv5urlHTGPW3HDeCaAH0+YzZHARzSrSA7cX5QlFus
2bvwY/E+ZABrtF9VF9nqRC1VlyKI0BldeaWMEupKfXRdMScorrrgpkLGnp9qo/xl
H2hp2hQ9y412AgjOG7PA/YHAFLOEZ/wB+/0Fr01TCA5GEragzuIFggwmOQdr+ME7
MSoNU1Un7v/qK4MlLg4ypmJAjtfNe+J/TiwsqSv+ZGwSbbgAyCPEhVDzC0zulgEu
2WlUSxBTuf9HCTNkhiBUhHhXp5d2L8WYFL20rT7vXrkokUrO0KxvDDzfBwmhXp4y
nRWaCxqBwBMHinzj1JXksS20C6M3MFEnt+Ps66zKvZ1KWLfNxzBd2jhWM04Btumu
R87y8gRm1IFl8To8pPaol95RY36WzUkjV1p2GWMv3EPzF+Cnm5FE6Gb/eLzJX0L6
wuDAfnAicr0G9nlHvQ3fRlIW2uDPFwl/cs8BsSC5zMwvjtx/X5txMLsQtWr1MNsX
GKNESI6rKeE5dhmwjtdG+Z64wQBuJFYYlewcU5mR+R71iIBuNVH4QojH57hPlFI/
U7RskBH+bEg3+4HAg72jW7o0SNizU/hN+aCdaBG+YWLlfXhSMg7/l6fvHYapplX/
RXgZfQQZi6Ih2tFnq09Zn2Lcd8xoUNAlXyJzqXa3WN4lu/CoOuQQqfXbBaUfyu+D
ijh51T46cDrFPYRMiE1dyyLTPvsg96rGpswzdowNgrAsztHqwD9r8S+MrSfOUKaU
K3guZnw6k0T6283BMqcH43S/fNQluN8t9No5E9duRr4r1YXktRS0iFzxENfXDN5f
3MvPdcaeRi5EcumHfrlAj82/1byQbkjiIK6cweA4wlI7GO/xzmMloJIBcSRrzqnG
LS9FIXD8o5iw9wVcETMXd4CHj3a/GArykrWLXYNcGpTE6oEJyaQAIs9qq01JBRAF
KCmOxd2x8p1JHusky3WjFf1O9cqT8bTYCVs6F0snJ58X/wKFHZhSM+JRxO+yXsgh
eX6QZldl63CdP0+chx5Gy5fsBXDe0YgyS4+QQcaLaRBA6kix1EfA3ot0v3EeH7ay
nwzXS0b0tbUg7XKwNWrdLiycxxMFQDptuzO1eo7mtnXIEIdTwiPRuMjWvNFn9yGa
WD8tVKJg3oF0Cxpy0xp63LN7cCpp1BLIeue7MdSeaJRyN38mF6II2ZcD0pPGpzRf
AXv1ZS+He8LjL0e+ubyvIsbBMVF6Zm6ELdbtqBL95HXg0JM2mnolplcfRZKlJ1Pe
D7e6LK4nSGWpCLde/erHcsbr80cHONvSffgyAZjD7lQKbHzjBpzgi4WoJnpMtEfu
Ietg3qm6Z9EczYuXK3PmcorAZtsxoAHRWQx8l83Q56cAxQq2xRCuWBwDZT3Ti5rV
4nLH103EHd4UNKvt1sWJ/W/Dmy9eQqygeBvjbUq5PoYM9QXFg5wAM3tKw99rSpMI
OpvVUFWjoIV5BwKNq9CqUsWZ4DRV3us2qS5MBAZizMjxzVKfhCc1Hm49hjwV+bzi
Pzob3aklHFct3rsvUSiG5xFkMBYhfjYmV91V2otbdRnGxbgQYirNe5R1VWjwtwJt
JSynoVhyTMED+uNOobzNskT1ma/Pg1CkHn2jxNz8eLzJuoNl4eMluWWzff+hGsvg
3XLRGXu15F+bzO3poQ6aSGBtpsyq4oDbcuILO4Qy6Hh7LE+5IUy4OI2eNDsvgsBD
QsFfzkpvojJkhvYL05Tu/0UXoFp+8qy3QBHiN/kCEUhOz2TAatJjAXmp5oQfWzNE
tbgjsorsc4PhiHp8K+Pr5zPvWhSeJECqEvbcp0A4sj39mljfBOScwOd4H/SxuD+B
ql/1ff/6cBdjBA6Ti1VioIXZ3+K/lnx+T1kw7YvpgIckLI+7Ji47HEbjXS/MSQPb
xa0S3Jsl9gtkA9iaEc3YOzCBKGP4CDBoqPm4eFNSqwLLCLe9P+vT9tolHsc5i3pH
LsjJ8mKKAnLN/mhsDqJwxcw4/GCrCmKuCgierJfaK3jOBYHYgTjz5Ac9kgaz4qcu
ZUGinjRpvctv9zWwMHDausUV1KpwixxCfn7V+v5hXH6UAKvl9YKftLGSKweh9wIf
ok7Y2ZaIeHZA9u+Ea+H4t4Lqlds0RJ+NY1BNtNzcdEASkf1j/crvDhWvGoD+PMG0
RuMMIBcxsSjNHbIrXFZOwIhHdypIdoumi/HfmbN6ge+RFrVOAKbkyUjwdZKnvw4f
GUh/hdhzRiCCCAOuNua6iOJV/6uyOXXh2d/NbZfTw4QnrgSZBqE+c9RUnze1lDyv
eLad/+77iY6hlqzpAcgNWO9VGUP3ya8H3wrdBw+q7QJEp20v+4A+EtiG9/iFxoK1
ei/mUlsjCflD6rvWbwoEj87GCyJDwO5dichlAGOJoVbkJf2OmQ7RKCtfuocr/v0+
+jNulpqpwckdgJK3vurfeUD36DKd03Vv6SFRNumP0+z7sQJN6DYY1Gp/0yJFiQMk
6EXBpPXJN4VmqOpTk/gfl/SBaeRJI4qU96kd6jaDPDufqzXIUVF0VdFgOdQbrDRU
inWiqfpYAXqzX3FcZQmI9DVqaXVXAKpa9zMcFhk1sgnnegzQT+nj2809mQvmKMpz
Bub3stTaMbHcmAmlD/1CFTXchn3fz0WOJnPdfcOVuyfKvMSVS/KsBRLeZq4QICTZ
mVmwHkG0T/2YozubUHvRUTv7vlgImEM/FCwLdWPCXjm3Gi7zthwk+7iECqkVVqlf
4bicX0BnQlBQBfmeBqHtw7EA1OxPRwHukiFgIdk5xgKteLHviKA93PuHtcQnpjmR
FLszkQ6nS2RyXwCmNQLxxrV8/SSxy+9m5+cpnCUEnjl3RU9/d6NvJ9iTIiSX0r1D
4o4gOyAODnwXB2Gu4jaC1ncybNA9KI3UlvqajnYcfepyYDxSYusWw2k2Etb0Yixa
fKi9FCjqceCyav7hA23/6FUaaOgdFgSg/D5Jyue01xLBHB+HwZ9vGpcF+CyhdLVt
388H4t6G69RBfvBTUD1LvOBTTtuskJakEu0Cv7+8AV10iw40GgxZbz8J+rro6uUm
zqltk3yvTPah5H2mq6AQetvfjH2bipaeTezwLv2G0joW9k+C+Xd1UanoB9DSpWBS
upmBVBeFvSLnEJzTqbw0EN38CFKcZYV9KRsWf60uF9S6rDZ3Kpvb8uiUpd8W/eKU
1M2P01n9ZYdhsrI64DrliLuWPfpqm4qDrnlEJS2vQyAehRXUaYJx97pxetgNytSG
RrimuVjPuGRmFQ6F54m7mGKIY924WZJmAiCF66lnjgMcIz9Es9yFEK/SAiITp1C4
iHARdFq6vfjC7B/b0QfwZ42MzKdCmJjnVFHzl3485tfMdSWL8MChHnghBBVtjU0v
nkZc9eRFh0+6yGlPJ/K4G8NXaqWDx5sNGEjzyT/9GvHKJOqBZLkBxwI7SXISJcLC
r+oRsypE7hETQB3WvbYKBnuQee/XNwupQBvSLv15M9Bt1rPiLZJl7Y6bA2/+U08c
IelRuGsAG2tSttUGSKWJYQuYb5Ky4lfZNRz1y4JZ1KVZG6NNFmnv7exNGY6QM3o2
6I/GLjdUU55QxETa34ffleLsvj3HCp7PXnt1BApbrkI8pBl+kdWyIvJpjnzN0Lsb
9finEyt9D4P94kw1GDnton3qhIQkkc6CWBw6VHoJYW9VRCFAz6Ywv3hjclh0sYy/
DUwSmj5VngPuKsWT5nYtgGEBCHv6t7kJLhf24L+qN4xBMTWqNjETMvDaxW60X3Gj
keh/W1dG2SKEu4hl/wQRC9UcasJpEvaR7lQuTpaDxIO4pw7rAOPGg30MHiidEVta
Ngc0MpU6aoneGCvFBM4/TW8j54p4bNumURRd7oTAAjduyy13y8GzyK1YjLPwEK5m
YfhBww9x9sqa+FTgU/z8CyfRdvrOWNwQ6qPURL3HezufFdzs49MLeAXPhSx3dtr1
QI8UHADLNRWu2mMumRn6+EOZmDLgGfbwJ/OO8BAccWN6C99nZynpe14yPxv5DzYz
/UtVHjkaRaTfgZ4KyRaTiob/MkFZgofxP4G6UH7Av7XNLWtaHixJtBfo2omVDvoo
jFrY8hTcSmh7m7qtW5cpKqRdqFH4LGfsx6QzfQnjVHuA8uHgcb7x4Rq9dDxGcCbc
cd0EFFRw7rpBsiAjNdFVpzWJVEd9K/S7xfpyiQ4t34dOjZealXRxKvFRsufZuUTG
/1lU9hHPonheb3yMLbpf8VHQi0Sevqzl+Y2oPt/d+xMECTVKmch21s3AfFBzsV1D
gWV6esMvHWBKn3/dtrwa6KqvdIH1B1tJYNxicMM0mh1ghqxWwvNe2pO9FWySwqER
+0t3u0tLKk6dw8dnNDaSkSs59XudDtsN7Yfg/VivHy20tn3RebML8zMRYYvRsQGC
Ruqfcb4b2Su5DTmv1ZYDIxBDDRtLPYlmLqWbW+6+iHtVCKz1+9sVEcYuUOh9gegk
1ENky9z2byuXJhWwUB9D9+R//P8Od350vG2qPKY+U+zZvTHNRrAe7Fq7pNQKyy29
KbgO0FAKqsL9awYVDD76xSntcrHifJj286k9Qk8KG1EIg61zR2yAmpetiwwoH95I
KgYM/+o6dwMoO2+Y3thIbhr4aeqIHD8s4tKWkiP+Oo3Wng2/sbDr/WwqZLN54O3K
Qn3k9oDiZ7b1qT89iNQcW7nYokj/PauVAkAL1c58cdbDvU9EyBdwKAPF+a0ez3AA
xP6A/V1Cfk5a5Nxz9Oj2XtEXz+dlpRY+LDneSMAwd/SGMB1V1S0tNuVHLM5JIyFH
Xp/M1RZskdlq2KYft82IQOXcq/53lfdevupk9gRzRF6eNlJdSClXQaPieGgWot41
8xzPOLrZg6AkWi3QP1NrMHNUqGfvYCkxEHdyZVV3N9COMIhNi70JnHWaymisPqNl
35idv843DJ7irZ2mVSgCNfV1oCHPT25hJ3jzAfN+Hj+hIrGladJLWI2GtDGLX86C
kaOMamZwLbSo955gseHMSm3ZnO++nsLop6ydzIUSomAuK4Fgu6P/4jrpuQIUU0UG
utqi8DUfHkGIRLSLx8hP/HuQvaWsYOqApTSq7QTrOZNf5FbWc+ej1a4SARwDOkHE
H4Yt5RMirZmumuWUxkqtkUYjcxLEEWW82rWpr4e00lRYuXxO0QpkZhKGmmEeBXiX
3cFODNcvqcfYFy4fJKefLCT1F/9al49fhVAg2yR0u6pm/ixoV4tcKMq9YU7EBo7z
9XCmuKoseVtLxPrhT/ZAQDl97V8oVa1z/gX/oR9XDpsckZqNjqNqw6fOz2AIXNud
bW7m58NRoAy98L531I10URRLpooE0Mm57Re7Q0prLyOzueWWUxpufQe89LsCsk9w
47l4TNJxfxgXXCeI93w+xaP/m8ecwkXAs2eFo9fzzdFvPZB7KITMM6hCgTWdLlQg
xWmraQ+lhsAX9bENBT147+wfNJEizFe797EcTUcqaOShJvJ8heIMNuE1JJW+nkny
L+YaHDdzWYa1NlgGsrTxbnvUTgZS46LarY4MEgDhUnDh+nN0J5Nls/nOtAGn296t
dKxf1o1rBiEibZKD4VcWLbWKfBqi2gzige+NQpPYMScZIPCt6AjXvhah+4XdNb/q
QWvUR4XuRRmNLcsLCqHMjOFcm7vYFGcaysRm3/ESdq8+7lcnn8aGCT1am29Y3gsm
1IUwN6k1Bcd1jTMBN2IgT9AjfEVyQt2NkFN0U98Pk/FTxyQiN+HSWxEd5lRlF5wl
Dt8XJDJgt4U8WNA8OwW3D55YAWMTlskFnqPMFOLSVeQ7X2bX54WwjMmMZvH4WVJL
8b45gdmqxairt2LrRSzBbN11XWkAoxUrupcG8NGrHi2VDJMlDsYrlqwvTWGEPamL
AJWrsvZDfz7X0Ufj2bUxje3whKoqGlnTyrHtvkz9NG71FW5BjgmAy/ZR16TWlaHE
svRltvAVQY3z1uFGuTxQ0NbQAqWNFDF/iuYcznz2v/WUCIWVaue0468yJpoh+Swb
lCgSoBQ0zOLxsU2wQTexI5mBJ9MIwX88eEY/Ku7Jh5K+USW5mA/TfFShIWko3hN2
6WNSiWF1+JHkwWFP3RoN/omaF+oh5hPwvE+mV7kOyVsHh3PWlUijKU0sAZ9qvP0M
XsGoovVbJcrZhBMvAnpClfbdjuXjqKGY7cTZ22awGebb+ilCl73EqJlDC/1EfCnF
UKF7RcjRS19L0sHX89YxCY0SLJHFUVUFTIcU3Zw0lThViZmplHvc0vPXxHqSobUm
ekfT2V1pjasrdVuUUKWEdnXDCQn2IBAiLQnsdfRfCTLQIJlC73oc1ReohyH4okK4
n8/AQXVcaVavK8eTaFlHJAEJPzz/oA1H1YgchltxNiS4r2ENBMtQWIGihjrG52I3
DnjRwMpw0Tukx3+AvbWuU6lbcBbbXwdUuJuGmwPqd3ltvc/Z9MB3EVPgZdahjaNq
QIfEhFqBMAP+J6els3dznhTPHaaRoiF/PT38kE2eMkqednIRpYyqNAdGZwrkZW/Z
Edf/4Hib7k9A20klxE3GYfdoXXyzq2t+8ikz2Kd8WM6u0V9eMvGAEqjLK9PDbG0F
qWx/nMsralk4yQTSTRffkUi/Tvj/+2iYMgxHBd7PDFtPiPd+VCzt4hTMAWj/NtOI
FtE7c0gk7erGaaEWU0DgaihI5Y9UQDD4ROjQTSNwoSS/FeId6ubSLOJxkRpoTILr
UbKavTz78DL+6tOqC8I2tjDMhZ975/bo30lea5+uO7DNK6ZlTx5u9ZL5Ficekeo4
SJlfV22dxJCmxLeVGaViO2SP1n/rLdL5FNmRugSIHCe59XCz6KhU4qX3ewcmbIwv
y9f+nsSxAk+YhSXVP/bT2/6rcdOfWid+sIx7Bbi4+rtiqHOLgOZSH5cZ3Tv6wyh2
IgCZedx86IWaxIsywkws1M6I3oa3aVyrQRqgnzCiABTzAGMe1MaK0cgGvyvoKTTk
FNPTgs/SRzr/5vxMXcID1xW1fhv/TLzbofGJ2QPFEnppP1FBuw2wo7gxaWsT81+9
CGMi9ZZy65Avoq2wI2Mg5JUXN8UujesAWup8XBzfzBSqKeUeiAD0qsX9GNd2Hntp
5BqaQk0XuX51zS8775atsyqJjOgdiIW91vJxC4HkHyzAX7+XBJghQ65IKv/v4hQM
/QxYlYDhDN0hUrKCfHzkk2MtkeimtpcggnI083q8yQompwpBD1PUR0QBox4Mfgou
6bBIbO7wJK9E4pnSoq0gZ8PDyX2976cEJZXXxmplz+UWt0Ks9qWXyXYkNCHaEMdq
I48fbOfjDHuYN43g3JH1Hc9apWxaAeV5AyJVR9Rq720TphpzFWzU2XuUbKu9Yq0P
MvYpizCifjf2+ldppSHGecKF9RlluN7JwoMJYfPm5CoQkTssFEnYjB9vJxC84GSi
NAhqe3JXlYkg4RIRnpMTQATdY+CGsVM1mhPD497HO8ZJsvaE3ke7cA36irI62b6z
2UF0whQyChlFEfmFW4SjgfD42bP+8SdMvIWX/3spw56YrrHi8/W08aw3OpYE/OSh
I5Bx6kwbxbBamSxymYuvOjF+sgFKY4ifKCOqgywBY7VIbdOWdQ42yKC/m+m+A+E2
fBui/HgQnm7TNsSn90zpiEdz1e3lsEotuLdwuLQSf8KOuRcSxqoFisHXQABV4LNH
RANTtoyr/2nbaMWuGDKDWhZ/IXeiiW3OvyDCWHday/tNzU52K3Scv2CcVWlYT/3z
3DCe9JBNkzumrI7lEYMweSRwlh0gnNl41qpuKShX3at3lvltKxCJ3YnqpohvkBRJ
bsEpjfWW5LgfUyuI0l0zxjn+e29zVIY7Go7hFXIDf+u+Oz52iE8kGNh+hiAfSK0d
CyGsX1dxAUDlM+hvWYGroziqDvMCE2DB5TEmG6o/6qDSk1TUctv2BEL077KGQBRF
QGUGSP6G6aomAzPb0YfzqkpX29qv1+Xz6yxVcDlirkF6FvU8tJaiGEflPB4sgg2I
62foziaQMzxWwAkytnlM7NP+mO0V3ySS660M777gRhdx89bc0UpeermHZJ29kDXF
Z98wXKNIEt8rh5d5xCcoqBiKO5lBx4WUOV/7/UjDTLlbU1Yo3Cqoa3Ja8EMb1RUq
Bh3L8lO2r6f/v7pObNtYtjJ0qE0GAjr29xW87tle1HzA/3jSLSBaNMqfL9eI52py
rvDQDhzhH5y3kOqRG/N6H5ISImX/mxrxrKFrjjYSCguFU0q2bOCopWQdsjO9Qjur
2SDj+xHjj7sIeTJvHYtSnokiee+WIb+pSr8xW6RfMiiZ/EbE21eRqKYkj648G2mV
bcDkkwNYEm4Awe8trWuRpvcy/dMZpx3fXdNiDceqlzk68ZHsfv+ekQs0tzWbfTZM
IfoTBiBgkENpQTBnuPCUKDYNUcWuHKwYSgP/su2Yjzo83qEWT0iZTSNrl/GZ4Ziq
C4xseD+vBWiu+JNQnKN97sdch8tJQztL8xydTUpR5R7o8rBfFmeD3jaaVs+6mlTS
MMFaoBSOpM5kmyBdw5CZqB1ZE94pY2kpcYiPYBWd71sp8bike7pbRHuVoFxZXG+2
Xew5xICsjKdXzu5Hxsp7xwdjaVtu02lv2/jzuSWR69SVm3KYxpZN+G70TWMCsl83
uxNMhFehYD2oAIqzJErk47S3jcvdaGK7TjhO6PYY3hQQHh1kbbpSnN7XtehyA5Sb
gtbdrr6koWZaQRS2Dely00dOEF1j+Q1a+Zrp8KNYKZPSEFZxZ54CSK6JBmM8J7z8
a+qvC/1k19w4U6oj0bKsGBORRL0Rivk4EdyjC7GVMxO3blu0BJHH3QZ+8IcfiuSl
cys/p2cB4cA9qgsVD8ZQ9du4ftx8z5Okzk6UNrZT8NdZfhwdBpLD/LFSKdbhdkxd
lMX/DT1C4AWMsKh2La81HgaPkLKGu33bd0x5nvKeVzxOLLNnuY3S/N+ldX32Phgi
w/Yc2Cdou3iNR0IOD62KLijiXNmdV+vc3zXGfMB8pXWKeJ5zGHfqVZF4K8zkURCL
RTPT2LzxROQuSCswkigidytW2WYJm7YK/HFOv3t6J9WTUg5hCWN5i0sgAZSIWQ7S
Y/r3NqcpOfTqLNMy1x9cWuc3z7QuLkkuOEhN8XhnM/pAtAanpwtFo6FSjlde9LwB
XplmHmMWjHvpglAvpzoHnIBStlNyoQxOK0fqKtIu1xAoAReMtH/SN6e9kUgFrWw2
dIYUG7RZh4XEtUUs1jaMOn3+aNHJh/AtdgPf9FzaQhVkPC4dOkGqhKpTxzYLOpSl
f1Ys//LZV/GZjLeXzwmYTfCQG3uHTgIpNTQQ9aNd33F26VwwM3OA4WBZW6XzasM1
NgoCyLBb1rx0eg7UX2C8E19bzx7DHzWSRKSjdab8Mf8IMyMVW5rxvE8BDxeUZkmp
sUw3nxN0GvzOtMCxlMYsqtH60axtGcjygzJSNnir0pv4YPeiYP4zdVI6o8NT6S7p
xsWaoqua0AN6UntCuq/Yd7UeyOKL48mY9pSv2Y7Eem1bRlVl2MgZwk4yDWx0TQaA
iAWKnmVD5DuqnmcfzWHLYlz1CzarwwcwGHxDQsUDwb+n/gihWiDmxgkFg/CiJpLg
Nid1uMIOU+pF9b0xMY4BFbaMBIY6IiBfs1G5p8yCH09p9i5RhB+1luBEUKeKacFN
KTJb//QoHleLadX1Fuq2BGLSSEoaqT3ZVS0btcwf08hXYlFQ4/1w+SmrPbxUSlVu
viYXeBfTdsIXQoFR37TFFxnZJFUTFtfI1JSUL82XXMb1wR4JPeLjU3OoELX514zV
LRez6vzHZudJxyf2dmqtLZJvGWqdBebgCEPQ5Zv2WQk2+8Bgwxf966OGc+GASO0x
aGUdsTOE3ENNk6gJrO6nBHjrOIsG95Fe3bDQmr+r8wivUOuoucG4Gmx//5hSyInA
vy1WZ7mvl60c7oKOGJenwNbQ3z9dKAQhzjEj3/gDuuKiKP/N2h+AzLsUUm4PZi6d
Zc04te7FmOUdp3YbBodtlWBDw59AuQ8kroVY5ktLZ4QBC4TmiNNkF97SmQ9wG2Au
JgXmaV1qUKftLo+js3aI/Mf1CfA1s9uTIOIY9uUTn7QkLUxEZPOYHogrHmONXKaT
zinUcX4DOk3ek0JgR5p6U6uXmxKSzqbhmFiWEuErd9nDlQxo7bnq1QdLx7O4by5B
JJgghx0waDEWize+u3tf7DxJ8y2xc5ukfkteZJm8PtpovAcRFyYHRD9iQ7jRIfXA
mBNeW8KLk1Mcp/Aluyhg8OrDuY9jTbAvZipxLAFSkWRnNYPdK2g55AJm/GFz4Boz
sKx/1xreBVbqXeRFGl7ZrST18pdo9kwDeqTVl5m1myrFbkytXgwmwJ7RsaFoG4uw
7whXZuy0ODuR9OQZrOFtb/eBCUJLFI+MwbO558ibEkekqwEwejrG5752OlKQye49
igdaSyi6VwBwNiaTHYdNOFg11nJYxWMtN0qzXVyjpQ49cK2tZeKiBGosQylicpXo
FPKCws1uJNUBktpmLmwCa45oPJNn0b4fBXk6TagkFC6qt6eNnj7oiA+8HvLcxfQP
LuZHNfI29Bx2cikILTxEpv+YqknG5dV5pLyQdDXtzR1OKnVpAWrq5XpbNJfO5a1W
jlmgCSueMTQ8PM1NLQaN8ROjNTRneWzCybk4bIqI6/fGaF52pcV8moLxRk3yvna1
mD52lw156h7lyUVCXZSsOkPKVrG5f3RqlPR1hBlZ3HLQfLHJRRvsyCAWeEcUhGDj
Yz9e2KxAANuztzYERoptW8K1Adhd0vJMJUVO9OsnczdZnx4tUNl4HirPwz77XPA1
zP58y0aIMBjA6HSWikUCXDtPM5kMmlI0Hoy9eDl1ugG85bbTfRfhb56O9mOSOCEm
jXB0KnjQuo/9dd50mOsIthYMOzfu3YOsyRq0lE+AcdLxp0H/txYf01RDNR1i5GKo
qWFhoxiO8mJvk/yf8ssLMPRQbYNgd6tzpJp7aMOooq6OMoYHWlqtAcNZhN+E7GFa
VIaU6qM3GxW4zGy+bFaPwBZTlWcY5P1JiAlw/8dglV942bgyK97ukGd+JFaTF5Gg
AEKle9DsVzyhF8eHFZMnawRAaJNbchRwbd57+MUY7U6rhAEUKUiBSJDmrxgAXIl9
uGN4VNn/3wOFOj7oSz0p0BQhGoCuQTox1fVXuPB6F+xGRlfNSpcPVvQLZFRdpqOC
rxsEw7460Ep9vQKh4P5t1v4T09cYkWeMU0RfhlKTRslwJiUxJ0mwf6s6Z0nFjlLO
N56U74IejyvUZhFUGb512XnpG+BAj52pqSp2MrwAeVAdkw8VlMVqzdYLcwOR++sG
xaHP3YTp4hQ0xi6PvYj4qNGAqjfxU6avNOwfaUgMiZayv1cqerbSbDeIxNpfVzuK
g/HoXKsbgxYhvBcv5RouePvyW6+EXt12zGt7yH6fgqor9iZQX4qNTIlKFnDyLsWs
P0l/0jgFk0HFf1KaSuJ23wz/utgSo97V8jddJO2KJoSrfcJVpjEWcMlQK9Dql9lZ
dKtlZGWMVC3k7o5NGWNo+y0T2BuPEVizvImAcLzJ0fATDG8b2tPBCJ40w5PGPQnw
0alS0j+6WCnv5AmiqTo8IvSXOokgUwjoC3WVAKMroZX9t+l1gAqd9dScxKt/GzeK
TfWGKlVqHcbwC+VzJimCwQ/W3avk+RDBPKr1CxdQnU+EDzlRIYN3led8mO71eGR1
MjMvcl95RA0DhIJVhJbyjNt6suZhY7aVDgyeGOaSdDGMP9iSVz0ZLsChfLQY5U+R
6qgcYDz8VKdJcoJnqaZ1v2qGNln2347JxcghZaNejtO8zc569aJuN60K2i9kSy63
GBQR94iG+g8aiBziK4IqOSXiQsu8GrkrBAByqyjkLHQh8Pho2GrmXdyAxsXlbCK7
1HlG25Y1/2KHn+jNVZgMiQ+s7DodJ4BmM36+7uExf025qUxhlnnlF3kKqPrfkWLr
oF/2hH396lvdf7AxU7T5BfHOYJ7o7xMre+i2f0Bc+fnEo2yaDXwqlNu7tJeuHfjH
dGYLJv9IrtlH08sJwKizLymX+ZoIikNR76iNRFaIZ3SzBmccb2EU3Njgwf6Q/4vT
IfFAjragN5rTPwF/BHDTjShg518JHq4MhWxmTs1HMFvJ43yYQ+x40Nmzm7noWxwY
90IcjLcJm6bn2QjBtV6D7BsL2t0YkZiS5gbG+aYG0xm9oXht6zZz/nC+d4BC3KVU
F/U4xbZ3GwwkOR9KKlSSWOc+j6T0PpCyB/KOB2tdhOoe8EKu03BttIXSE7+maN/I
9fdvnqcynD3fCGaAIsjk26J/Ua3G7T87zDm20RY+/7a6whor8ZvfA+zgQ6xbhO6t
zCoquYkNkScsLCi8agNOeO+v9whPTPjlV5CWLirqLffzg6PBFoYDSaXAs9O+XRah
2mCXoiemMcfZGJcs+CL3rc0LOJdCCdyWYPJ5e0dPVec7+RudQo+Kt1cSps8/Gj4f
C3oJD7wxiUzbM9KdDDJsEyb4n/LcmI2Ivoy+n6BY45kXPlVCCpQbnjcMgrPNp3lg
T9CyXzgxulY+9Y9yOPY/vgwI5NKe4d4orlB0riWKC/4zbF5l5GvEUZGaauaNATRs
c0Yp4ueA3lNjvjYOtRq0V5KVB7bJJmV2T0EkUXIINBK+CQrST8SPhoH4Cm4p+Cf7
ikHe9zVq/4lNIte9BNVg2eQ2+5Sww6alFMOtYO9PWFN2la29EYja1hrHukfW4XkQ
0yseO8Qhn0gLg2FY1QHfRt0658SBI/4Ir2zNXAaYrwnKhU0X7czyzxBQLYuu5DPi
INrCE1kH48cUKiaE+gXXt16rqPaPWHvnIkTbRTCujKqc968oTQRlV+cTUC0s2N4t
T6OccSSqFrONCG9wl2apFcRLeMWvU4UnTsS+caWKUq5+wamQraQtCnlIOMX1WemD
FXCWErCgjo1y3Oy6ZKj0t1KyHvLY5911EsmH7mXmOHqapm5qXlKGAyhoZlEf3+r6
K9lAkKIySHnBshQwf9QGc9s23wV2VJ8mmsYpqy/3MT84ohwwnltPjvPzL3b9YYso
QB+wggpNHdcFEkjp7SmOQ9p5WCkARQ6eJneQY6EY6toYgOkbhftC8dfCnaN5mFOf
g/9v75NZKunryq2nnCjVWEW/TuF1ukfCluRMxDYlVE5Bd6EReQzEgwIVbQFh+b5S
Yw+/X1WGLWPe/yhnwELwMTyETm2yhHOzsPe8Lml8k0E8QQvHHXE0DgMDiz5XuoA5
t4pNTFin8lgv6HUmb7xwUPzCbUxZWsqDh9DuJMM/u+bxA+XVvXMW0rFTEXVPHDqR
BQbC3jDB7rGX72x+N5xp/yfTiKE3zxY9nCswaRjB38i9TcjN4zRp4l3xsTnkx2BY
m7WY+63SKpxULonCoEPW1wcRPau7ErvxkG8UiZnEggl8jImUC9vX/8EuvHhaxb32
ch5jiycEl/Rpp2GrarxE8G/C3dOWfn8kBgjxIrCL5eeyi/vpaGPB+Hx7jaUZqgVw
lrSe1yUHV08112SD/3Gcokrh+WXRaKBXa3ZVaxPovhJ0hWCYWyXDUtisQIpvvAMO
WqQVrUi8rIbjlap+Wr6oqWCQpu+mqubyzkxD0dtx2Mqll/AEv0lN3+8Y60ooZilN
QMcbUxv6JEOyVlAyLR8Luo20/KE+P4Fl0ujS4GMHW/HCV1OnwqeByEdtgnBlWYBM
k6+CFyI6WMsOP1TOdLw0vLgYHQsvKvmcpiYuar/8TSnqOOQ/IzDHRQAaKWMXrmLQ
dhjE0tyDRPT2ZuZc8vod06gxquGBftgeD/aiMMo/5P1lGxXxTShCkSoodfyG7MIz
xIIyF2JLNu7dh9EzQPBUOSaHkhtfR1rxRlPxUB6vMr4+rkgjcHLlo+Z3MLNQYzYG
pmpxrifrhoyhMR/oCwA4W8Hax7dO/r0OoMtjWDmkwLotQd3FOHxWEhhp6q+3djB4
jkmBqfUOUgRcMM3Fr8xH+UHJ1mfP0vfv2XbeEy+TJ1TUgs7KS1rdkXvp+pxT0A5f
jShuDFyIFYT53a9wAOliD6J1JrT50KEqHlXxIEPr9U78A4Mqvc6gCJO5K+sHT7ev
mEST0rJSa/omkd0Kn2L4CLXnIsPlP8OXmUDGZ3vN9gqfM8uUBzYJJEEGSz5bsU9c
neUZNiE7filJka2q0v0U8ayiiatypQWudP0WOZhVslbE9zbeyyZA9Cm1yym5DkSj
NePNx97qwozOMHD1wLsK9Yab1aEl2RglwJIZ14iO7cuXtEnYv5CroZhBVmS9hUfA
E2BQvGouAIJNx3oFANmMHC47uqUebxUvDx1aPZWvmwmFcHHmghcFJ9wIfIvECO7t
ce2Q+6qHW0C/KaGPdJU+6E/D3ln3cpf3YsCzdPj7hKGRbtClXMWrRdIFmfCDbium
fKj88FGJ9LLDTIQ+vwDnysFbJXSVukprVEe3mxwXAlL1Sc9w3N3BNliZsISf2wDy
TGP3F0vw+OQhiJIuE4W1GL03FoB+bj0JnvM3V93OSTJ/xYeSgUGNI9O7DHo8rp73
gIS/d33bS/4o/Ty0YsuJuMnotlB9SZBqTHnarQZV/TL9sGchrWmQm5ktK0b5rqa3
sgAz+m9TS/9/1k/xXuxLBcwXGN8ohbo9dAC0dp+kggTcWTu76/aKwH37jJdOFZfu
T3NsFb+P43XdPMUWRVzqcqpByWHEn4szhuUFBFCsO98vTQ+wNvAXXTYPjsxz+GVH
iUNPtYKlVlAYhiJO+HWu4O7d2inLC2H0E6iuqY7oKMjgyh4BikXbxZhaw/2ashdW
+inOpnVWtuV3bLu5RAk28zGZW7i0xQQyynogtIYIe/jJVYZY2rVVm4REWaG6G9T3
fBGgT+27RqeDtOdYRmFZWvakJpydw68+tnbOdtbHrjfOeedpFlnYMjvlSDeUG1FB
g7hvRu48xGjQ9immP+7v11q6Lxgi7Bn9lAtIFBBjucSDd6Q0BAsOH6zeZexuaspH
cIESSYpeHU7u8VF0RpzDTtNgcbFH8DqMkhJLkbSnyD5160c6gqMc70qAVWjIhqwW
9eqFEVTH2CIX70ciK4Wog2TBxD3yFffMQft89XR60p3MA1MJEXwkWDTqDmeEhv07
Hf0+4X1Be+Hw8YsWqwIHZ3r9p+JkLg4xdSJuPEHfCa6Yfdp373sE06sxhD81oy9c
l8qKlvWX0YzAXJ4suuHmIDWfcpY4vl9/0uNew5xmTJvL1ybpa/qygRdrrc+nyVDz
XG/wn/7M/qucwPib9O9zITKybTjkVEw0S0lhWHakmypohDOjIz0kVN6tGqQP6fKi
EFkPWWLXxPhztwAexYT0mZi91MnkQE5nBEFSKPPWz1MsanRMPb/CdW0cxVBQ46Hc
ATlZgmTraDYmlKZ/jcgKz+to1fVL8mDmkShA5FEd+mx8h4M6nRwnndMpMBasN/Lt
+sQxomGn3hE9qVDhlj+1kRwafmbZFDXOLLb0ieoCpOIhAUmxwy2DGuLEjR0dUzpX
mdhyTLyfLoXXVDCdI2zoAayyDhO5hyF/o3puxa3mYWi5B/KYCZ1mTZocThuc4jwG
2zZXPCoj5iyyojgL+/gDn78yJSmzRtDu+Fq7GOGyMlaY4178C4umCs7q42LybYTl
SDUuP2fA2aihpkn6VeP0HNcO5HNkIKcBp67xtH9jAGPk++znOSpO+IzkCPSaz+Nw
2MD8q7CSzF8L8S7OAHn1rIfMhmvS9CzQsVUSP/KYGG8z2tJQcKUCJkESp3m09DSU
uZbCnu+R0MKdwvA6b5FetFrkN7TMw0vH6yjAmsmq+ni2O98y9/M02ixb+g1kRgOH
VuA5hQaOVPhFbNEj8umjEIPtm94iNclpiVQwTSaabsIgk0BnroV/OqQsldK0WhOm
lRpP9m+NLqIddIbPBp5Ll/JOgeRPRSCgGFTjkMj551fVI0Jg5UBIdQ3pLVzYkv4B
9f7XnHrffXOcu6+TrAQ//wNsP2il62/zMfItgbs4R9m4om8RDhkQII7sIFgBdPdi
ruI1MI0ojfGvstWQ0fVw1bird0EYOLwPg1TWrGcSwCzzVGXyMdZiwWPL58CjXGpG
N/5Ht5YC0YZahstr+yTY59ohQB8xIcSk1dvezoXSZzW2yqRaltXQV6hmIUhG4nLq
iPyTunX73AC7+XxpJrvHUc2bJfddPeOpOfi052eoOHAmtnYGbf5AsykI2A7xT4kQ
V0WRDY+AHi/uSmK7Ma4yn2nRnRuQPZM1xp+cG9+UtwCpQX34WIhOxiFMvG5Xlpeh
X3lA72I8xJ1/pJRFH2xtvIsIijxnM52CYYhoP3sN73DEIWPWEpIbk+gShhfTsSsV
6X2bMi2cZD1c8airtYkhxsbLmE+xGnptYi+d8MLB27bFnmTh2VtnP89ZfhIEZlZq
E0CyYmBF9NXJRzZ6Dt/ZjZvu/gpTaBIUzv0/R5kYlLdPKIzThXFOffeDXFDuUiGA
DV8Gg0PMXLePXJ+o/BLq85Ga/m9F1kniWgYbOiIcEORqaKaFRvgnOPqUBKFD6PHF
yVUHLKGKW+Aj6YQKx5NV3PBs+A/Ymy73JtbtKcO2ml2o/xMSA7VUEN1H6RiIIGVu
NrjwUx0+lrkUz763/l+xj919e97Qt/owuvsuKKbNIiyUGR9iNIHs+L6naliba5xz
d7ui8OFy1NRzaBQxKBBpkriFYdYS2xlejA3wYn+QXGKXzW4qoohWoEfvzRR9vNbV
FPbrEUcL+9wENi/+PzSxPNdWkHyMvsjwOT+iBmAb6pQ49A918wEEKh1/fzG+hB0t
hprDpLh1qG6SkwqWgo7d2E2kTzlXWdkomNt19N/6ooYLe18kqARSbjUXpZMHkcjN
pOhe5wldRSFChVTtbv8YMDyb7HcDblllIdKC9MNsqKUPzYk9FNDs2Dli9io8NUl1
PW9oQ7/aMog0erwinHbS6vh5oIGOa2QhJ10Ky1uNOHGJXTyxwGvOOy366CLnfyZZ
hHHSrSgVSFKutNbhCtUUkSX1UL9WZmLd4Wog9yKyYyrfGOVtb/SRLvr9DuzTXDCy
zKqPPlOxAko4IXjdAyoHSMQJXA2sse334z/pb9gvrQlDkLBA99uCIcWg2077Ofcn
eOXa39rIlw5nRPra2x9AljkgLD/CW/OeNJ6DLK7VJ930QSx59SjykXq54XIWDs+B
xi5vqhtTH807qjo7rrCz37z5+3EytMhqSYs8SukU44fpOD+yPMdT8BexEu1jZvSE
HyZpku9I6WNe+Guq5v/PRQRNoAH6A9skPpHdiHyD/ILssumSLRHCc3ZUPOLDcL1O
FY4YOHVLa4p9XgAYz0wC40ukM55xzFmAciQVlA7CLdeQc//vJ9WeOZXx+im4asop
Ad33aPa/SoIJLAkQCpseAcQdtrqod20gkqemtx8Xkea/UmE3mbEQ6uMzQdy6cdH6
a8SIf1jw13pSlcKGorjjadQs4TgncIhjHTR7mLCJvH1sIwS/H4NgQclP3KUMQXVD
N8q8z5qxmcnrYUg2NwRo+1yNiE4s5fIzzpKwCAUb/l6SB2/yu66QK8+3iKZ3MRGS
RASYFJYdZu4nzzYT/N2yLReff1BIfIiSXXyeKeL5+MPOpkRIF05WzYK4IonULGQZ
bOnL48yv1sStOOx58tQ9XD9X9tbe6r/4qPCeT58igfHSdEAuvNlxN1wQdmlBNrP1
9BuMnd6ypV4tX7q+8j61AILItvquEnphP01JkxC1VddGAgg+ramT4BjpmgZNEKH+
8DsbsuAxvLeaIhT7ykWrYEFUkmnAI+BQBt6P0gPmcpMP4towu8vSxA4wONf0xTSU
lRY95p52OZf9sx1u9xIbTQsSqei2bPh50kXJ/mxKtdvMOOizJd+ld+1eenBS3BN0
LyMldYVfRDMDpzum10Nqxu7Bnb/PWct607y28kuhNtiz/o9AhV24elnCKTlUl184
gJFVKW5H3NtWBdGRXbm+Ii7QCgyqnGkk4Yw3M1bkSbNv6onQmD7ZANKGn4XdCPCz
aZz+yCKSq9Wkqu8bmGcL8siNdGjjCW6Mr4cp2Ar6C8C1iT7wyXG6XylwBCe8Fd5D
IEjAcodnrvYGfPEp45djWoKx5CoBYS1u9JZSQYoa4fGYfp3YxSAw1rkKNwqhSaOD
piCM/gS69tpEKNt68T42g8ixnNL6mshNUB11mR7gx4Ys/k58qSxVCUYU8h4WpLrL
SXb4eACRuz7f4VTpOOsm0+sWp+7+PnYneAbg6Ah2qdNFHrSFXdNlzBqVE1VFJ4cP
EVYAJq2YZ35mMLlywh/yPitS4gpdrN+hjj1JMJI1/94FMhe5b5PtuA8I+Lg9zVkl
IqORm0oEx/4KTHRO+m8NNdpgkrbdVzwJDkigm58awyxDPqqUWtcqFGTe3s8qfTkT
91R3b5+Tw+AVaG3StNUUXmKD+9fz94KckehscM2w98vqgigFIRhYXUYjU0U5raO3
UgY0Z7mG+Uamr41rCdln8e8Qn3um2ai8NXBXGZnPHHFylus65ApWaTKdilMVq3v+
iYcpoKvn/WenFiu1t92kzT2locYK5JUkJqM625XXwwYIVv0kY7DRHwDH91JJ5Ud/
rHw40oncB55z40lOShE1i65u0LkQf768CSeLJNHcKYxs75/741dBRKaJLzO99CQy
nMy8F9JsrxNzlTAOaoDwZc5AMXgBWhdeKNzXbgmi4A8Wur0d0D18L9GIyf9TsUgV
+Gmy9802WYCzkIb4yLy5NJwK1+pJSFMLfw4jGMM0Gjz8KTLuQ2I9/Os1PiGnC/Bg
jKbS9Gryg3YhCv3BonUvkUgtpOWT+qKUzzkuBMBlAe/ueZCILHJQZjmlfSv8m5VN
2AHrZrgNdmdXjPuRB1U1xVD9UT+QFpq/z4UXuXuEpb2md16WN3hFeAUW4fUyWJsZ
CNudXe/yiTSOfM8wf5RMxRR+Iy69EKUQ5eRL/wARs2SMrP7g917/TwXXO1xxuIbc
WZjFdVPWIHzWvUGq55MzYM/g5n4PFPXZPaOvv13w/HGy4Y76K8UiUYQkOnv6oCuj
iDjXWfYNXstVxPMzwCD24hH/jtqfQnYwQiqJr2f6gxe3ifAWVoBkY9O29gtRS6V2
9o8t10GuPoaY9iRfQosflYqBnoXkN8Iq0Q2SimIzPMqudXU+CyffHe9XmrVlewlD
nU/xfYMxmoSk4z/PNUnYCU88SyV4L2L+IM6Fj1Jzw0CluA0FBwauovBLoBG3h0KM
k8xqjT/QmVBC4I6RRTrpZqsOivsXXPYguCIdfkGhBbMw95gFMsgfnK45lzPPq2vX
TJZ3tcifcJfpNqOYKoZDUgbfCt2hAzSghds9NSpt0NoKzTHqgm+0CyWqn9mTicsW
N3yP6nxp65Iy7wQUaPBtrttqw5ZCmmET0kRNJsV0Vspyy00KasUS+2aRhdA3SMq0
XMkzjyJwOLgV//IudkyertXD9TKngIdEgzE6ctQvjafzdvUaoaibVEqBTJYqIBFe
ybRy74K5H4J2h97FcE9qV5wILU6jp9UtsTWCBY5Cxp9k515dIsT3t+7BUt6rpa3H
vVZoHzqUnqu/7LqwqonSEviJBJb4qZBUFpB4yGs3mvPre7GwER6cSRxlPcQwgbZ5
m1i91X92+wr6yVHiqf81BfG16Zogz+NG/ImASnJoQr0Fe2LBjJBNePsdQIuVfEtr
uekuKWL442+H/f7VhFuDnrPrR4mK8XSnYjq+evRm5e8RieY0tT9+tc3upJadh5mp
4PWLT54jqs4dSYyzFj5E/k6Frgn6bXWeLlhvyd/lCNxF571BXZLzp66Dt1zGQKqo
PE1XCFoJljd8noD7xbNcS4aEchUeQWFYNz/00cBNrdXPQjDIhRUTXTWKT/aCkpj2
Rp3X5i9Hpb/UpAHS2tgeToV6/rk2bkOOm76ntyt/cTig08pzJTjIthaXb5KECwwg
1n0vFNtWnbXy6oO5Bwv1vIcbG2dU/MyDbzEpXWrHgkY90Ph0aD/S45tzSvj9xPJS
es9AAiS9OsJNKo8oQsSb5hozld3RNuUyGOLreC724CQjnGD6Sauysfye69geDgfb
CW4YDTBtoSTjDsTB9Q6OWIntJ26jgRjVLtuQhrB+XE/6CEK3PmH3nqNMC9Sk3gPO
E10Fc3ayzZjd+cUQWpt+GGd2FY1JwDu/3s70sTNzcDP+3J1wCZLLz8r2AyegTTRG
uALYWWTDrXkPmF7gNfpq6OsmOPaXqvYAxM20Y6fUOuEGtgrj4XYO45WJgVjT4ls+
AFZjw5REn/9ENe4bDN4a9PlqD/9GnXvG/PWwb8lRo2gyeW7VGQWR6rsLZVL6jkab
6aIETfeDT7AxwaTfh15qk0jykK/7GWsOsJ4DaJzT+XeyIc0LzOxSR7778t5qm+aI
YUtRGcUE5Vny/MeX8Q4lyc1uLUSYwQglbytE0noysqJRRT66q/y7cptB7QpGUmCp
m0bfbbshEIpVdbGVIZsY20Yk5/klrmMKCSi15XEFSCqhcOyjlSUCidReW0TqpvbI
rr+ta1egOU/je4P1TlJAOt5F6kJ6gpx9QdiBvY2YjBFOmo7nOcxEuA4bf8eN/KwB
3a5mZPBtYNjAKNS/N0nvepFFk8BmytwxEwaHUx03TlIbxwE4EeWgHJ3b0GbSRrRL
tthCAUC72boIt9cFvWkiFSVMwhytvoo9QSon5BwkYHjqceQxQJyRJpZvAfRLNEUj
tV2GTH5RUIC326Hkvibl9eJfSiAjHQkUNjX8K8PBp0jcPIZIa7yv/zuW94EIBt9y
zMhu5CPIVBsB/QMIi+o+T+//ViCjggRytvLrpaIHbPUOrDS0zciZT/On7ThqFL52
GBfv4lfB76/AX1z3e//pqJpPMulmzoMKB+SAmwwov9+cLbo0PoZJ1vFCZvpmmY/+
IjhtOWz0bZuNfebEz7p+sjhzttyeNpGl3NZY9QCArKSvccdNkEBN1uWBPtVK0H26
9QyVChRuTHGOwVfpyK8tAlKXA3PZNdAPcEkp2pKnpvykXZLAQkWEK9Y+6cdA+6z1
Uofp6YhqEbuUA6GcILPQxAyUWmZZwPDeGfYbUaCtbanPjS3o8/okdScvQ7nljmGT
WByADJdG4krcSaXocRqR6IVuEnqQNssCPDX9n+8AbgvDNCEtIgvrKsZQOv7is6GH
k846CoFohHejD5DL+dPg4nykHpfWVEceFPk9K/rVfOUvZ0huznfu3sQQL/MwhjNf
ds4L8i8SqwnCIk1w2BXWotEbcxfn0CKm4LmicXQfSNlh/s/5FURlRuYIiHXgvIat
M1wGTSErtm6HI5XZ4TS55Xqv5hqSW9NzaiYxENAcLYwHuP1KrX4S8LZyaeAxJhKn
+iLqMS9+r/osT62u9rQIzU8MsF9yb7IhgECGEV5wDFrRV2oUmKjy6YnlSQfFIBeM
bLfgGQRrPt/GxRBgM2AF00+AzCq8jePkwm4rcGmyci3QJrwP78Wra1o6W7agrxst
WGrX1AhqAuKqzO48IfQb4ZOtzexkroEEdGcBAHO8Bpc6xZKSr5svq9c3CoicO8u6
kVwXUgw7coPp7Y5/DMkSAfOUnnsfKSlhQY/ma8O7AeuNiQsgxC+n7P/zIpcjQu27
hW3OGP0rBh7aY+imoGTobl3p6e4wzfBU7UqGp+b9ftnJscfcHWKcQF8K/dVzePV8
ScGV8UAgDeJZgNBMvKIVlezs8IoNBXJxVkdtalbFMwPskqbczcqVthp+qWkoGY6W
XsBy8HlZCQzjbjWnbPEbRCftSKN9SqwhJPRQgiMImXyHOCuwFrFPJ8VPKijfNdqB
ysNWef80TGhOMAWn7CPhpKDfWm53TQ7Yt+WGzliuIQ1srAB0qJ3eTwlVx71A6oxE
MaCERKeDJ7KvydRPonijVf92VOlCKjCG30nl2PEG7NEBDp+ySvzohD+j3b4aAvhx
rfzAmjog+ptMIAcv4GnrZJpIWA2k7bIhQLy8I/LOKRwbx384xUvLbzpfqOGUfU9P
dIpFyEbQkULGgy4PbmOHERnxLhpp5iDq/WsCr5dqbxfeYvP0FQsTkAdFhFWjJvA0
k5qdp/+dmVdVcB9jkkMfBUgnBu6Vp5otV0v3UQ0XfdbMwCDE/Un2UDOCayZKRGfJ
8unwjHMao9oK0wI7wGVHh+a+w8YYQFee42xHVutsBBcReDhwHz9w1xd1evDLDziX
Z3hqwVp7lVV2q0diY9PaF7jsMKVFx8G+pP2L8bQUyvMN4E8E2QPeiLieXi6cKzNr
t9xSTBuItPjVocQxwriOd4W0Z7LlyHBfCmEXmH7WVMiyoogbta4nKWqcMfgQhzlO
ez6TlKIqcAUdfApRhRR0UjqCNMS0O9VXOazhnGtEzR93u3FD75ftWyIUtzycdhoE
IlnHsw1zXvNJsNRm6jEvdEsylgHGtVVUKtfi5E/1M3jMV2jIxfwSCY0tX/uux7/L
+sVSI87vzpy6ltr/H/0wO1veEqqPWK1DOmH8cUFq5QKv5qiut0oP+LCrPaQlVSj7
gj5Ukj86VpPviYMx+T6DW4DO11nQIcCRjy1Mq5kO5C9xDfH+SiNFeJK5CHbRnb4U
cRVUnFxy8Q5X2qO7sUxs5UQ3UHOqYDC2HY7KZV272lMndFPOIyN6aOlf4M5708LL
CVuIFJVbRwtEmse64A/EZw4CDeqyxsq0xmTA8uTAkLqUpuNVw1e++YZsCNJGlFFn
NZe+eHDstu3q+ELJsqKZbni7nWOSb/Mns7ftONYR81yJEPZJ4X2L6KGc4HElVhb9
B9SxiyJZjbegkdvoLooTEODiX5SZj35Ysg56qQr5rViBq+Vn72sRtTKfio3MIj5o
7SeADwZmlP/nESDg6GRWFuF6Z6lfFR8tNXAKqjyqZqrKxiXf7xNjG/WDPGUieCOC
UhvUapEtjmHMtJCwVcLIF1kmz5Dbk5GVq56s9BJl664lH214VmpXy4zHG9zLU33w
G43C20+0jAEpNGE2zG2//8ovhHa+8ANBoi1b7xx/7pw6mhuFbqFg23qyn3eclNmf
4dj5u+z/SrWa79pG3FLL8inGcY9ycDZ8I4uhSM1g1SVU0UNpab1rKyN30Ji4IXTS
Wfz43anPV/R2oIuXDuufJUoiKDl1zrETP5dLDnisq/vimi2e+CmLv33/lAxMczI0
sI6856dWZwjckjOLeTROJxDZBBUYSzwdL5xhxiEE87Vx7S220VHm4XHHPViKjijd
jdMnGJWHIOu8sq1eEt611kTcTuPLBtAXumywVSVuRpS7Jofbxft84Mh4VXJh3WPN
++xz2iMEboXizlptpqj+/rRwFxiTTc1FU0NjjHKVj3i2+sBoVLZ/tLizuCEvGYYi
McmcTQGnmNiecN5hKryvEm29dQ81LKB9FCsopqqACI0FCBTf4evgzz/FrabE79N9
ncAhIxMzST6hxCw+4J80fSxS6KdVpQ1FLU5HwFSKO3CMnEUTxvcku+unL6C3nXkP
zvK+04mKbL1yFoIBMYYz9dMyfAGkbqPO793f82A09tANH93HwupCcgMoEFLYW5KS
sKhxfxDCiLjwKfKF1gWkm+X34WiVoNYOTe6S4EePYY7KiSItTCDJnqqtRoumopKO
SBkXkyvm0lK3c3zR5gTMFGpBe4zUfJGJIwKi1lLEBEXKtjWQ3ZK/6ZFHcYbaBGeT
PwNYmpbMflQByNeMNKYAz9dkkUtQedK+hgDqDrcnupHneQzIsjlIPpO9PI8InrGz
9nbnIFRQMCPn2CEgHGqct/TXlJ/NlkjIibZVHVOkSKHVABXaHL2t/guH6exGEoHx
S9qan4Z5ZtMVh6GuKc1VIHY7HGzcEP7HeBTvtM9T3OkYJcQmxKbWnfRH9ak8nDER
YtZo3lIA1VcJGaxc1rLRR7xUnjGr8R9U6bdD+ynLhz9EVWXLBga51hYkOuVAm/e/
gUo3QidrEypLjdeYY6BKBxmxc7sapNqCA8JoyMO4QQr0X+H3l9SAYMbcvFlWr1p8
v9N9sv6VBTQezYov0VqHm96BiPmjVNryN5riwzWMNPRZX7/oOrj1PnYG/yQoZg2j
vSkSUd9dHyoTWcO1T6PoPRKFOImzqSxdx77CrQBrmm3DW+HFgrttQcAIdwfAsmVp
aErGSrztuDU699m5d/1aGPcVBfRAtVEc7og0WGeDyN3wE5/VVp/C0Udee+K1XDzn
m0siMmGnPj5IwxziIOyWq5qpp0tQvoIAQjQzY/c+JBTA4TMr8wjQELbQAJAF3y1i
/vC4JDW6QBrB8ud4mMUI2secktAChQNk+yHdMx7mOnhE3Y4A8yGuN0ASpYs51hmr
4g2sqWhnV+44H+FQR9suvbqIv50Bqth1bTIrlTFJn9lYY8/hyE5SXeI6uTScUxos
lBz+BBjrgRGq2m0az4ixtfyMRuMhpuM5m2bEAB9UFz76ql7bGaetlk/TOHBn+qsZ
gCSI2e5Kx/06lXQ3Ox47PzPiX4tDnLoLdkJWv3HYOG0FALFsQXd/xrb6S/rZP1jQ
8jwVTixWSfWzDLVOJKyomxLiPkeXF4K4J9pzoakDANys6ZrWp7sc/GgTYIdkEp5s
ryK0+MgaITDkNBhgAz95ImCcqfgFWntZcdQJREU2AQNSAhWZp6O9FQUu/bB/dDis
YKQKV23yR7E1oKhRKnC1rH9b3pGXKwRT1hGFWuUdTX4V+oSHVMbXYKUR+fC5diAE
22X1uG4PdUboktqT+YmK2QjiHqCYjt38byF2NMliYtWH9ciWwfh0QAK2ae6wI7lG
B97gpxhw6bIkqi5lxB651SX5tF8LTfiQHXEuFWrTBPHOXm73IxWpEkL0VWybEi4H
eIoG6D+uQXfqLfIs1MW2BvjveV5Ge3J9gC1An/rnCUce85I+GNcwF+O+iHMQzf8k
APfkudWa2AtDX8fD3P+8fNfJhk0X5iOUqKkhjaqx395lGyLX03DOLI006Fde0BKE
GeLjGqSiSbNjQNAOvbtYgGQqdJznc998mqxl8hn/jky+SITYZ9wAFtP/ycGKmJUe
yLZs/Hm+aFwpVrzx/KxNwwJFzC2OD4PsemGZe3dTVw07EjmtOA25+DMzQJYqWOhc
3VskIrfLsG0o16AMJh6FHdQoiq98gTl1ayucllE/kD0RopLd5dt092dyeKN1sMaX
FcjxWfx/3tsfnGP8/HPC6koo/gFNndxAzOrySzrqh4CRfUSCufxGbTynaTZMl46j
D4l8KAwuD21QoETym2IsEmBCrN/MM7x/kO/KlZlWIwSoKE46wW7JbAYi2ACs6uzz
cgF/5gyZO5KBxfRMFNX7Y1gNpF/4EKqcFtEHXoU0FZDwOkEqLTaREyhqKCQFKL0A
c2dW0qD3laGI8nlkVD+JtzSmqJsSGTBzB70MJ6MSQasbYo8NKddwwUik0QxUxSMc
bfWyP3BPuHNFWBQK7cP4MkV4CdgcABg83tI0uvz+RkXDwIinaMkUgWGhEmaPAE6/
YIy6gJdOc2KtNjya1aCPUaUuMP/AjEkQMX81t+YSIu+qtQONiH1QEYlshdOOCRg7
Zele66yTMDzlzFO95ul3MSy3w03EQ9vQLibG6Vwb/+uGwiusqpjGFvJ6TT1iw8+P
jkez45yl/vT00N7bWoeNQd/YnQKAyYt1AWtBdR4D1B/CjGStjz2L3L2v3BCTyLA/
1xaHHp7RjwQMRK8d1qh3JfDHE2cxsO+LY2m2vlTB8RqJ3ffzNGyXtKcDw/w/VRMI
p8VMFJ29Aykh6GHUlIpjRyG5O0RGZNHM75NcJYWt5cLmsNuN6fwIqba7EEnLHWnu
MMJnOlsc7JaUohjdgR9GRhLFT2GzkUhQyjscCOY4noQRCqdO3A98dCRTw6DL/7xl
/uQv3iVi9BC1uYGVGDNUOlRFHUq4UW5S+6fpt8qXapRLwnhmoUGVBAl+8kYuAwlO
udRQj9P+ovF0eLPl/GE7JJpysUzzoYrqS4aauQobmv9Gx9Wc3QrvznCWd7c1grn1
8FWyVBUbD5tEPyWYwRJv3LKEWs6Mf7brB9sfKwtZuPHzrZIHAh4DlMFGI6RpHOmY
rW9HpvuDFoi6hVZmXONWed+un53kMhu8B370m0Fw9jP0yCaMCrfX4bGVqU5RpJ+D
h03EgRgjyoy9+i1wyuz4BLtcsiRCTAd9ry6Isr7yqW0CtQf1lQNbi2RJOHrI1ZVA
3fOVTSGFUXIcV/H6RiVjg9iOQETN6IEBgWkgq8zlvXpRGzNz1Je68aMzftTml8XS
t5nznqzpg/MtU5Mbn+iTp+ZNfISDzCHvBPaLSkgzHQ97oBIV8cwZJiuWYxW7NtXv
7hRAbPDYRFFgg3eDM4ivJYEciJD65UWMmttShf7okQ6sBTNrDqnljAizV59tc4Wf
9BLQQw7cUAiqJlWAkQU7kdIrEJ/1hLRq+mQgRDfU8lVu9pFtGvYgxyneTdbwhjQb
7qL4eeYOmNlFqYlQm7dyzRx7cRvnSMXQdL36mDoMkjtSzyERL3gT9dCCoLmk2TDz
VTGWxt/mZ2Dm8wUsW+N6Msfuq5sFPET0GjsSfnEo9R3PMuu0FSe1R1OGsicFMnkE
S55WHhnSsqsGc/LsfMCF0iO9rFJwEDqlyMdj8JY3Xo50RY4reZavjpCPJ2BuXs+e
z84+fdX8C2+BJTx8XBr4O6PN4NZFeDZa+/Vr3y2wm22+44Cgc55DQVJ9yMaMggUj
YIxuwJmiPSwW+hZfhk8qEURGhdr2aHO8DTov5nceSVMfvxDSTd7zu6nJ5uWCoS5q
4yUxnU5ypjjf7ejV4pdyWe1Y8md6OGAHnShhutcnFc1LsqvoIZ/bHpQogCvk1zyc
dN7nYGnsXfcNIYXx1n6gFIbs4cNpEtvEwDlQfXX9C+hjFBsZLa7EjFSOSUe+4kYO
joDhMcqXrGJN6C90Aqb2q5P1kUZM/kxS4tzUS+6s/u4pGlISuk9UbDdV5l5KSObH
dFmGm4j7Kt94824IyU/3GXyOPHyoFV91uKnNeosaeODOvrwaJ235A0ZoPNC9ZWft
tMA+ybNX2avbvRSwgA3j5TeA+onque2E273SJK85dwSlMqtM5M9XcMPB5hUi6p8s
fxl67lFcAioleFK4Jb3Zc0YuyfP+0/8zT8oRUVXZI8olB3ncsN/onSIMdG6yMH+H
+NxFTcsG82aDF9o9KfPin86kpGL/T5F+4Hlo8c+JI8MTJdPOaDCGt/QeyU9svdZ6
AMV17j5wUn+YQbybJepJi9ZgpldwoGey/Jb5UhLDLaiu3XDAa56/kGNUAO/OYtRX
z+hIHGwEJb9v39GYMlT7i/DJbleZAr3kD1AmUlbjPG2/150NgSYgaRV28RRwafb0
BKW7x0L57CjvQhSLavi/mEXxozwgvTLsYNXf3Urrhhe1Ak+ffxj7XYmMyt1fmWf+
xg5L8Qy8IAsVqdpn5JayUN9Isi075lFjHeIc4DEIpimtJV+gnEfV6GvEBuok4m+J
SFVtnGBTnlB2dATcOJz2r/K9wfgmMPDks4P4Z8Id4gMjK20LfrsJIWe8nZV8A2uC
gGywKt2qV7LSK9WzEpsgaTCrZI7p9dp+O2pscUGywzn9Sw/u/8JP4XsYxNV+zhmM
dNRXDa3PfmdOgmrsfLk2cULqeRZE7aKvmU5a8IUmWucdTzqHI48spuPhb3nvfp6C
psOyNUq1ildZPBAQ0voPaueoHfo53sMPt7PYgVGE0gmOCngQEhHZQzXo9TTQ9Ahb
kHkuh6G86ZJAETvyPuWxyow6uGCMX5p+GrvZBTL8zWtVKr7/k+j6Y3668zU3bZEU
Q5h/jtwHcsINZQFUoWhG1afEoFgrA9UhrGiXcks62ijaNHiK48IsU+lwv9bg0Xq8
saEE68HdDMUcP7NQbFFGkS7fgONKZi3p2aHTBvHZWgk4faaH+qTle+ya+H+qQPU0
PUzFbj/kvZulG+xBnKQFreb5nNbLTUAtOu3sSEXEgRnJVcNKy7dux47E6zfrTe3Q
3Yc4aGQgbP2Pmfp2lMdqszCTTu81VxnHoQFRVwC2F8hrNPIC9F3+YibnA/3mDsLB
5StfnKaB+iLPoBYAhYIZG8XdqYaDz7OmdtR30q5Ggxfk2t9VISXtxvaTf+5x7GtK
622Ois5CRtKpZVQI4RFrJzjHs9kZnAZ75cxhZoqDTQWXlTjGw+m0Hd2itrqIgO0p
+St5AHRK+r5UBbI6Fyxk1Dgqw6ZboVTdHdjJA+4soRGQ7+FODOTLDU8E7BZs5FZ0
VvPPh4+CkUEyF77jxzsdnqer/A5WRV8uWwLNHbXabdoMhK4nhbRn5+4zNN0NWvxb
ziizYUoyh3GcBG+Zd4GmfrEZ8/JvvUD89c0l/OhzIj+PxEr5IZT9Rvw+rRbD5sbv
xR0IL345FLcmt9d+CAeefYgJ0btGjPIg98L8enzctZVtDpfCPR2o4DXgoI9uDUGN
IkOVfYzWx7iu/gpCS1b12+fu4BTvZ9/RNd8zh1My3TJa8bqSeDqa7I74gIqI0vW8
NlV200Au08c11ouvcPyTgQAltpQJuScoKiRa2ZwMgCbiUahTFhyRgDOZqfRlEhV+
gEAPgeQQH2DHuXQi+kkan25TdxiyXnigROmmUDcHZAVg1HBaN0QTctqSK3a5tAxn
Hk501jA1KDM/bLt6H582nZLfQRz53oXW1sEZSV/MzvDr+qrRNMaa+za5a2r1vOJA
Stmz68kzSL4z5zGiL/ImQmt6LUotsTSzvhPE84bdda32QH7o1niSrEB0EUtXdBUt
3g2Zy4z108w5V5XRWvgygKfzlQgCksliBKti96r63P/MEbaUcPWo6Upz2A23jnhz
DLT525s/DbdhiJHmeDw1b+7NckspiYDg6P8xEgKVHlECXZMLSBRrz/hyRTYSL4c3
xDRDmp9FLKq5sBaLKw2v09lqSzGogau35w8lR5aQEIEWvThKsQRsSqC40PD94E0H
MNAjK5No5QsisiR+NcYT8xuB37leg+cswaKOIBDe5vLzzynn1hJzh5X97MlinQk1
WTcqHeQKUwzCZN7B/Y9HALs2Fbrz4G5ti8H4ZRIp1eaLJIHDmgm4sSYdss0yihaE
0wV52uTsj7v3I6jybz43OsXSmGwG3H05PZ4FmeW8/kDew+YMRXJ3u3UyQvTAHdkt
7nMpOyLTgCD42rzZWKJkPlSxWWWcKwb4jrsM2YpK9Nmc5UuVl4NAClb+Zj3kTbeo
fn7c2f4ASWqq+iBPdtrr8J0o33hpQfTaFCCNeTPWhn1FYyzakr94FIlg5ZLsE6UG
kGUKlRDq+T31TQzdpRWGAtz8QuDlf2ZBnGUj32kJKBPZIRprQ/NxugqSYMGdFKP4
aOHWAdI5xLJwohm6II/+JDXEnzwb2bcBfSWIlF1NrzE5ldFo5ha8R3IYJkGVc9WK
EmGDuwF5bOjgXJs1BtKbSJHyAu1ids84wUDU77C4VyisxRX+uTlAlUvs4a0LbZmC
KliJKB6MUA3OIjmvdAoTEW+KpY31e3HZGgdL8UYRpeodlixotCbPp/wwX4iJgggZ
48NcsK46mo67ZCSUSJrk+ZrlBrd+G3SLBW6M3y2VL8wEtkCdWJVBr9F1W3AdOaxk
xCSDatONj7F3jPuJ/P43ZUpthnf4dBuc+T/W1E9aw7JV5lLH/tO8t0SoKpmWr8Fa
tl8i3qW23Leo0WkRW1QYWAxX65plqy4g6RmwDHY3qVdmEdSz85PBLoEZ1zGSt7/8
UjpIx3q71VDtFRyWfulJnNcLOK3KpWs06LmygC43mTUzMnOPwks2rr4tFKAe7+uV
g4BQV18VySLaxTU9+m4dwBQQkKryjw/Y6G6yK36Hacxhm9wkenC1wzyO9t0nKhfu
hFHezeXJgzsjYQq4T9KWZkoworhH6jz4QVNbWEVZOOoJ9KyOUlttJDkyqCMqpNY6
GGx69FrrOKApwE0RrwdtMl1gltpA3zMiZ4sGszMWfp08I5cFSTNcrCLnHCwhUrND
XZXcRUYmH2qZInFs0vvyIdffnR0U2ZDID0/EwjpYXUn7aHPgbdTNbNg70m1GsiGz
C8rnb/2QIsI6yAIvfi9jledKi/FkSAQAEtA713rZOP9ipoIhj8KO4MRWbUKQPMY0
PyrXEq2PtJ+/jl1eIWXygHZPyHOIKDyM019Ywj7f26v1RZEtpytlnX76MVXJ4XIf
SqxQw49yxd0Q2PvPD9DkaG/0Ey5Z1Kp/JCHaPPbGfe+g6lnK8EUrkzPxIPqQ4XTh
g7n6Gdfs/tmjUnzSmXR5G2pI0jmwYWG9Fx7vKqSlBmnOrOcJL/LAxFVv3HC4yawW
zH7z808bvigL+bPoOqFz6RzY2yHHPGsdUHxCn95RlxB2uNQqQCHCcRUxI3j30Dni
VDGlOYeTpZ0WAJ9/olkmAdfZ71tE4xi+qcLz0cDBdjXBS3Zd923BNIaEtu8eLtPj
G45QpiTQHPpJXtqRSFJCSHxyzAv/czopqbHpBBVXYebdxv5zijsiJP+VKC6I4gq4
kh2pBTul/Cwk+iB0Upqz9oWYq8snO92Rnsaoz0QizqQmeTMk8IQS99vPvzWbkrya
K/2m8Fxy984gag9deTJGMZYnIsYcuROPP4B20o0sIiFWPn7k8y7fBMrlx+GcU3jt
54yJSevldgMVc6pmxA5a4cUsghWy0FuyO1CmTa9ultiYz4jrumYQ5gy7VjIqaduB
37KBeXjY9HixwDsk6G5bYKETG+a9un56oTCMKLMBvPFlNzuWsONJGzPF094/zclU
ky/5GJnicu6kblbVkvp0pTP66W1dBq/uTF0y1yJud1YdvoJ636r0UdjLl2OwNafy
DB44KmCcXW7BND4yslfhqRKv/pW2GHVtxEaaaIr5XSd6gjTjpq1TLkMPdGI4wQQk
SpSg1OZttLXe/QmaDqWfjVVjB6qSl/HjNUi+ydzRnuqYnqGzEhVQoDb0pmzyJTj/
I+X2AKm26drP0xOMla8yc+1lfgXGV9WahW4BnQPbjzn/1ivXSKpjAhH8f0TOZh6O
5NzCc8/203z5qYpmjjuZZQjVDdVC8FqOBTtjQt+DbImr/LVxVycdl2LoFiKEGKs9
hpHAB1K+aKGIyGbrOdCO4y+3GzL/H46Y8op+i4ODtCPeBDlhmUBbHDkx2FKdQAwg
IsSbAVlfJEgQL/nmdxNjivbrKKVYdCJ1b7QUqHbRMm4WnWLvOCMoJf3WgJNZ9I7R
EOmnLGOrNVqzY+u5tWFt3ugpYEK7tP0CPJ0efAnEnZRv8Tz6J10FfFdwBmF5feyU
TOCOrxexzMkQOsuyDJzCT/ryCL9p+8pZtwsPqC6y3uEyF3US5pJ/yITwIDkmpqeG
fyWuTeVjXz4btP14gIfu5RRQkMQZw9eCkMU9WxhP/Ms2OtK9dLJHV1/WyKhqL59L
NXkJk5kSGeiAUsvcF9OWnVuR2C8NRrZEkqbA3H0Yoo2QfWLtSsk6maJB8zaNciFh
WIxPU+EJSsJEcvZVHXH+NHh9PaBbSiFL/sBbyEcq/f+tcvC6bPJhx4c2LcnBrt83
5oYEppKQ5RRtFwlNkUg9SysplTRAHASYw+1sFKYGhxrDUzhcQA5pekmF1p9gf9GU
FbuYqzMbtWi8il8DC0XirUpK7DVNMy4DEfYFd/HspViDddPVTW2s+xEEExoE2wrY
ufSfCKpEgtL/HN82Dgm357woYTvBwBI847M9/9nN+WNUOn3quLb9OrxGzCtlXSw4
n4GDahM69UPBzfRw0G4+fqWZs00Y3ALa6rzVUGQDA2XOhbNtpDxNhLN8BdLAm9nN
sYFqn7WNEHbfXegFNP8rMsPEmBLgWz/tdYZjq+5gE+L1U9DzwtCIVNoODqQDBUTU
SuTVsutovDLjopF7kiCt5vz0tyBvohbLV0blL0r+C0NwelgI8ofhOZlSY7LBn/SL
dwCqeRU1kl0QjmMvsievBxs0A+HhE44JvbmWOJCMOlk4Tii5nPM6QZllibukgR/8
uYmUpaqQmOA3+z7QXHZhfB3WxI2lFvY9OZ8+Q6ojZgK4Bo28NIDw4dpEXLvqxiQV
IH2g0eMWZ/GImgnMmcDolSyYyC/BiVRE1ROBBhXRAB/uR3Wku98exaB/CeLDAJ4B
K4l8LYY/ZuiC+u/i04pGKm7+23QpvhWI2XcUPejkPYl7Y/2ecJimo5ZAVoqBDneG
4a1/+o+hTYK4Xa/Al74J0qVO1pu7gZ8XphPHZdSzUbDhMwKNSn6F3C12EWfcvgSC
HwoYbapPA7tInBybWgCxt/UcILb31R4Nmpxpx56eJ93yjXfO9txGyuc+KIjfl493
RX5gT4aPU99ZVkuaFJibcXVdJwtQbg5iXevV8ZYTV8imnkIH6CbZKFfZFM+y6f77
r3iuqbFda/z+LejmV/MMHIh0ayjCA3EI9Irb56DkVUAP6gRoQQNU9cy5gzXfP0qk
mHg+7jC2r8S7JFiv7A7Eh6jCifcbFJU6LstsGebXSVVYQu1MxWvAfnfeRWlsU5sl
51D73QN+iCw2DPn7RPXYT08R/YHdXjPmywsq6DLbHkvd99RP8DozYqclUfygbaq3
KbnRRViWxzgER3UxJwU9rtSYjfwjE97Yv2RCva+Hn4ynaYAI8ASwPoAra1CcDkEW
M5UFsEfNYaUK1Z7Aa44LxrWgduI0DNCy36aty5do7Lxi898eeGUyO3a5uOVtb0yV
xsZ3plag0tPl64kBMR071bmZLZHhLfUjmasrs3gJOVBAPXplz/2F79cF9Jo9nrDx
+zTWgZEgLISRXibQwrdCpMmmQE7ocomquFk3Pci2DxYhXRD2q26SFSBeI8EB4OVl
pf50/gedzf5hMNtcTumGi6J48wWE14XIMUhBNkpOXfq2nb7QbA8c7aX6QkAubNu0
fkW0pmTUPcuTaPbxYzpDHZkyqrZqUCx8aq1MUpghE+H+Aakt0rnlY+7gLBz4P6sq
dfOo/O701m920n6h6aDN8jWCVAxg1R3vFRJJ9a1WnYsrCPcSv+Zoks8mVPIH89Qz
k2lPK+fS32RkHSpdU3nr1/bteGKE5hMnzJgu+Hw+hkDrKQU0R1n0lVajrG2W3cyu
WfWuLrH/aVTXuERh+GluWUkME1EZcq1JOYXx9hyNkL1NOALrRmHQTl2PbP91tzlr
MF+MJ2OJZ6ixB0bA3eSoqxNqtUAksOttmD2JseaYZ6LnGbEhrIeKCTmzdqoSX/V9
au2LcPY0jOZ3IDAa2gR4q0Yk48QvTb1y2jUADxOp3n2i2Ada+Irj/XJeNPmXhE6Z
QNtuyQ/6h0OV2wMVEnp2HQMALZnOVDStWAbeA0h61aKSe+uT3jAWjMF9AMQjvXw2
wCai18SE17nGS/QrfS+e3CBV2875qjUvO8sptN31OQv0uxVuM5Ess++q2kf0QI6Z
g9jraB+yY1HRlbUPTODM++WyAXYrljfal7dZ7xDrdAyJdXMo/zADo/Hj3p7nz9kX
joSjJbirFD15cs2R2ocdrbrzaciaZcmqd3acbpfMlYdsfM5wMaoWl/AJLje8rOdX
QCg60yo/5aXejEGIAalsn4SyCx6/fBAekxlKrnnfSaj1VKucpsgTGhmBrEkRrB8X
CTIbbs2sr/Wj6tJ6btvLDc+JfK1QhF1ojyaSPKb72rHKrWDuNLH5ajuBSTiqnFxH
3BJtU/2M7YAAH563Td2VU30uoVAiQvcasQiz57JV7XgnR01BBZRvAEQBFPbkQS5b
pS7gdCZTq1BFFWvz1JYRuR6eMdFiD09//n9W7Vzu2fUSElg8GzFFqAVahT6IQv8M
/QEvdsDfH9GaVwR3aHpxrfW6ZsL3ABNK07eiif2kPRR2FGKOO2Uv7CCwJVSc5HEs
kX7k5mvecoNpMOEUmX5chjWZKZqqNAGwdX5ytTbv3MeE3w+kwbSq2fg2yWWIF13f
5BTNYUxaYdYtEx9OpI2RzT+F319rwn6zngByKOFmfzDvKcYs9HgOaSAKnjetCpAD
oBQQduZQOHyT5HEESNzYp1bvw5krxsKoNa8ncLoA934xsdD8sR7hnZl3gnt0gh/2
uQS8Pa3x7EslieLmlLN8W3mKsqsmhSUyBpzAILqURASg458cQKqtLmHCOqfsh6Xs
+kt/PZN5AsgIf5yb7l8S8S7bNSlz8NmIYTn1z3Dsr/dow8elS7l3svpRNJXtjwB0
Ni6yTMLAE1Ihl9Z3DqmwixkUU3ZkcGg5e4CD/xwPbXyvMzEBV9ZujuekzNkONAtN
hSMvM6389AwXdPDPfY8wVEyWZ+NpNID4qCX/VeWZHctMBQuJFC5RjJUxNriLjGJI
3kRP4q/6RuuSEq8pe7HW65ea6IM9UvIeiWH1GyTxR4O9rajor/05zukeYn4U8pOc
oKOZI7W+jFX6NER7IT2/5oGm6HxK+92zppDVURa0etokBGvHXgFLBJE4pU98hIdv
pE3WnVMnsSw70uC9OHesoRN1lx4Wic/yFgNm4PP6AHl3VYVk2RRn5Mn9NH8iEcnF
jTMCrJS1GqL50nOItJeBOBuN8z0ZXqbilILaH++7AGIBAkSgsVqYK3e2y4xFbMXC
SeCm3KfTkdyPa0QreRMrnEGxhpR9kvCWG/QLz5pP0neDQynacoSTViNuiRkmuDR8
xfFn5xtgZBYtIMAVefzXKr2MCkoEBaFazO1VyQnJG/mjmArTjtprV/i3f6X/2TL9
b28JjEijR9z1AwlbNAI6G5swXoMkebNNv+S94wUAL1dWnmLK2OXbCK3F7EDfd4Q9
54MTBjIJizDiE/7hU0XUDP0eI6z+Q6l/+dWsHzYVHw9Zjh8Ze8HvfwaBXxKGxH59
xVWbH/X+AJc3pmRSC7oBJ3pU6FKCnlq8PKl18KNJtfuC4x5JByjHDzgDsZaabIIL
P43ZFWV1aEaXI0Aj1w2brpa+e0APeEE/PWoML+URXJRGu+ul9Sd0MDd61HYTjNuL
dyZFBrPB/ZQlbhipp0HLyHilhdK/oyHd0LSo9+AX0Dhr2qVcGeoVUIuN/IXGsNLW
xjb1D+r4Tvbwl5l5XVfaaAxn0mao4T6kdOvzxc5/u8/EL95F1tDWAGP6CmOeXWvt
3htAYE80ORGQUzEJwIY4lGUfsF5k1uLoaB71bVZxn0EPj0XlNDaFOHoRBIDpCG/o
4wgvNckabRhQbqYyipX5WqlpJo8r8K2Qne83tfVHvr1V5MMig+t4G/2lWuJ/ZQRp
CRXQZ/DrtdaLFbB6AzbN2y5CkwhSj5li+XsAi5AMAW28fhjc4fOR9SJx2NjhtbC1
ksCYED3Y2WUr9nxsLl1c1dIHIVamrWm+Ek6HzfcrseFNhUoEugRqm6eq3cTcYbkP
Jwxvkt86ejNYfcTA0uaUTwswYCftlrxxvbduXUGnhwvWwa15pBCP/0fPyam2GOIp
lYHnuESkKmbazwt9Z78/2aG9I77WWvY4HFryoWeVX7BtGZ1i484rSki357RKOpVN
g3P/q+nP2+5LuntYKD81noU4Ubzbivvo/6PxN3je7037e+kB0ka228TD1g0mxmFN
gx3opyemLbDrtXh9P2nPD1jywo5wDfzBg+CwW+cFX6xkPBCYFZ0G85hrnXA3rvP+
dGC1jdH57K8haHBBw2gorPsLxWdEJtUVWeYPX/GAWL6+Ns5kCmqEJzBJNOEAS0aE
MK/gZf7hnDf36JDB0vlyDXB0Sar8W7NkEdjZgzObB/kboDIEbB9H1Do+KG3gOj/z
nBJmZ8nMUjpq8LVcXrqKmbi3s5n285Gss6jR/sY28Njspa/0lVFDZUrcCFvg3UWY
fGlLUVMGfiGySz98CFZABlaTV+ZDgN9DdVR2CP0ndB71wag+4kAp4VTN1l9gEJrw
I1el3AyTwoDClJRpK2PmQhGiRoInzHIRUtMwJkTN7rSVMYr9Rn9TZVpkhwDgKu1E
x6bECaFSxR6yYlVyeNFDdXmebtokjNMwVZAvQthmhQJ+SmFJLxAcX+usaMkVLgn/
94uljNRtjtN7AlGa2NGJqiQKafvMbBihJZBVt15ovWkRYXP2KLgYYA3llnmfHfvs
+OXC5urnMv23n+uzTGwqN8l8pbyhRklZN0QhjGBbqEHwkFGAACj2vLlBav0j4oaR
ixN9lJiCAnBo0a9Od+cXAyxwffCqz39ZWbxXXZSpAtd8P4El6Iy64m+ECnA2BlwF
ZVkxH5g9roGd6ctYtdx4PwYpJ8s7C8vWSAzaJuidw4VESAR5c76j+aotd5s3WZB/
Z6eBJKXnJ8e143zfjrrmyfwxOpvH6HtYH9ZMev3Shl6hY+hAZYO3Ei0GExVmrBIp
vcMFKvx4K1AmJx+nI3SuHoBLZRV6VXV2zbWTAtiVMiaADZReXdcrjo+qx76BUtKg
1ccL6ynLzGiafu54noYNtVAI9aoYSxsGnSayv76iyzeHQ7Q9B8iJkqnGzo9L8xxp
+tSJ8ELSwSOCteWAunswhQV/cq1ycGUKEWg/P6rS/7zzwWYgqhuRUT2t15QpL+ge
ICzSwAJAnqKt13sS9WXZ+y9l+gC+pwKZCSlsdfrsQaw/ljcu/dq9wCPBlD7GgC1h
YcvVqKPji1gh8zm0i1mGOu9VOvk18euYPGHM/Rs8l2u+A86H/gG5WnrmUa97UOh7
1n3aTqVmptEnFzk1SW0m+qhyWwHoSatKdsCS/hIZCEoz7AbJ7aKuc9P9QiA/dfdn
I+a9uUd+Lwi6zfXWzLvnPwtSlBIwLNt41JHedkMPCb8MAtzvfpgl0ilW7Roj0itk
6kaQjBdj7whOTmC1XdrZschjhXGPot2nbUeHZ7Av3SEegy2od4Rvak2t3mzUZtlz
Dm46rsmE/2XKzOJ38IN7Z2O4NnoAIejhgWZt7mVx8WBFeOBeGWE9vQTS5Sf7BHGG
tCuxZ7lWJaFVhhd52JdIZ7OsGIpQ+KZCrbvTgsJRcXhFQWwlVaFBCPqlJziH8Sbv
3Xjpvbnas1rhtc4SW1O3s4+wlT4Xc1vp/1kwTTj+hpwxWQ0yasLgDuMld5wtcDJ7
OUJy0Nhr797NmTNY6EXB7grOk/O52ty/4RI7ZlV3E/vCBzkDqzI+Obd9cixib/uX
I4snIPQenjWETIP8bhUTQcVmiNbNoiI7cByuvBsm0HtHd8OSzurFcP7fV04AFeg1
+BX8uN0kOEI42xN9jka+U1Pxz8h0TCVjI/tIHPU+ykSB+12SnWmKBfj6pZP1b65v
KdDdVFGe7Lw1QIhAk7AmrsDYZUa2Xmr+dazcSuuep6ta5IQYdOMWatwmL1LHnBe6
61+u/PU+PWHJmhAgxzajhjptZQjdA9LJU9WP+EWHIfH18D97uXxmhkdzaxdZe8PF
yl7l+bfHtqW+sQhCFVveaZEm4lBG78Q6rppDhfGxxqsVSsP2XCEAJrejTBY/Kxim
p0i9A3R2XJ/pOrMmiU9O5PV4gocASYxCnrAj26yBnQym6vMmfbCeZBd1ylUu8Sjz
47T7ioVDNxSQ+P+x9lKyPANVQHXel1YvmsUFC4vGgYFZ1RLL5VtbJVJPD7TQllIh
AWuFs15DV7A/vNDZXc7NobTII474vw0GYOzQvPZuR+r29fBgLsCozVLvQtiDB6kF
TUm++DBUVkxt2GAAzX5LhHJxS79OkrCmvnd5mIKRarb9GpLWrOh10mfi50PdJUW5
Qibnial4iu0CgVguqpI/p2kWZt5w1NS7VsuSl7dgchXX/xi5ukl5HIDW7qBk67Wk
FdRqGEoAbzgIhH8M2t57bJZxGXl3YN3GNRiNpk8FKqum4/e++RNQW6bM20dlIrbz
jBPe+lCHwL2M8camBaAjGmKtztY9AA3+DebUxD8pTvHm3rIJvmA73sNaijgl0/2g
/OhgeIoip8ehLBSdO+p0nDPkI3O+vvTW74PxMxyI+z2TGuqE5HSC5Qk4/4+73uuZ
hL8+jvijTMoHFKFIOsB0Shsm8BAbsD0N+63hcLaJxCGnnGrVdcZiP5aKq5ikUYeb
7w6omt8/vf0FCgxabBrG5nligDNphbkB9pygl6yIdlH7mt18z5gfaWtn8AikPGMI
YVmKDdYQ+dkYP/1+uP4ZVHpTdq/hhC9cAiwvBUlk40KuJSzvaehC9U5rUD3YtTc6
bSK9JMSDeX/crO2x4fJSVp8laGdkgejlAIXpA/dw0AtJs/kTPyAqSPCv0o9+fS3R
hWbwC01hyfA8nHRzzsjon4BhImxNGecovXqCwHoVuX2d1LcaW0ZkwGkU3zojTqSi
9KrFh25XiOZctSz6PUyWMKWB0KzCMfXdb1g47ZUkKxWiI1bakBtVewJzDhV/y5su
/6kuNag5cPPtkxI1hax2ZPPXJx7WSgn/86V+KUp2IaQaHxqaUVPRztL9eEfDyyV5
3Jqu/Po8R729Yl8Z4dowSmRC2l5h3GoeVhEqn3cNsUbvHKpr4P/Ko2oB2FLYsQh/
tkcRHsxSqAJrSuX9dp7wMSnTWMoOJaoac5zRDo2/JAOltiTgbTT/OAk9WfSUgC3K
30/A1+xkpcmXJqdsk7qxTjLqDvkm/9ICjwiWJ8f401fSv6mUER3xFXjIsMYGIrbe
fQ8jx1UCQ5FaAH66FG7DMX0ENCRUySNdzKxdq/fdPbGuXYWrBp5AvToLny+uUCFX
qjFw/6mg9rVbeSuJKHCA8F3a/VkgPEbmFjmrsL/05nHKkGxLtQlPMxfG6Ye1IAhe
6LEIBmTsxuwu0+lT+awRWFUjIkCwOTwZGCUhwFkjeV5NvJ+ufgi9bOqCq5Q/2aSV
91Ejh72T0UPZgwefn1rlLrBk29rUPqEQFeMezDUkPKj7U50YA+BcbL1y5k+sJEhK
HTdBwSr0KhDo0G8zUqADFW6drW8CGRAATa4guCpjggG76fH0Pq79GsETrNdzmgns
y5L/oEcDtQiJSnTD3DwCazlrQ5EdUDEgjAZuxhFXig7BK2kR2NxMSiUjipTuZNL8
NqfzMyXQ4YcE5vaFduqs3BNxEd1nBbM024p/jbSJ4uYx6vpYHPODFnnM/Vsz0TDM
Avfdt7wiNLJrXR30EtHfBSdaEZVzU2RaccO3cv43WXojifE760hMdejATBsvPH25
ILt4SDgajL4SAvrX8p+++YpJ5zVnDmTCaPAjnPUrkxvHK8mhMfh7YHFU7krY9Dri
NowLgwMXdjngoELykdTMIL+Ex/9qAOHwbUqYxMzyykJNfX9AG8o37PY8eszL7FSH
OKJVNVh7qOvj/HWrR4FGKsbBlxGq9IG61XM6I4pUJyfdayZlFMqYqflOB3bTs/ev
Bnt9Hx6i/LDi4C+7pM1nYWgPjUwIzXUo1S6/cJ/B0o6OT8IwqbZpoNL0FDiTsMh1
VGHHXpJD0p6yogagZ6BRg04nnWCCNp5cmk+4cSqdlC9aw7zp22cSR7jgZh/cNwRI
mSzG9gaIW6jVXGIT9gjmkXuZcpSNrACDCgfVaoRlQJMCeEr9gX9QzOod6fxMo0gQ
IipQbwABj87lN1EdonUJ1k9HIWyscB7hPQyEoq8aXb8a6Z8+WNcAvQghUJ1RSu9Q
xLtUW4t45izweeDb3NsgaabdisVILj4mnNAUWoLv8NOOA7iq2qhIoXjx8lpEASHi
YnSI+DNQJeDb/hH0WrcbN1ghGkCCGZ3fGiKjgHXICG7yNRQhPxpIqI1vYtClFrsF
X8ZOixoZxojQrlEmTZsLXdhhcM2y+xSNXifaTB5xRqH5l0CrN9Pgb4rjCjF1HVca
3pyonqrd8h+0+t1ML3wb7/rHKoY9feqAedLZE/iHJqVaQmHYIza1Um81eT3rJoOW
wy/m9MJgNGT6aFRZA9SawpcNctRJ1H4d6XaqN6oZNs29599bZyQuHduUe4++CBWP
dfGPFKkojxBb7n9dnsZk67sd+U3SZlBitZgvDbCLwD78i5OfmFdt1/azpNpp2cHW
ZnTF7NPyHXukuydPEN4orTIR+3KHJx8Em+CKa5DR8EWpZfrdF19j4cf5B9gdAOho
9Ra8z9GiW7ZYFFjnbf2sd3Qoc03erumQrML/Qf6K8X1c6NhYDlglD4Afabe5cQbl
FYWjNvwKJaJNF6TzxuYBHH/ZnSaOG7YkG+KdATtfqpcNUnSxE6jqfN5sueNjzyyG
ZPDJ66b2RO690PTaV03tvSFeAIXCv4qMlxGZdlPAMgoRMJis61AWJkbYdHU4rB7j
UR41H9n9gK1XMvXSNoNQzLM0k4vmd5T8MNtO/EzRYoOqVuL3sA0+EzMLCRIVSChT
x18o2cN2OMxAboO8RRiYkyZMtWRbEnrzMUzUi2+mB3QSUNtehczRVOlppxdgj3GB
GrjqYaRhfo3b0ojZ+AIeJabEp/jicT8DMe1LctVmgEsGbynS3l6W+SOS65TI+PEQ
iFJmdqDr4xC0nndYdWTcUqUYZow4qD+ELfMcFRVfgCKNot+4zLwh+jnzM2SugskJ
YBs988ULWXb3hGgZini0cMAxKMb6iWQwvfUT2+ADL8NLuNPDOKnW4tWr3TIhmtIE
tioRBZtG4TAyOYp1Ere6C2KNdo6WQNGSiCDnb42HwnIJ6hKSYEdYcONg7jDTVkoV
5pL2kM0sdY5JS4N69w9jk72CAkPvCFk8qDh/TWWEtDikk+ceRsceX2XHq9aJ33WE
NAylYzQtlD1wbR3fP7fjOjuzIjmNHhjW3QEPJaLo9furU4mVh8el7NbJ/t8eoUxC
3ZhFXF1xZzfjIdvh+Z7vkj8PkMToeYjSAzXb7SiNNCkPnRof8knQDnLPHzaU5tJQ
89igFNKehicHFdVxXt6w1MeCDVzX62xVgUgHGj34iUFEZukAtCjr4qjPv+Ze9NMg
Y6tbx75/v81OM/lell6+iLosKAuWEy7TYNRaPESqASWrZ90Mwz3I+ikK/qBae/Ef
KNcIcSSVZy+rZcsZmQwJNTFSNS3kdoLzgY0t4sH21iiajX1SWpvA6lYJnDGP7Enf
zHRnyvOOR/rjUzuP6RPHMyCFvKKq9edY/mAt/ZoKc6fB4Pgm3rULO+k3A6rRNqL7
yla3uA1+QOutErvJll0SKuaACaMPWpdARm2hY6WUGrEeiLXME5xa5ahHW89rqSH7
9TAS3K2TVjhRoRxcvNQcLM/xm7araNEONgIH1M5u0gTgsM1YF0ir40swdntPXX2P
ACcv1x+z5a5PxoV6mRRt9Bt3tzwPs3bPU0wDrLoOzVpO4bDQ+b+JzyQVn8GSqtON
2+3OrIHE49yL3jaI83PNDLZDjXwC/DsAPtDzcvkxgPsWFCafskTUChKSRhq/YtKA
o+Z/pAij4LajU4lOIJWeMtD/2mTRzSbaJRjwdutujKVOPlRfC4QcOW6iA9vT45Lu
co0dZ4HykxZrGboNJEE4yu/42uT8Y+pMtYtlcHAK0v8nnbGY7nBVj7OCGhqNKXDm
BQI5whejV6smnsHW6tcIiL6LQU+d1WeODtMoEWhs1WbxQ8j3cqpuW6Fr5V1neHEW
gloEopJrtQzOk2mmxpZB534/IsknhWJPshjm8J6WuLo70UtBe4U3JLL8wZ5Q1mDM
qvOrrbVBB2YxfPdyHQjL512Rep5uIrOlk75x5NbJN5hWdklLLECTC4fCACQPPGjP
Rdhh2g41/PCxFqv7WbHyaQOBKK+pXlBAPDWKDztLpq1nME+SDuMoTvAEQ0PMhJda
uJBkQHuTSgMdyNzFi5ixjaLJG7FXiOwvFXBYKYQ7XlMn+jfeqnDaishdxPtfJTM5
W+7r3k96aprHE5lEXoX6uqGMYWcX1yJboBmG718bOfW8emt3YsqknSSQeog6xs9W
8PI6UeGCiBD2t7JGEutKKSzCdaCeQfupvJLDxpxRmog8WbLiFFHRxe83mrm6axxN
DArGMp5uB32WPZD65Opk5exmGVb4H0QSgt04yqDZJ6UrR0v+1QJiG/q7pIPsMgAk
bNKnGbN+QEuRqQRWm5yPvFFEksevDuuXSi92qENSsSvR+Klj+TVoAjm8il0xQk0v
+ckh1JiJN6Fqj6TnXT6cAt39U3lNdUJtpoaKMDUrOEtCRaj4F3j6LYTwkAh4geAT
wY+rZ1a+0mdDc7RyJvQT7WDQRYedK5nWVjjo5HdLTy8kyrVG/+FJkMnMSvgU+IwT
Q5JRL3S9DWSDla5ZIQjWtGuyPxLSB9OHhAKQS8IiLA8Q46iLXlJPMkLG89VLeLD4
JDLvigfDr3mpgkHdDt0m3WL2IsBNlr3vTqYOL1vT+HWNqleOHVEuPok8pJ+09MoQ
J9WpL+vO31ZlJJi/Z89sGHydQOu7TX65i8m0JkMyVZ/1vp0vPPWD8LhoI31H8O7D
Rqdzuljwr8jNV5Z2D50XuowYi+wqqGjyjZaxeEiODzmpfCc47V+Kw8H+nCk0n5QR
5Ajj+IzoDnSEwF1fUo/Fh+Hh2JdVfa4bMQLdVMX/+l5EXWtTe18DunbaTU+jvTLI
wsKRBbg62K6aZtDLUhkl3atRvW5vomk/GJ7nnhHMYLbPU5DLoiCmjWVAH6569ebm
Rg2oqORplTnwPJT2it9M7rm7FP3y7f3UY+uIgit/XUNDL/zCQ8qh7TP52JNy52ej
AiSCjmanrS5kmJ3Ek+j9Bf2rSk8o6IvI2kU3zKd5+z1LDEwbk/2mFLPNPcm+3q+S
558+18nMn2BlpF9pgaAbujctJsMv6LJtbr0paCQpDwGjc7GkZF5EnqG3LmoQOllJ
vy055w9PqJDkN5P/qqoR6bZu8Nq0jxShcPZUSBBC/cUyUpzYiEe0MMiFS2XjJI0A
nfWZD4tBvLj/QN0LeSbA58Y54/oiSu6XhN87ELEw6NbNtLlUPr1gIeEX4ZgRNJMC
kqxUBFZGQMI0V8uiQp1eC9irGHcx1ZXap+35f8Lv76hJ39PGXJK/yhkMxNF4YmX9
+Mixb3Ads5TmQ2FTNNilqSqp9oHNI9v4rtZMkiotn1sktLz6JczoCfolEcRtWbtf
cPz96Mqp4cKIwpavRKGabwEUZlDkbFqQjZqQlx7HI2ndaZc1yuQIZY2h79i1JCvl
puLOOEuNYHuqcvoAdGC88w/PSxsGipVzxTal5ZNS+fQzsSUgxV0vVwyPLXKYBs4j
6Y1vizTfTjgrfDef0ZB2FRMSm6uuRp4HVRFRECyaHcMlkpN0abSjJ5IzDn22ETlT
kC3GDs5U+IbdIda6W/tdLfRDEXRkp09sepQY9J9BhMWBWCevyeuOVbgFUAqYTwcx
Y18aLGcotev8cXubxuOU3gPJit3tqCWQbQVea1AjM8qTcY8HHR+mNTrze3xFxxWD
58JnigkUOt5neJ875TGNywCNtVyl+tjpBf5uR3uRMWsD0q0+PlYK9PSU23pzsEn6
ApTUxlp62MrcBg74aAWB5QOD9CB+ESrrcmnE0nBhcJp7w8nTIwgtPcH2om3dxA1p
15e87bX2oWzewfxbrKaTod2QZM5Z+MHalZm6ZREOlj19lQ7jYLjLctndkv913ea/
1IPlQWMWiy+trFDc5Z2oUHswylQb7IGivqjucC2BlyS3ZIDwM6ZkgQO4RVyVKfVx
WJlPSGUj1Bx2OiycpmxXKBJXLit/qKkhzPX2cr/y4lQUq5Z50Ifiy78PSnmJYL4R
5GVNbPaRwsH+9mTmXyw06Kg5s24X3vG8OOQ13LJYJMjCpoYDImfgSY6/hzoOfFec
WF3Rc1/o34Y/+PIyHVEZC0FXB0gpto8s26fmwVALlMcW8EbnrmSdgIC2zec6nkVi
qJJT17u/6ni/MaUNHTMdEO9xOMdG4rHnlhVmsxiLLpYnlPDeo5seYUrCJAyfbzqD
5wg03VNuQymAOCEn5tkGQQ8wvDyPNd3I6DBX+6oNzJEybEr9/MOZxFeCVb/MV23h
M/QMQaRQTcIbbgoK1Af8s9hisFeQ45S2ye+4DPZOz3QBcZbyoBkgbOWQ7posZ3tl
zzfhE7TZQ8MGGBFET0hnS3UJcgPO+lwrSbql7GOW1F0OpOPJ+6T89+00K/H5R7ZX
cMWnQuw4kU7SXe8Qg43kAzzhAG+VPF6c42volb+3jdtrJ60kBTu+cxyUXPc+g/uT
7Lxie9acJY0D4HBZmu3VMxQYl665/pgH6uLeu+SZ+hqpXUuIm0bgbqEhHU3J9PTq
/Yr55dY+z20tcWWzg47e/ow+bW4Z5zYjbFRM6OdnisPjjAYLsUl3OHOozOlblrNN
pgNYu+DcQ0GED0A2TTjID4ee8xMuPiGjdrMBbg5AocCWcuuONr3uZajpSEqGD2gM
BDi1NtXt91KGRDUe14exbjFfqtDruNWjrJDEe9Iv/3R+T29BAUAVJoEf+DxRgVbS
WncohoQXHf1jo6MopyZFJ+z6WGMynZNNyJ3h0kmY+2grXu8GKQQYyufZG6rkl7gB
Qkfu4kMqiYiEJPEu2/QzgYRhWg7mJQWT4216pW4X1dnZv0bkUh842tRgxuNU3B+3
C5rSy3LD8pwVbTPY1Ib2gQjC2LUx4U9XXsssdb+QjYb4ip/i/rJwBKvUomgCEIg6
gLaupFVRmPvLQYfZCunXPruZ8offLRVR0wyjrYUqa5MujdfdFABEanH7SpxL2iyr
gIlgnolkB3nq6kHF0QKOKypoPZLZwT4T2WkBss1JNuyNDLc5lPCYmg1IOzp5OBRf
7yOi8Fz8Aon7T13cZ7bqphp5myE1NE1dGaoTDbfB5zy5+LmEkyyF8xcN2O1l5uQW
EK9j6z5mUzIu94rub4o837tswx8s4b2n4uoQ8oVdi2QfP/5SDoYfgu7glRadBTY3
74ptMKs1m5VyyqYinaES5Tm7XWK9xu1q9qABQovhk7Ic+VyRhM6Eq6zq64nrQMRg
K9wVdYyTTFwaCejLjpz8hMvbqi6jBmKbwaM+Li3Lns6L5WqVFW6Ho69n63Lesmdn
EM62GL7WBVa3LqzJtEfevzdICf1PBzli88u2yUJZF49ZdJ/5ftzn83ZjcuEOiEb+
HqlDBx1XLMTfTU6eB7DqgDeA6juRIyeSkFpWHxPsWRGdYU9MZOVwObVZ0BS5imu0
nf52aTREgYQPdUSAlGZtAWCcoF6aCpId5BtRUckZFs3I0RJrRlmZxyd+zUCcwuOd
3v/AwnNusXfmGP3Rgb/fSVYrYdP7WuBQLnWEDhgjAJ9FEI2iGg+GpRbJxi/3UAUM
5xDZIUgF6WMgGRGozUfYs2gCsP3PU6BCPJUKsI1JmJNux4OeUO45rWMVtgZqLyTR
0SimJabQyYOxmFdTVkEVCSTUtbyhWilc7A6mG1ZMSzIGt1b+JWjGzD0U7bDhPLcd
1wq5jAkvyQ32Hxi5g9FENf5WRJHDP0LXcPjy0aOajdW7+C5F2TDwBOcWTZySuh/v
uFtbc0RdfDFcuahGdfoXiJrIEdc98bUk1Y4cLyVl+s8+qMvNSexIwVzaXSLQ4ZsZ
VursOSxrT4v+BOjwqo4h7WwrrHHqKlItmkDHVleGojn16zAcZnx5wnLdsZemmRHJ
64Yp6Nj0BWUwZtCa+p9Zhaz6RBPRQcppLBXhXglhIGTSokVxA8B7mS8IZOnzl/i6
wmBEpglYRfIHoAviay63NDu7s8Gjuu+eCpn70JXUI377kEtGhUJu+uvxaMOAmLmO
eEMMMZjyIqcgp5VTCGONFa8b7hbSDGkK/qorVgSvoFRYUha5WxYOruH6kOAa1FbZ
zAGsAEg+Gn/qszHzRme1qyfEXXfRVISNv0n2gIJbZSNPwKvDwn63pJdJgPKsYh9N
+9TykFpbOVWMtKtJqDZTt/W5C6tsNlt2enKmDS7/pCp7S4/5A6S/fPi3r8CCpsf/
RIXHJjG6OzbYUApFf20HnfjIc5eUzxO0F75BMy1eIoQEagyoLMi+Gz9clGPDLo+d
P1TerdQD98bf9c6o6ElHE3KmPmmNIRjGJ1mwA64hxh9CV1cQuX0L3o4M06GkPZs7
pJTSHlISL2e2Sme0Z/XK4I6BXF4TXSf+D5+KZqkt5pXeJ+hokl7l/UAS2MKlXZBH
VJXb2PgtOBUm1ibTeNH/4JxFyjT/dHStMJ8Bfn7C9XUfx0yV1C7QMud10NyCCFL2
SEjOqUk7MqsBXp8012KMJ85H9z5AeoqaXFHBN1Sd34RxHiMhY5o5QtAGsaXtqF6V
8m187ayUzcHUEdrz2aquWur/36ce6akRSe/uStrFyt/CExJxchXXY0MDA3BlSVfi
a8frbpbnhz3Un2pymrLIasM/RlPXBLTnPF2ZNpqZsRgAS+niFiU6p+bIULWEUep8
PMWN0bkZpPA6R5uHcEROVazFrwlw4rm5T4oXH/JSxIIPKW8YhL1UCOJWyPtImqB/
rpq/+LOwMpgpIcOVMr7PWvFJHqzL+FlGtYOTqeNiCFZcppAW/TKqTihckEFPBx/O
HcP5TBoIflKTHhGIrNzYcShowxazucdbsZ+K9LdRDCXD3w0Lb8+NMo2xgWs/0skI
fGXdAeuKl7TQ4zP8Xe1dw0XsvJCDla9iMfW2GWZt3dyLuIH2ZX97G5tCYMfxJddJ
z1Cm8aCDmEFzNUfrgfRrwAVoFSqc6NTkFBE2X91bTEFh/aBkX7mEgyOzrAdYBlp4
mUwVM57Gmhyc5Ir1Ju3Cju/Dgx7QzCwScToVjPEervsTNHcfhu5lOJ3Os6lGFNH3
TR7PoAb9Y0A6a/Yvt+tStvpYzlbaFIow6bRql2NyFONhfHEfLmyNHZgvuY/WBaKK
l4ANKAfjrfzFeaIJmEhXt+CEjZkdjKZG0r+lq5BcNqcr5/BXvzk9BuPDeRdNHWIf
SvPvBFwUUzmZoKfgKfpzZ7QiyE9qLpIZgILuxuilf8MpLw6RKCBOrCtsuJlOVUek
LxxRwK2M3cHhifvm/8xlDhymCzxKXGpVYOwY33ti/gUy4Tbt+eSN2e9BHi4rGAt7
+VXJK7wsuYo/fPRcAtJJmFBM1VSk76z9MeqRd+HtXWqL0WHUtO2EXWxkQyixx77p
Z1LnZVH48H32GLviXjVjnvkHAOz5jN92rAt3wqnEt0or2D3LkBETUyk1aIdrYg9m
AvYAxjf2lb9CSzI0W5e9qjVf0e2rokyRNX3N2wDqQQTdXWHKyW+umJcfLSfL2ACy
Ya70zblSSnT/TU9GiPdCUYCnWo5hkI1p44GAjRQ8bVxdvSPKA+iwNfeGnB1IGC3T
T0fyuajHAh7BhGUQD2c9Ssr50wDnTmDj4dIOcrxchnYD9I090Lh0JC03Qx5/Tq33
956niCi57vY9Tp2Okj5wdVzAcDu2O/zQtBHKl/QLxhG+Dv0uoUzf/iaKI181wRBt
2TtVSXI1y6mCWXVnv2excVzY7YqvIGWt+dPtnzUaGSoWHV9ZYdx4kGv2XikwLWst
RZ/AaM4M1jRxpK2454fnyiKiY8PmFw09wkShFMHVTT3psV+KC77jP8A9JZX9Ix90
OaVLkM43ybNhNO7EqLISnKDe4aQOZ9nGzy4TEpHz+oLqhbQveAh5ktHTAuqFOg5r
qI4DNxrG2qyfqRBONC+cTgmq5TxzzBqJJ7b+WwSj2zp+Y54WVzFE+YXE2YXwPXWX
Yj3Yqfl2DpTjg2+c/fYWJdc7M94TdQ3X1h0Z24mpVWkdB92grbC3rLxhHGA0nDwK
yQzWbUjUwMM3YCo8E5s2FPHDtDPYxs9urQo2NLFe791N0yeMR/Ot0FWm9Qu9dneb
VOhjf3y3tjCuDmje8tUrOQJABJ3yoPJqHj0N2Jd5jpwJinbovZt6hZ9myW7/R4uU
a5EFXfCg/US2rSC04nVSwTEtk4dWuHIQiNbfnCKrZ1MnAR7YB/Mx4IFf71uSxgo7
EGseoTv+JBHkPzw/h18izalh32oA58HVFVSbz2yNKTPSyYxqRRvA/dRD8suqC2pB
Spq2X5mVaXWzkQCYbvK2gK243slYzq0iufCftQLGE3Rh6Lez/1eQhhBidBT21SQc
Yw92mcPItbcLorv9sTzpZ9GjZ0USn0xHnb2Dvy300vXmce0JsDfIkQh2KXAcyYoM
gTuu8UP7aybLcmsPvxp/NF4YF+oYgzjmjDqQwJUx3MqAeK3N05slgDIvu6PBMjUO
lnDlqj5GV0G0JTmOTdTOmqYriGYizB181HJ+Zck3NVoGzwt2MEDgfbKpNCEf7ymI
ck4wjgIv1Pv28IdpCWAZ6Z8jGLB6KqnMISmgBPF++bSvpK6y2rB6N8fVuq7IzV4y
BOd6VaEb1ss48ZjkDKp13GSV2SqFVbVfYBdgvmF8f5OUxSsVqlene08qJ20Dea9r
sli1nV+3XOlpNoBFKPKniVmUVmkKlkE64aboxUQb7+yCz2gFLAcwMq/lNdtWV1Hz
wCnrtRe42EDh2J8no72xs4bPR/A0eP0b9fCtPyfjj8t8RMHbtqcG87jJSocCynta
+KA5RcBjXfRe49SUzyVVYUVy+Z8LCkn09h1DJfNBSQUh2KEEU4+WsPP+7IUYdVKp
lRzbQLoXAPDxfc5WWmDpDS6mpO+TUZN4zbVqNYejHm+yIFQY4ktqFupSXMdWhqXt
qui9KCLrG5cHohg1P9B7ICdSTm0ZmIO17XBrAR0ZkTMMbPabVpQVTynGOwbO3bey
R2+4gTn6N2UiDHAm4bJ6n3gpED4xsu6fatbsyItn86VLXmtkLPa7XfyZKLWZjUwC
EfkEpKFr7IoerEJGDE+XVpL8m0zyLQ3oZixbu7hBwFUWlwTAYNu5QCg6twiaUAkP
NsFDyG6MBh4VIhlBAsAv/1JgfjUfvL+O3nD4K0AM0FaBxwucRfJRp/zJy5n9lOtN
aKlIyjvvghQR2DVtvox5ZwHJ0cGz3jTimPCO2AVXwdSQXHv98lalhrandhcDLjtL
8wybiZtMfztcJO374BIy0jQoa3pQnesnmw8vInAoCDVM73KDVyq6kSUki6NWvACB
9XheEsZbkj8VgfD0JFrPV8nlNAYgKwHg6DfqwmLGuRtP6C8qJp+QaZh6axdjLSCM
BfTt6pKHMfJ7G01yqYOXcRUcyvW3NxE+uhnoAWfakZqW23MAtV1LCPeGkG1mtLjz
2arBmF9J9jsc3tiARo2cLtzm9IrMOZt8ZMxhLbkUXdxwOtT1LyO6xC3OGLi9aV4Q
anKbk+xbSvv3MuMTxoPYF8y4nfl5cMiQI3oKdUXhKJXBJoB9QPGxxdlPg9ywELGS
3tfN5m7vU6ATMmexQWUznW5RWiJlEpTVLvtep280uPOF3OKj82GqCc9lOwE/XTRm
/1mFpO2jzdPgwdJ32z1+BciphghGpmkb5GbpAuDqYGwtbhCO86wu+Uds1VU2Vtfz
Ar30kXs7UfhyQ1LKgJImLlE32T4Vc3vDqeVq0pam50AlMaG3BSL9p96AfGaNkCGO
7YhhaMeXFNFqPvE28GFlvYexeFZ+zAxnXwEeWIIv4WLf4oFi0PdsTv3CHwsMa8GQ
kg4gFGWDea+VwvbSR/oy6iGESlkHerD7Mx8B3a43WFYlOf8Xa//yNYCz+7F19NcO
kXtdJmKn/MolxbwJnwr3zG8Qpbi+yH5elWLFANAi0HiiWz3esQGA8Uw6Y5jmyIWj
qmePy7jzGZoJx2EExgdATKoFCdZlIlJCCBS3OfavXi3dmcTAyI2OFdmXcq5u+JY9
JdDdZmCJ/Mjm8D55oSk8IyPO4j8C8A1AygzZ0JlFrxbSvYwyhDMiK4v0YQmpQLqo
CPcVtSnCs+e+WbAmQY0rHwdutszsuYLaWxkcFzNKCAjHHLsMSQzgRlVnTARpb46n
2VDjARXzOU7S1s5mks08fxG3Hein59xDcdJ2TfAxvfbCPvLCGC18X4hU728sDwC7
9W7WNYZceuBCYtdkKR1RS+Jfp75KKBVvyNRBJ7k8E0qp+C79aH6H0FTRuFxvyDHB
DS84LYnhB6/ht6/VPmIR1q2DzBbnTw5nTuDYpmZT5WNPVWOsl5LAhEiEO5iyd1Tl
n9oGi1SffZLWsOx96b2TMu291/9cclxbn9GRCOyT0Kw/p0hUTx14TpScuhfa6mJO
uHG+im3uXFmZ26+0L8zvJ6khbBWTywb+3h7k8lyfYMDZ7IvYETsq9saVebg2sEFI
ipMUywrUF1cnmC7pz3+sGLyaWElGAnfP5cRB6AAFiwdMGmGiNRoReyIw5A5qeUeC
SxIDr6TIK9lx5TU23jXypYXV8TlTWHofMd5CvjjXTB3wFn8aQhLZKIx/MsezylKh
O100EDsLqfuPDIZGRFCjfHDICdRWQqe+D345bB6kaphvRFegrxqJBDxTHl6K95hd
nHyHe/Sb0EUIteCBnN2qL5+H5JcfBhC5vJr3A72CiAN8M/e7VIJp6rTo5baAR5ef
341YPBQ5Day3EUQFUkLJB/TQaA4d1n8fcYXEpOeeXe+4FfW4ounukwW5Zac8+3Ts
H51brprjGdGGtpNfEHFdFeIei2M1fKN1zz0u4c2lkBkhSGJs89N+l1jzxO0EMPR7
b1r4cKN5mzm5dIRj/4A5rrUQZfwJHjHYFqvEcuhCjdjnU+AcRGkv2xeAVBdWTRLj
+O+/AADtAIV0xj987qJHkR4KONs3HAtY9CpHUrBgncH3pW9bA2A16VQ4nFWqs13L
r6Kzuc/6AXju3rHvbLl1CzdObvwmMSmXHQPTrGmloaIakJk4IB4VHqNjwpWj0pds
jMuaJt3H5zNV9bPs/7sqnB8MXCaQmL3vhmtyMLTDdN6KDG2W9APJZ1OifVHpIoRI
eXHOFxBwSTly8z6on82WuPrh6gt136qR21iFfKnfZWg0mlKXAJN4GLLyG8fROjYk
UfxrTJc10OukMKUrzjvUlqO7QUtF3w8z8T5Q6c34ILd6cE79XSD8Tc+NSfAB/ubg
lNAZeP+SvekZ5N82Dymn8xpHD0eWbFROzRKO+6WwQaJ24WB/EvJ2iGsAGF6if+xx
arrgkFc8GT1TUgm6/veSsBkEjx4/aPZYpRvnmDd6jxZcJQ+UV3uMl4EX65Wu5YMs
irtLpH1GRY+hD8onF2klgrnTKZP57IInwEvlswlCGWiQWBEn/nmjlHvtzqj747RU
MDRsJDSWI6lZHZhTlXlElFiszJ3gQwsTyAnfnYFFFkuQ9hnD0v5gwwEznI6CtkqY
A4Z8+NgodQSw/S2LVQOT9udsLmxNc4l4d4r8JKcxRrIbD/4DkmP59AC9U3N67lZh
cpyQoi7QDuNJrZz6jwi+sZModr954PDIpX9m9YDFAFQeT1wQ/y1JJ992+MQJ6gzd
bI4bzaUwbxm9hgllJ81U5d4ctqEghijY+3kVBpK+7EQk0Cl6tT+2tBwwtYphY4NS
l2oqDI376YPYYHq7iod45blFdZecARN7H8d3xJvI0rHEpt6Um7z8xcfud3bqoby+
FYKjdIUteiOK2XZM0RO7nQeMJcApRMP/83+TV0+VmQZY5KuSSyTwNAbfTB/zBkTF
qf9qKTskoT1Tn30QkiO/l5hXDn4ezbf5OP0cm/X42EzojbDEtYO015N2LCAyBTqI
6vTtgMtupotxHE2x8X3pyT3tXjMeloNjgIGq58wVkibuKqnpVejovk8sMec/cvxC
sljoLwvjHm8FTsDIvRpcA9DeXeHpUtMS3Ntm/mPlTb4NXpIJw0WGM/NYh81PK+0x
Ihp+dXGuFaX+yBswC6pKEnmxINW3fFXn9v8mCNZdA3wglRgEB1hUBxx4xl6bOR91
xDhV4mLiuRVmtDhdmh8GPAl2mjbkjvbGo0lOriTKf+kmG7UPWy7VTp3wzymsYXqB
CrfkINDuEcGNnZfDBSBHJ9K3oHIUJgGSJoDDXZc6eQMcme8ugMl0OnJJlp3MQMjD
P2IW9G8dziPSq3ERHHXmvSGipqkbug/LXTHdwk1NaMIRpZPJYBtuCttz+Gp9W5LL
KmQcqxa8eAGxB1/l6qt52tnFbPVCihcG0Yos8rxFNL1JFh0fjyJJXUcB6eVNdH60
9I5IzdpIbngsHJD7O9U2xHY9IvEebiYHAokZfhTMV9pPXvGkvngnm2sSeC/m8R1y
B9WSVp7jlbazRy7hu9OjQjM4Gh202pfrScUmNJ9ShKyv5LNQDnqUnR/I0FJCt/He
p7hnB/+nYERVbokS+sjo15mqQMI/yHhAwT6s4XCZCU9a6k98oM4JkR1zfhn9x2kv
vAt7eeFZV9fEHBtvFLhGPKh8by9V/FPS3cS+D45RJ3xrSzfzUMFjXBKp8lVk+A2V
14o+Y/numTknuO6ke4fo15T0vePY4MbFyk/xwc47JPAC30PKUBqCgPNMzgCBCMPM
kAKde72xuAktAEgKf132AR1LFyeArTeJG7+IAag0Y9Vvvje40DHMtMIcHRVGCuJ7
MQaSYZCCPt1ffPxgpRL+tmsaMJF145f6nRp14ivknZXgzJO0CEcKKFDvVeJWzNQS
JJkHT9sX61wjUR8bNc1LbuVBLnnrE7zBSKRGh4kZSOYYwLv9ZzZaZ5ZqzJrNPFv8
nvp7+8WJ23CJjD69z24Oa9fWberz9XBmEzO+h2Akf/JuQO3K/8eD6bAMANrPQ0Mz
9Mn9/HrWXQ/1r51D1KeKIyY8c+V6fRnMG46vDejlbLngO7osLaVkAu1dSrRFk5cK
IyASNGxwfUHI1S8eRFqUCvv6qgii0XmWRMbxQCrbCpQTFPFnvXD2WA68PaU4KUv2
hy/qTi9lEIMgUiOBYxHH2pt+sKq9JquNjXtpnEQhSohvzNiO5OD7FedeTu/dYQSE
dxRlc2hrApNkMDFG9lKJJLq4UjkEgck5iQTB8PsgM0drCPZMzkO7Qn89uegc9SpA
+h2dPFcMdcVn6T3ycsuKU0oaBSjbdneXOjBhEN9hpGz/baY09b+UoHN1PtMzRHp6
VLkxwZhjTqj6eCu/fuCmvpMtuTI4zVW3GDBSJfKR/qj0nTLGDEXIdxfQzZ9aHVyv
0IY2Ntlp4khvVtI6FoutEB76/HVjvoa3zdqvX45+Cf9vxA4pzfI6v1gGQ9XKDOhm
cjKIj9Lx9+/7iq1nDBphu50YXXQuZIvi9XMKQiiNdQo8iUaaoOmpuaQmdxlFeM5H
b2eSa12Qmc/aQIogSb8S+wINq0Yxh5dkn2cXrFCDbxg5YxDF0bclvlUP9S8KyBOq
Bsic8/JXrh5ETZzEg7dJkp6nTnrWclc4OLK+hwcyK8jwvSC4cIQ3tFChu46IBVa6
GB3mi8pnUn2jR6bV3ofmGDB4M7uwPLek0PAHXyU2Zl1RJpp8KbVlETp836zphEfH
ymRDJLtP1kMJZtCFTL7tsPq+Tql+posB9pdMXLK1rFZreKwzK6dDHHzYTXkO2fnL
HXS3Hx/HF6VexyCyUlNIyiV1x3b5S5CKveARioNrVzojjEPEMr0SqlKbAMcsIdkk
FjCKFALB4p95TzuzJoL9LyR5+UJwsU7oRq5d/0dw6E4kNadwT8h8SscE+xIWgAYb
z/rcTwv91XI8VvHP1pn2s1vfi8S206hwb42Mix09XHrCor5e7Jp6Z39bbv7mX/M2
SrpAwO/6ewejElIPMBBuFc+MYGKvgSVpSPLIRQZS8FLOoAer3BQHMR3g9HN7yQeO
ZicByI9Y5MYF+SpPazOmXJV9DqcqNiIbLZO5+JEfHvwh7EzEMl3PuQ2qkev7NJzx
hbmb4G040qnd7sHf8o5lAtpLaJwrBkaJMn7EunzNT4gvSd+9PG7dWwHSmGFnT6DZ
J+YXiANb2ByrFiDOW3u+VfVnecrl7Knsgg2+beDQ/DL8hS1UmVLqJywCY8rK7j4O
Y/jFbsnrRPbvoXbx2sQwND+Uetrkoj/UZzdhwSdvWpkS7YL27HNm6m6Wx8lAg8di
Ki5Fy4ZT299Q0uExVYAMKssKrj6rkzbMYTWsHET/QKt5/jEcmA+4nzvl9BERBz1A
9Z6NFbc5tDtyJBXLwsv35uJfa6G/QsPqynfAvzvX1ufDU+dlySMohdU2QQvRD2Re
QHKNG7mm8WcXGIxwZA1Fb+GdeMWl1lRVkfeQmnO5ny2u1wkfvaEYzsBtF+ZNdmj3
lUqMLe4TfLd3F4xPhuYzadjK3Ctv94Gpq2xJSwKQLNLVzaXFUNWLC4KD2zqHFKP5
CJOBJ61jEiHiwl4D8BfeCJKToFd3UpsMymK7aYI6FXX8UEfAtqcfZHibESVoVDbZ
Hx74uV3ssCGB5BIFTafXjDfHRQj4qmaYnqkZsFWr6TBB2ilUW2KF9A3cUsijw2oz
pb+WeOiwMZVcxhHs1w1robknGEUIq//M0wpIqTKkT0AfBIB//jiBzxlravCVxTnF
sAo7ZAm+MWAVcCMTJ1gmijKLCq6T4hBpE8W5B78EaRizkiXlF8asbfWsUlCC+XYy
EWWDr5TC+1YVOkZaeYORsbKgPhPrtopxxfEWDzCADmZcrjL8Ou9uywge/YGmfh/K
IRnb5jUqUl285ZgI8Dcm+lDip+aCQ02OiTevceLv4d5+iD9WN8/CaUWBMTMTxePT
OT18PfO06ahvBVxmpyv0HrLs1OUBcsoemF19rfrl4g3TFbzwd4pQojilAK4zdgi9
q9UAw+3kW0eXJHvfsfQojhQz+94FFxMs7ivRL1tU/zmljATCl/6KrtfcipuH2dzo
ERFoWQ2u5DV8D2myMqhWfWx7Uc5RbIasGDrPwvxpLiRAoAkDj+FftVOG0aZwEprT
o1oNpOakhoHPZ8KPhFUgWlO6l/YAE2xduU2y6YMPrtB05gutCz0r7P+IlMG0JgMk
rusB4P0YA/OiMiVfArBfj2Q4KHMjNtWeAITH0ziPhGyjKnV361NZmt65Nk4G5sq5
01VJnWRQbqQul/FzFuDC2Uysnr64It+uHrvLS95I65eP4XHDDD2UqeNj51YjCrhH
cA2D1F96Qd7um9cBI6GeXoentxzcaW7K4UlofyU+9Qau45IpxMuKxwI2FmU8H2NU
XHfLUDPOLd235kh9MStxkaw/B9wrTe1Gvqjfr9gJ/0FcGimcUs+DZWY/UaZY6iK0
cOZFWbMzOAGygq0BvLGc7qeyFHAe3SxREWAs+Li0wu3/ipiKU/D+EosRczqXo539
YL0u3K5kKsMULXA2DeLksz1bfX84RkmntoUhp/uIci7/b6I64Se9o9CzjjMLdS93
2yFWiaovRgTFGx95xqK0u5uVpLRoKtDSdwzNYrEjIRGSIjMhtSatvb35JITueC9b
b1xfvbe4nxjUyJww5jjXbCxRKUEl+9Ypt1qY/JW0B9dWP+BIBmRs9RJWrvAyOxw8
9KZMWcGQsamkT4UwFlPMJtYu8M6StXuQ1ru5gkWsUzdNm6G7LIxHe53HLCZIa3Xq
2R24Io/hR9d+9+B/J2qFIiuvxZAFPFzZMz67T04hWYgVUP+XVawmy5ePfYpjzdmK
LI2a2PDIN4mp/djl91SC+4C2vHHrBykzrf7BQei305WvpKz97LtWe4GZZhBnbAK6
ONAqAHa2gz//ElRD2deHXIch6sWCG7O9j4KImD/M44jJefqWgBFk3dQbzc9LkjLK
FFdz1QjTyK3EB37uuXvAzrpz/1Ny6pcHcFxEEB8TN31a8VsCbix3TLivMD5RhlU/
3fKeeAcXjm7ExGSVUokLoZzR50FdKP+GPH5zb22TzY+kTxGStFGqi7CWIF0P3X2P
gIUA9TGC+D47hR4sBaa8BAafiGVC5lNvWniQrfMn4aGWQHvDIS3h9NVGJ1wbXLPv
K7QtjHBCURbmkbBGubrD7yXDEl6c56x9+lFIac8rw8S2dGFCN5GCi9xu7z3BNcmw
i58Qb8DsD3AD55Te1lF2+AcYI3g7TqmR77UTACVvs1E42ZC/phcqvW3ljlcmkEmO
L7vKRagDF9oaUGc5y3N8UQe6wGU8cep7pFfuztqaBEOsfg/3FXePXhk/xe4zTeym
+NdBaHZInEC6qOpoqAxcG2X9Y2Q/WWX1NJcn2w5Yfx4oILcCt5T4ZWd4cnvvjsTP
CFhfz79TnYXE2UsLedts53nB5fswiJMjbXsI/WKS0rYwONue/pXgYYrOcda/N0+K
LLbxs8VDGzd7obhx6zO96HAPc7xnBvdpk+FzQ5qwSZtQZk8iM6wJ8eD8Z+i0HbSJ
OvXANmOq2YbEZEjxUYkuJzruVhF1gnDjvvg5nu5BuWykL4zyrFvJ3Af4u+b5wDGh
FyWxKV26gxsIwL5aVAiMxNDlg4XVthucoSiMVd0W+5l6Amk4Vl+whTWLCYAXE3ko
QAySDk2TQwsF/fn5V6HdFSimIOosLCwfomXS6svzgXc8QP2/EGd6cYaHIqn4E/3u
B3C3trp2OKuZf0sMLmjZqjNYopUBWdGTHhM935sGPoEl+5LdWSrKlYSbQF0+Bzh1
f6jMHwFzP4uWcmZOVKVoGLKu0xGcX6dhhtWcwQV+l6RIFeaSNb4oaVaupzwawNja
Ypa+Y34/xI/nkvebT/29jFKPUPiTyUTNkTZ1uesYlGbXEomW0YUSyh5+y663OPZf
IKP/1nIXYhx2i61JizNgjPpKYaGh0VP+0iAjCXAY27oAb9Ki1j5CTX4mbx6HnVXO
jE9XN+paN7gOh2dl+3IxBFHTEMDAiGdoOVTQ1wX5H8KMxSFrtbjN+okFozOsAYtB
A/XhRix2K/uHhgIznAiT8eZV+L2Lau0DPJjPdkvgRwnOKgjm5BMHb7OST3Lpz55q
fwl7EPIAsiuqrs393zFwntHj/wrmezC64gHEGulRIPK7T/ZlFUbNQfoKZVOa2Gx6
Yw+TQmDkgU8gGhgBp6pBvl/wB7lKXqX0uyNlE6efgsgz4zNcN/qINAaeWywcE3MZ
K4O0rBBrhZJYmnZklnnaC+22ilWCccBL3eJ1+hSE2AdeeCVc+T8CfNO65XwWpAjO
Rrv/yeRtL3keb7FsitTcJnOGFmI0iL9HULUhcnR3kXoHgkp0kF2wRrUClT7wz5kp
7Rxq5ROpoCjF9icB1Te3EpY6xKRW4EemzyWS9Leo20Ndjtr2Wdk1x0A5PuouQKVF
vITfHPk5wcUTQmCRl6qyniIjRJ5z/fNxk2hi0gZMGlI3+nnTDayrNB2admLIUtIx
i1MP4qpiLj3FXZGorVN/l/31wFmNyiIOT0Um8+HJVJal8ls7IlpvMYqkJlc9Ktzg
SJRr4s+tjALxfl8OhZ6HzxFCVxgTAddvuf+MCe5R75exzpm109l9PV/AOP7YXJkH
DBQGJ3MsJwWly1R2r0H/VNuQKHmMhAv+FMCkkfKwspTc2YJBtHA28TPItPUmS/fJ
QiVmqyRLYXdK3mKuiQfOPfGt0InhRs9snkeOV2IVFToSB2mq4w+C9etz6EFotyDF
S5QKViWgWbhfEW+PFH+3ql+OUkHnRE5mnrCdJTx81cqWA/v8PLq/5UvNCBuD/05w
GdIyDoa0VHzCY1Vde5imZDzTD3Uy4kZ9IsiQB9KqMJMxJuNdfwgYdxumsAsUzzxz
3x2TAipMKv5l5ndhPAqj0RJzMAOSq/YXwZYDhl7EJXJB54ltv0GU24LP4JvItibg
VJcaQ20vMx8rJpquJGLpbWRnU5uVLXNr8sGnnpQRtThxNWClLZNQLCAHYhTmfBiE
hheK8RmF+WAjITr38IKXSffPMQLpPMr7iBUhuZSCcKMG7qdTUqiLGf9qfsUHQDQS
cSqQ1hV0hippa333IDiNs0CZIHQp4Bpc+MCQduHwUuubAqsh5becM0tHV5az8ce1
pVlToHpBvUQ8H2KYkWNeK6Pg0TmhpeGvX7QthRYAODeSxDUzJ/rmPnQ8JCt+NA6L
AD+iPZDxYWuWr5Ek3KGVoZ1tM8giQ/RzV+ezG6sZGlE4ErfpxT+T9pTwErZVguxv
6WirECjw4EVHzZVpXgv7ckWipgkXRgW1Wk0fQ+DLPDy1rVjPMfPY9PihUYLpg1Ld
V/oXb0gH0XCg130a1fhCd+PdGs5blT08diLKQuW3Af+/baEN1pZY+hS2lUr5Boxr
lQq6v61fOseckMjAUxLRqE7f1FYhatiM5r8b2FejlNUSYHlGHhJZCeTVhGRrc5zJ
fqgxYHL0iW7PLcVt7xoiPYEbC6UpZZrk+MK+9iD8l8eNWN2jAQCj8bVcKWfUXW7+
3LBsAhXHt5fNqfe8nZJe5QvRxtNjnt2aJjNWO1U6CF6c9EiHsD7+xpjVxLGUOUbW
kMNrGRFDue9bvyCS/vmEBUgQeIvd3m24FOkmoEHG5khare9Ja32M+60F+84eZ9fy
QNK+ifJZ1orG1GftYwork+JwxHVzEmQyMLTeYOZmjQBuGpcGG8AOAGfIaSDj6aGl
cPPpAIf5cg9IYr90hYhssIWa/KCtwTtIKOqJ3OIlbxAL4INeO7RwiY1T5OjE36k/
eUmGn+e2iPZ1ns6cAbxUILfeTWLyUn26c71lEBy668pf5U3mz7qPBd/3pRHa4okw
PzCScZD/HKZ1Znh6otV85k+JIA99HLRIvguowQdZo6WxpaFqDQaiBPU6ESheTWKY
srwAOOvESVzUu+7BiWQPz6WmFLjjmV0UbyPAiCvopXVcvrUnLpNN/ipv360l4fBT
v9CRRjLvZfBSmPRmhadmsUfsxP5NO8wDlGT7wB29d0uANb5PmzH/C8fx+sPqcce3
RwohhWjh/83tkc/ilxCejqugCI4AmScdMctdu5iws91Owv4iaD5yIGzTO28+QLLY
fuDC/uA2cjKXCZZaP4kbufLCGoKPbX7wLf7BSgs/QZuZBYz0605cAMYS3I8qZ2Q4
qXnVuL7VspF70LlleqNljGF9yXejiyV6IGPMpt+28DU3YikwrK+fkM53qD5+lRa3
/aWGzTViVQfHmtgZQx98rZKnCVbr1ZGT/uYZIqjMLu0BdIabAo6Fz99TeKKMCnOe
QJ4EZCfCX5tDuoTG0opBE0DWDxIYj1I6TlSoVwSeal35uMqZkqCSZb940NzTxeTi
s8mnYBIKcRKGVJfmv/lrD150L2efiqhZGj8y84kikngY1C2tylmJenaF+9zddFLT
lXsZKm6vvLWLoWUBjppHi1oqS2kxpTppT4vzbF/45MiLNTnm7jDb1m+MgAiS7sBd
ZOGu4icDbcVVLsOqNFgKwXkb2h/kvH+9o0PmG/lgQV7vflPd7itj+6mmAZMYLjaC
3sMk0+0Fe8q9DPj+BV9/khp/vNYFUglravYS0ug5Maj21Pg1rjdCgdMN2tmcTK4V
kRZpMPW6sfBiO11icJpjYwXZiRbcmxhIBhQQvxEtvmWmgnn78NvravuBaZVzfRRG
AGLn6i2iM8RFogTtOrFdJwIALMVxpCUxdL0sGdfNf0H7exlrr9gMlfmbJqknhWiG
l8LsZmfBolr3L6JWXNVeNTojMtHPnhoR144UtxsnhmV9dSUibHxh1MneQb3Trgi1
0Ddn1dy2ZA1zgMxULt/dfoZVwZIQeHI56dqg/1VY9IyPFj+mfdigWPqMfP0ernz/
KrTLizZgx2uF1v7M3hL/zP6L2Cmv7CMbwf0brmhFny1E4FJSZI9suEA8sRPdSOj2
v0TlgH7A205Le01Ovyti00KYGXSCF8JAXgtQN+iCBd39rjB19mHFzRhoYZO+wrVA
95H3mMDfztzw/ULlJwyTXPZxpveOzMDOlB9NHxjyxrwb02lFUcO0v9zUZO/3Wkzr
Z4VGteGQ1ScRQX236i0eZyKuz5S4CMaTVsOfskA3zsBsiX5kN0+mA36nNdKzVTry
2HrXu73gU2QoU2RsjwWkQY8nrLzp5pbnaAx5ANAFiLaV/br/bOdRWUS1iMzoqcF8
rfOPFixdsbAnAdA1E3CJrAvlYkDnzO3L2FK05V7whqi9HVFumlPeCc+E4MaQx9Ks
THS4TUDqCH4ZaOPZ8zPRd6t1ZP5HTj/TxFZRZHl/iVNm8PSgyPF3ZRM57PfbXXua
yu2C/pOO1shNFdOo3V+VPwFeBu8q9s+9rw7XieVHGuIGTzDtF1ZrqA3AyR3/STuM
4HyH3kG6MIaCyWz0201Xs0sNki6jEc8AxYc61KCW+FIH3s9ricHsxQG6JAmL0OJm
PeC/E+xbuNo2al3R2FZ4WzJpv3gLtlrP4J0jTdMD9LA2HOOsFkzNQhQcnyNhYBRX
0yXEvKzXCnM/Avu59b+ckgOITziCPdKg+uKM18O5xeoWGP5gsT74NdHL+dfblq+8
mfbBev2sHra9GD4nvJqSFkgpY5uLaJtDbuiUjUMJOQH/MSQhNtPCzBY44N5dQysp
POgay08eflLX7FuRblhOV5WAtczv5MS9Ylu5LwHwoKjT4QvicR7dxG2+mLa+lW0V
18WUm577oNHPUXS+ke901mVVWdFUNGVOLfEbzwq9zpIoP6UQPwb2pkFaBhRiKg4s
Ur5MJVIjf91JGDBNPAaWPLmjCeJs+1UbrkZjr4NudR3OMTIgSxJplZ9wmAZshJtG
34cE9BA5zEnBvYKYbxJhDy0HBMMAO1WcUsvFaryAKnYYkQUBZ5/4FQ79QVusvku/
DwAg5ddAKpqNJ5vGS0yfQzH0uRyatPPQge5qdxAecx5p2T1alXoAEPWkjR8a07f6
XUsUWknL8yptBMhnGc3nEXEgEDiMLX2huj2pWZkawU8JXXShwplIh3UQPgqPIMIQ
6xNIwEdM9O0OjS9cN5kXI95tn5x377PyInruqpAWKGmAPt4gAg6Qhkidgqxsq+jn
QH+McfAxN6R4rvo12N5qyK0TrQvi2liGUGmbZa9v7VFP2kUk89AD+H/tU0WXvkle
tFZ5C9hSBiO3tHidN+WAfUUiqA2rzVrd06luHO1oalRCpyaLlxKMuVHUlEo+1TAG
j3bunC2CD3elK8vGPAzEy5wbd2felUoKLWos0evdbyNsgQw8L5R2JPkHvez8+pMY
l7U66PJkULdba9DyImOQyZ3heHesisCMBOs45lbcdHStoMAQiCDTRQj6DItStyEq
/J4P7Ux/FvXpaaoX5OVCopCxS0UF/TA35XEWrsu7rvusFnAHuS429ixP7G7qFGHU
2nw+J58VX3z9DJLlzgmrGi48uM8k05Yqs2dQVGjBsMlwCeU/2KQKXrsMbhevYBNK
SEigNgWNRRJNpF5SZBfPP0G3fIRjK+pIH9CWYcB4oKQDbTb/sm0gvKJbQO6Gzo25
n7P3DC1ZpQkbz6VUchmLwZwlJMSTlpfzq9UlmwmbgStnU19Xg+sd0p39boajuTy4
w7LC9Q4jX94lb5zL3dQ9nA/IRp8bROQPNDNcX2zKLnRuW0wrixbJA3P0GUs99fmi
H8PJT3tQ0kgYO5FuUuhilNZBJOwZ4U2XbdPPlwOhw7sNkmaXOQE4rVkX3ZXXUeRP
XHDfkYHZdKB3T8SfWL/LokRX3eVnlkva9VRZkz6Qgj8gt61/nnemvY18p/gfnFYk
kqDcBU6bZLVmQOhylSWRTtph0f1F2N/FXGdgCPSBZVqH7Rk5STTkLmNBWljn0DPJ
7npFQtgskmvOszNtu2rD/aN6Zf2Xhg/bpx9U7cWGiUqC1BP06vZ9p1vIrg9VSZJ8
JUdMfFFrJVI1zylc7OsiZgQ/YHORQEaAzAQG6HcA1a7+Lu5qEZC/ZwEUAw7/oA9y
N2OtFUEUDt7sqn4VcKfVPjBM6Yenp9XIPV7S8d4JWqYb/HWGnMISy+DOqr9nW9+a
rDC1z9MhLfajuvasTmLJ3A4er5YxZjUA1dzwPgCmEJB254XDTu+ZqR93JjK4x8+Q
TkQ21kjLfFMsVgLrcMMdmGUVtMuJA0wkv+6VjJAFj5UrveUCB19YztbttIZ2PP5W
O9reAWz6Md1avuKqnyyJk/EDE1As0i6AHwLbYDsNdTKJDjWuExUxl5v6F4AIGY0t
y7BRfXDIhjFOnWDIBV408mDCj/zYsmt7iISTmgFWj7FS0trPy5WIwiHp4jxmZKk1
6OgA/PMvJFFMg+ynwnD6jxNtCS+99gMFYH3fIYbO8WS+e9Rj4T45y4iYVfL21za5
RieVoOqDmxsG2yFiQmPfXSUqUZJaIonQsezC1Z4ZzOvQTSRTHWlQochwfuJzQvpd
HJFc+Z4KZ4B2C8WdJkP2HQVCI+6hzCU9c1rkrq9zrIqzgPk6skn7GwSQ2+7GUl9N
vkUrjevetoKA4lZ2V5lHOIEYxzjEIjIjjxUio1/06R6oTAbsTd4cJ57iUUJ0gmpz
05i0vV6wcOD/ocFIob+ookIa2pN2+istySU2TwH1op7kJaHtwZs5OB1RBVQFpFq/
/F5s3cE3HkPXBVmf1+qqQ7UMeTpZCK5xzqiD4sw0qN4C9fET9z726X1Ml988aESk
r22Ru25uR2fdABUIDDXEvjTerlFuGlF8ewOS3B5mJeoEOMtRTvYBxoUsWsZe5mpG
2vBwol1sfhiAahOe09faaea6Yu/xu9HwzjT1bQQBNzSaieAD0K41R6qrytPRHqG9
nSbriyUnJTuqtH8nI6/6Qbw83E4WdbpWXrz27zyexcGbsBbbarIBbKwZY7ObMw8U
REoG/jfwekAqld/z1SEOgb//R8y5QbWgE4c5AbB5If/g77pGKjs/h+4hlf2Llpvz
m23SeR3MsEFkjtd6Ubf6j3TUe0fhv9cfVSCAuJ+tak8fddZFk9xh2qOi+XS+uBnx
68pjFfpctYZcUwITWWFvbyetKtlTMVX9kq+/AMw0CZgauuQoCQdQG7YZtYpb6Ygd
rLbD6YRVxQ8citxTqFda3HX9kXmmbiDfDYFbThhd7XNA8nB1Bil8cxnLw0xpo+yi
y025bsiNgKAN+lBPDiMR/sW1UJqI+zYyUwRmSUrid8keR5J3YTm1Ss96wIcF0ZAk
rhBXJvKtr5sZf7JG6qCSrYm8kb4oYyuZ1YAKl/uJMtbxQDh9CkdVNVdofcOqoA2L
eAZz2ZjkYolbFA5dxNFKU+nw9EhwfHGaF8l9Q9vl4WFQIab8ldnqaMTuseOKPdNU
N/fE+wSGWC/w2L4ZGBSdBg0YzsVqXZt14wBUJRDvUF7cdFkcQ9w6a8uXBD7N6qsp
/ITeQ2dbZEmIvUYPdnzu/oenJdT5vpn1aYCUY8vyKUhwHex7pEm7609Cw2owFVIX
YYoD+8Xjc52UHdlVjtS1xQ7ewvRBja2wKG45Yf0o7Fx/uNnSmooWobg5PaiSQeqm
joxjP4fCEYnGjfQ3K1BckHRCOmeUXHCsBzIaYTkikDu1VOaLOjoxQW1KOnrRadKY
CZHtt7I17RPgl8PI+2z58ldZQkGsmky5MsyAQZmeFBCIlGBA1fpZbhyVXdRj1krr
UR+3XZzTA/LyOpo0v6nCAsw5rZgxFPWTC83nA1GdPybHgItvn9HKJPS2NDfsbzoR
THw7U+FZcvEf2/S2hGeMxySTx/Wb1A20zF3MeGfgoQMRtxz+OoS2c9IgovtaJxmg
vHMGLKw3za8zFlwukc0VYXEzlsQs15n/NQXpApEfA2CcxUVs6EzldMzvFc8Rkrda
yiCBZhyCpWR3FHvF/vTTYNJ/CE5PjmeqbHdTHmbzWR0ynpFbPkPYopfLn7W7UKz2
u1eYn4bOPzqum371CsQAIfTAd47oeSjZsQE0gVi+IACSuuXLIYTnqtEM51g7RDAZ
TAJDaSm5JkLyg9eAsHhfF2tRPB551c4Ku38VBRzvVY7bmSWq7+0lvB7lB/uFnzLV
A1QQeNt7RofUW6COzEr0mjsRUFVy5JOpB1LcLmxFUDwDu53BvGg8fD9jb1+GagQQ
tTPdvPUvEhrV8BkHc8LGU7FFDAq2KVNptguacjap3MmirLzBkE72vmy3G+n+tZfr
696/XhI5kl27nY+Hlv1N/bltudMT2E/I1Qg8OMh+f4otVDzlt6pbfhDvPeYImUzc
N5H+64LhSdwLxxDdN8sD2y92Tc0nRqNIpFnh9mSP6XM65RDICvTmf3zaidyr64Q4
p0Pf7p8AhDeg8KcE4MTmf0/CF8ek5nE3ecYqakXHpNjo7XvrpkzBliOTLKbFPmxR
7vHBMAcCct7oJD6hT1hg5fVQrxra6pVRQJslykCDR+e3hkLyY6braxq5sigN9c8i
162X5JxAC5/nazp9gBRgOR15cuSlpZW0OnJ2oH9mq7VxvB38GQ9VOjDI7CMlEEqT
s/ut2uCXRiXf8k5dxeGvc2eJQADmIe9x2mfSj748CIvIwDyWjpCUYQEjP44/spmU
QJsDw3ZoIpATKTU2Qu/CDsMfs8wAFlgCJFk1PG/6AaBcgjw9vmoyr+ElAfn3erKc
RGVO/l/hGumMm4/WFkJjlNlUtWsL7VpexDgE8UQJHOVJB5aoz7UiYrQF4EbjtDvZ
ECaJOq32y6ovZRmmyLKsoJSkIZ47gKRAHAYkkDi6hjTZhfU3X/EW6Wgzn6A4UQ54
OXZb5J1/hUI9nYdxEk3ZTeQiKHLwmrZAPKTFFaoL4/kowFmJ6J+KluqIEsgJqVCw
8cxyd6D7BO01k/Ofmzigaid3r19SXGyne2cZfxSn2x39qUBIDys87b22DpxIN6HE
ptuCJY4ALFm3NvcHIBdA0xtZQlLBj2k2rzEQbp6ZuJQ9SW/DfDMX/3qhsa+i35WP
HF9hbXqSPTVUr7BCyBKqMqnpR6kHUrsqe6za7xC1J9geWjEXK7GY0JIWdhvz1dSt
eLxnk39fcLyGpWJjY2KFTmSIv4op/GTtJQc/hD5soDmHnfubo/O0W1/FvKfWPYgF
w2aGLvowQZGqlg0REVPl6kG0E17ULYcqWmaQoXgDGy4NmLCqmxJLewjXdF5eTIMz
upfTdF+XKcJSUKcCGqCkz5OG2le1zLArjVOgBkSntPbPPdtqhEP3iq4uSvY/TOzs
RkojH/FTOyj4WcanZWJ3tlpgzTymI7nWH31dMFDMnkaUoHle9z5hLqhytXTA9C4/
Z+v08ZL83iyaJdNI/ZRguBOXBaNbHJsTLKugLrZ3xdkDMz8v9QOei4cQpv5+GIVi
Ue4uxQsXeR0D2q1yx1wWzhdD4SE5wisz8Kn26jfBivZQZoehNcJs052JWD1WFLAb
b1iui55zfyMUaoUSB46V6aqrffqpxkEyIWKs28A66fdEUrgY4Rk6SJqV7e1w5zNF
ekAxKCKBUyC5P4MvnYlEuAOYpT+HIS5iJynKhxW6rUkrOSlgNZZ+z+/ISc9QuDh1
xq03c2T01KctANSd5XJb90s44VT9FnnPEMA8DwobEm7gZlkO+Nswn/I72G4t2ocC
0QzraVENzi+e3MLB0HXGSmGFvzc9XgGAbNN+WT8cPaONEh5RK0rDNchs1yrzBPWa
j+sGu3RI+j/EFC8LKlbEkturchzLORPl27RMB21mZYKZnE+l1APdSkDc5/LKSJim
cUNdcWypanWZtQO22JFzntrjOisVUR9qHbc+hUEysUD3uO9NTobp37FjvBXgToXI
Ijpoo1XSovN1yk+Sfw69Wf3OJrfcP0DMRTQ3RcLBp7pugtRql2E3x4PV+/5rvxN+
NNTpV6ekPNgmdWGlt8jAUV2fU0ACdpjMIqYUou3AkWmabFss1q5Svl0nrfACteYc
lHslg0YucqSjo2EaMYIoNSg6HgDzIQ1Po/d+BseXQdiKHWj5ZoaJeFjkuyvROSOL
EF9yXPF5hwbRxMWYdinDOz1m30iG3+SWfnn+c5c6Qr1tY6V2WNMx7+/tznizKPdi
v8x94McPC38vpjQUDbwLIhRaEQ048gD15Ru4y6sb+UeyUcyIiRVyjPDUNaG4jDow
WR0Xe8INzp0x4DhHNcA6lqhnoFmg+pa2htlD1gAonYxl0t0La5h0D+6thRJx+kdt
nm7cDW9A/mVJ6ENuBatptPoWxcbr+J4TIJK9jcCke3NLR9hlwmX/EaAu9Nhlndbe
4Wg58fgMpX3XEo0emopMf/4ilCSnaXzZf55qhg4eRFh/GDh+IevBtpA5VxdUgY21
WkEfU30Y1pRXiUEvurZDkhFkhmHdKK80ybttOvtRNodVXInCVxVyGmorYAmTLUtu
lheA9VcmcXMIGUb3k9kHkWPkoRq8feBl9yr481lIbiIfKPlzpjzsP7sewlD8uNce
dZrh/F3TlCIik1FHLyhV1xwN0/76f51WYMlWlJ/F/qsDvYKCS281aleDEYcT/RvT
JJCPxM8/LZioGLMY3E8SkUnCi5hjf59SmAccyqJit+kbP2ZP+BYihpoN1wjk+zG1
h2qpyxEQ0pHqOpouznDINLuAGaBNYxQuaKUc76SytipTM0A3O2bVmC9W/WVtBwn0
dbHu5x3udlPCF+EqiUINHHKvkWt2WGA06q8TtrIHsXFsZlWhEoEe8lAO7vJgDkcP
WSLr6onRQbhGqvZyiLukOPy1n3B3Ohdxabp4OVoOeHIr8R4d0+LPGTeT4TPwFMhw
UiuH8El7CDhjvWMhOWs5c3i3VcuLg0O/zhZTgRyDFrLe5YaN+SSppBdwuWhcRBIb
XHp59VoRgT6IZQkzoeErNN2u3hJYf68wKBjokoCdnnFufXH/Cbl20eUOr4j+IOPP
EqmL4WIUmdFD4aopaNXN9Cq1csBVev4YgTUBKfqlEIKUFO6Ylpfn/912kGgw4kZq
YlOOjY3iI1xYh/7V1VfwQvRSzqOcgoOT5PGLGnTkaQMH+blX14hXZlMOxwnaa+X0
3bxrzpPGRcbWHPyU+O4r9Rj2uWXl82agy5KdpV8YWbYdJIXrPrkKNjQLrT2s8z8l
3xE+h32T5ZyqtK6OMuzWGps6YicbKAP6UsKRKjXRs8/xIuzYFb+P8PWQrMBdHBym
z7rSiqxkV/NXngo9SS3tO5GblNAKQ3RHi1Iy3Qfcz8EUhZdIV0PIkiB9xNRXbL0C
mOzWDEdTr8kdm7gHYnyLkzAOmxY9nbjsnld8n3HA65lxScT0jP0Dnvw2XIF1SG//
6BRH1XcipIonnWKiupLQZHvmAYthLmEhsdmGFKkzoyn6CqLRA5OFIjix2gGSDekZ
jHCxRr8usXnmoFX/hS3NvirpVvKOStGPdNS7l4UmHkvOz7UVvJ5LaPYGbzCBle/A
mmRa02Kjkde/oAfrSFxxtNpERkPtVtTHWrg1dwpygoyqfV5u9lzCGMpQ22UrAhYN
XKyImIXdz2oIyEkyF3Aqb3nugipT679/e6HQVyAdAb/cpZJASrdydkrpEI2JPuhr
JLwPVRfYrvj4kd2t82iDslJfUDMQrNCJaJy86QhN+8wlT65e+benFaOZERKh/FEF
35H1aAW5v4KGgQnpyhuwlGRidy8KGRidACj4RKEV7fJrrHXz5bNM2pvAD1nVJiEa
XJlpZmd164z8NTpQwqwERL8bWKuzMP1zjZoRiEimkTsZ+qdun/10NV74rxNB3elz
JCt1TOUL+eZsye1aHuOwz77HjbJuxy65X2TLgh2oQlfMabmdAVtdD7B7PHWzJu5e
PvLYxRsIXrq8vrkC+X5jqrIql52WRyW4SRAhnhdidlnWPf1RcCgN/Zx6J9eyb5Ly
NLcYB/7/V+os+d8xWAUw8ypwWOYhK3b4XVLjNi74UN39xb/VwEcK4XoM7EhCTE7D
NdzwJh9zR+SH93jR24H+n3pRq7Vdj7IYiaZLjrwF2tJInrZsbM3ocXaWNGiaP1IJ
chedS7SndaDJ4PE/S53bX+T4w68WozGUR2JyN/aRJTXEy14VFP+KsdkNWTEGF1Mk
POJxDFaqgXkH9PJtOtzHRAzhADdkNcD99YQDz58KOxpIba4REeWgF4+Iva6xx0LM
ZdfP/YYif25UsX8GAgJ9NoZMhQQP2lMIEfkhKm10W5zKne5raX4YZucwYbOELiUJ
VcrV0/5LE+CsjeMylRnUSShk1n/WGtmDzceaOxCYuC6rsN+/BW5e2w6lHFiL0qBk
nhr/ID/f9SSBBK+4VVf6frB66iG0rtzxiWaN/RDogArO7/LWIEyggOrI5o3sJAik
sEbEc/gJWrLF/GdmlKfBJhIn9C7kO+BT8iQTqDgOvJ9Vy6sLd1QvIOr29Kb6Wc1x
ykaFbrxycX+nBIus6TzGYKA7F//C5eYUNzO8U+mWQl7o4p1M6h3Iyq80JPGSfk57
N7o9At6FojJNNH0KR0nACIkZIyYeaGgS01FlrHhOExgrr3pbO3lxpTaUAxIXnTMR
1MxpcqPRn2eF1OZcZVZnv5jPbfwX5jLkpEcJk84vskbd/IelxJl/9xBecbdumf8u
ARaaZSQTjzaDVFjgsnd/BvqKl7iYX6wzP8OkM/uo+r194F+FaWN8Cr3IwC/fDBiX
pv84fzgzlgmbHAHpujpf5mP4VRYrhaIZ+MrejNJz6J/dmZ3GtnqKXAGXoVxBts7v
7rQyWLXvZdS/w43YO5kRB143KG7q1xSWFE1/0Ps2mwTPYXwO/i1QjXcer75EFA9U
t+pvDNbrrTN7VUqchI1ToOHSs7miXNltxvxT8ZGbZbPpMWWfH3pX/8q0DF+8NXug
4MV7GjKs9pUxmYgJEsQKMPjhZdYBPvGsztXNNCn35+JrpWMZRSY8ZP/tUP6VuGBM
rZJdxgrm7lHTQmHPLKrOO7yUv292xaQ9uzElWYLCCZ0xoVecEnrjBso453XRvY6L
Wc+64b3zYI+Nqi8a61RUHzks81c0jB3KVm/PrV+jQHhTJF9PceZa54WbHaqs+8UP
5S8DvdiO7Uh7JH1obcyB7IBITwQMxMZ9NqxQ6j2sniukoE9zgBpBNgkSOOmzt6S0
siTccj/0nkqMnNNCPFPeGVyZPVq2NJiv9b0z+IOwI3+2I/f5qTT0tNtd89RkcJz4
IG1baZZ8KptzZebaLTxtnc9W6C7DiHz5Wb4k7xTF693Nf9a6Z9zX1qgWlDQ2xuHB
CtASSSqvP618hr4k8LzCTR2OBdEproo44Uq7TmwC4onEjbWHFsiJiARp0q9Q0PuL
cTOXebrZgw8XyESyuit63cNGf7cOTCN8JkhZ5TAnSYlBvjWoST9w5uen7dGjT+Zu
Vomm9wl1DGNrAZmtWIPcEnAVnSrJJt+ekGni5Q/qk6ExWAQbFH5nwTTLDM1T9D+A
A1+aZylfPG3UJXvAvmgSGrTi8LqTZd+fRa+OO8ce8+g1U21NqBRLxgE5c2HbOml6
/3yTeopQjIzlzsL3tsIvSFEE5nmsd+BqXfL906Nx0cYZ6cjohv9PcNLcBi+TMBS8
x/+aiuSfx+7D9cGrLSzUFWfJiw4pPEo6wx/+JnUvCvMXGjKEASJUdJV089+B6xzj
MVeb+suVlbiC0PSnkrY+Fd3/xWnfxAKhpE9tejttwyy3qFWv9Bogiw6U9wHPdmh2
DQJxPNySDcK6i7hpZfIJiJ0tZT8OENEnEgOKGgQvOt2W3ikkNeQRhEXMp0GMzCT6
hQ/U+k1YTr9PjJIB30n0g96yX2pqXErE5eK7OSOQrYbPKyYmN3kfKwz3Vs/aGvWN
Ai6GT9tEWkSvMi8SAfkWW4XDafmFgBkOsRgvUprbngfLLzLICSVM6NqI1KqhCYD4
INp5GrD+m2JNbbyBttRXZZ/abN/+2ibUZo04jM3KXG6CuW9c9TTdGminYa/F9tU8
ElagBBIjNVBm4AuZl4ubbqOhZuUtl8azBdEFL1GSyCtOK7GGzNpFWTL0+HY5BQTK
iPk1BMX2b4qtAKwh+MKgo84dMgcI+ryjF8vEAGDSmCYKJaI+HYB/vohlXE+WJH6S
Dbwcs6KhsiaFNUUqDT/c5OZ7ftcLakLIW5xGmOUCR2/ExVs3gu1cYMpDru6Ihgqp
ppevWLowcgIXCBXH00n1Bhr+K79W783FGgCsTcahFq5LshudZ32jfaXXwBe+CJ17
2aFoW+8gyIJP2Xs3fQ+ud6bN5H+x3fgAeu2ivHNSaJUbdlbvVk4JYT8zUJ0tN5rI
ZgxzqveBmk6ywrTman8eQi6SV2xtD1/cI37vDVLF78n+rxIrTrfwivaLLp1VHosF
se9gpYUPQ4M4RmEk45vepdvmLr2jSrMPD1I/gY5CSUmjDBhbZwq/IQKWHmMGcuGl
NjI2lw1qjsNYxLy7Fxb67v3Ma+erAAGr+dZifccXu1c7DLcloIrZNdm4b8BgHh21
ZyM7kCoRaaIw6cQsvU6cjpGMtkcL5SHG4sSB8FsSHmbEUVW3bPFhlxrHjHqsREm7
PHMg2RaxWyoL9FMmQD63AYTxMJD4mHTVeY25b6ln/RfTTQaOS3S59mIJcKQZzRAh
fXrna8Q2Yia083yVk+D3m0KnzCxXHq/6HyV3daLSNKAyj7cZKZBwBwbu6kdBwqeE
uDxu04R7M66l2pX6eFi0k4VmgSHh7vUtsF/PU4yoedY8jA1hNU+b63oQeKLg4hJO
+3qyoPlHp7Obi7BnIHourqn+cz31qka44xc5wjc3nHAOf9tCGPMml66A1RByYG2d
SRGw2mkA1HPhjNMJFyLZoQ21OPkMwwVJPd4NUL1e2JKv8ud/ndWPzcVAD/r6bPZr
2x1/hq/mzREAR4pSqG9PZxCWCxnzIt1C4rUR4vxBU0iyJ8kGtjvudCJcjtzNDGF+
DdCfYnI4DdKMN7rb5ZFm3WzriuW89TOaHUoNVX6mXj+CUVfkQHhRTzt/1cBWnnCC
d72FnLeTWSoroGdYf2GGaRjBwdxSlPAtMrOKHGI35w9BTFIBAkLBE7q+bSNuiewC
961rw3hiJQHR6KBkSpENM74pBu879aSyYQpV+aqUzWZxWRuZdnNZ75Fa7relhDO9
b4W5u+0JO5ePMFd3XdOD8T8a+dogBaP+RL2IX1jcAEC8lsMOcX9soneIEZ5qq3VH
S0DRGKlf2nZNx/Y7gyEAXbrmPWe32lBFGnPFtYKfHWX8cKhocwDJR3nF2A1ifN/I
JA0IC+m9Z7egiv2MlEoaGzGaiuVc8bcxROnZA9p0v9Yxgm7cVJaFyssEUprh3yJy
mZPNUW65BgJ+3bGdntA+SWi1Praumx+fOCx6qltCKxYNqBSnM1n0s0tvm7+2vffB
HoWZq4D0oMDsLCyL6apRT3XXiMKdOH1avMq0r2KgMwUhtrwjxzYGyGuShRqLftno
xsUCCba/NMUup9chrfOpJ7IJkiG/5SH81wmy7+MlME+BPKr6O8/cFqmx3ZYOIPNf
1N+YaWduk9mjfQbk6ELjqncNz1LvZ0K1w6onbTWPYJ0FVP0EKT9dV9Qt0Yt3Goq1
wToUV9T/AQVHUOY6CyXLkMOhh4veyqBxfaMwUucbU/OO9J2aLqXBnVixA8tVqLFS
XiBJkAlX4VxsXdoyS3uxG/JcqduPh7Ou1mq87U0JkDqg6PTAEzpzonwWB+BSn6Ga
cMu+ilrd9niBaoq76tIQ3Uac84xH4eIk5PReDkrOVJgM09LVrb0zvauxzzfjpjT/
jeUP051J3ukRSpr6M+5DYFvRz9ZwICKphSD7/EuByS2tnboBNAQzxVaoNFs6vm2C
rcFK25dRv4Wli2yhQUp7U3DVguGK+XYIlMdvW8PaSasEOJlvqYkFdEAsv8OOdPVo
F8uzWoff+RPZDfK1efTEqVDpvKk3gFfmu0tICT76L0S+1+1+tMllAOR4krtjq+fG
5pn8w86pGFl3AI9W2/Q2K7y857CyozJEW3c/4BU93wXFH2LkY2pzNIcQOQJ2C/ie
45FGUWBy2symYTJtwOK5tujI/FvRhbHd21hxalI8i3Qc6Q004cU12PIwxxaJUsip
UdayGUplLFJg5ZRQqBng3SRNFe1EgEKZ2+SUGaB7bJy0Y8vyRF1UFLXp3eC1CygG
E4OSsHCJafm9fC8NWTeitnxlnaTl1NlrX57XCItujl8SeSS/lwLtcnp+bC0Rpu/h
syUR3nnpmtCdmeaBz4AYEcAU1W4thSGugfho+w5jVRMlv51V1fGkEeVRQ+9Nt43c
kOD357k1tObfY/wxHnYJQlghLfWhjnFRT2HPdCG2dVnLdOQJ4AQKjUoPeL/ixJpa
GnY1Bt9MCDGmLYWK9l+e7DGYWjp4I26jFYY2UJqTLJcnCD4KABFfaBZ7p4Fyezk5
tmF8XTcPSdvhs/XRaqOBj/CVZQpsJPVG35agTlsRDvYgedONsrbUMNLOYYTqzWir
Ev2gD0SbR7suLVoeOQbIz0gZ7zxtjM2I5MNkuoOEx/MOJpbIQowg/hir5529jsN9
+iKSSKo+D+lNbaLImOrLkzRvfeD2ruRZYz/WXgJR3K0L0fYkj/ZXhYZhG74yXOqs
MUgt39YLziwNbWeBrB1teiHakECo0fI/APXAb7sd8Gm5m5XUMV0/8q7jUzp+LGRR
yPZDVR0lcqF2gigGjzybsoqMhi7l2WDgn+LIUm0BKvAeNIdZ4szkB98isp6M580M
919ds42bL5J3rwz7lXTb/ZaV1fSxcNrkW3wDBzSmjz/QNw7CBMZZxst9JyMn030l
3PlTjY52Dse/4ng0eJqSp88oKLbHt4w71V8YNmzFiaHhs/mtzfBm+N7ZK4Z46B9v
nW5teHmlYmBWupj4c3EwuucjEskOLKVgyCSVJKW6JOchwYt9gfhOK8eHM8OKSWo0
AgUl5xhDBzGhrI2RxReZ/pZHbbxIW9Xdt7KioTU04L3na90lDO56sax9BULO8R/3
gEKcmh3iW4BCinUtoD7QhbdFt5HqZHmNCZehldowPAbzcStZyHeM5pdVH+qIpp6Q
s3j+3bnn4HWbQ6ZiaNXAaicM4My83fxa1/Gw6iJq+e4i5lLH8vDEBbK4M9TcLzvJ
l9rMHKluxOCmWmbGTpPBJvLywGzTzbRcM+Y/YJpTNSM2GSWrmYbBmRqpHIeQIGOr
8swPIuNgeFo4du5FFbQX34GS0o87rlTdZY3lDkNjo4SnYE6vXjJZyx/J6D6FPkHw
xH5mfOO6ke9cPOku27CZH2jBZb3K1bAzz2xc05CTeieQqFuNUbggBDgO1QejLF6t
SPsY/vs+Th8xJjxlFERddM1w+R8ohmzVwXkGTPGi0LFKXfX0WBnOPN7HvsDHmvno
RJMjgVJs6QXXgk4cBrB6HCrJJmU1BcB4e8zS6AHk7Cozy6AJMvpHLkiO9tBj+xOs
XK+9yiDEwsRPRlIjhe7cLKqz5nOGhPgwTmosNt6CKN4gbngK8wxVInYWrFlcLh2Y
BEVAXbr+yU6uPfa6vLCIFgJYJaSz+VUpCEXX2ect4lqbXy5Ae9XZxcc38YeMrh75
BHTws/XM2pzQK765sPygflpRhC7a1rq8gR0hZjgVCzk+Bofii4sfLIHP8atDK2FP
EOx6gKBqqdSXrOHHhYqA6f0WD7GZsevqf3M4dpBoIRJlNbzMEv4iPQlJJ4KRH9mh
6M3YX+12VBR3/zNhh3DrHPD/iCfPMG42UoJ1dkaeI148xI88Kkh0LaWY6zJxn8Ao
KmJiEpCBjMvBIXW8w5Q1FyN1dfbrGtZP/K+dkioi47f6kKs/ElXqkd4r5onpvLJf
eEpaWWN+5n16JgLs6JCW7VkKej/4UwjV95XBTQk58awMypSO1mPvfmBV3/HQ3V0N
tW9H9/yK1URUMvTgaqRgGRNGSZdN4Hl09Ic4QhqmQV++N7xk60UjP3K4tn7h2BYM
TnC17SIyW/b/GmfmTnYAimJlHXnoH5BAgssf+8dlyS/fn8YwZNXleT3nHGceqF9j
XPyDC/UsfmgoPegez431SAdRycdrdHqU1ryYSCPB/xOY/1Azq/foaKjmDy5VuNvh
8d3mpPNsvWTuEPKdjnNeErJfiH3P2kduv+OKdDxHkNkOc6V5HYcEyEcgIHyUUoIp
xaDLYOLoum9RsnE9FgKQZMe7EV2kGxDjulaC8NKfQzzXAzlpYL3pAGmv9QmYWjcP
gSZfrA7lOazD3HoJu+iQQeuZr0olVp5E79K4Tqg8J2MRapm1xeJ5i+Aekbjpjy93
0gFx7bqvyFM1vQT+gztF+41xDeUa75ARsyWyPlISqbiVSwJYgI6DXkqBXUG1WBkI
9wNheiVY9gTn599L6Q/L89+EkleBuxUrS6m6JWwu5U9tboVtfItuxGVfXJcELGL0
6vDoyHm4pJZy84kqaxe2QpjnvaMzvUWg+5IdNgGThyMzbO/jBw8j2NFtlsGRLW3t
YIWhHD39zRTGBktELaoo2/NGMJ4jM0+nc0byGpwlCeOF+5DytqEzzGpRwGW7mYVO
706Gj/7niP0uMn4sg/p4k/PXm53F0PAr41aqa0zppmERhiDqnBaWCgLqzvPo9P9V
e5Cu0R55pnL7uANak6BsqXmA41Z26Blan+xEJs9qmDUJ9rzdej+rDMgoBrMNVZ6M
Eh07ysOvg1RZPJlVODJxIK2BpjQ27RsX3UUN9Xp6Ur0Fv9uHs2rYS/YB7CjavaWg
xCXvjcjE+HWZAnYQ7QPbgBr0XGm3TaHeL7po6T07yOCGqHrqWQIhwEm+waIlxBHy
oUI6VwyTXdPXy4HyYhygv7gmITQpefK+YsvSOhyxfSsxC3ZNE81oaYTKEcdaCI5A
+AIaNVS91Uh8g+bOzO2HW4/s9tOzcYlENqOOkoPgcEUuwkQhrIz5qYVF/I1jVe9M
YXJzb8atusjSImrXDZIlr9A2Z6Ov6X6qsw3g03wZOqlbGic5K0dftT1qdUDI7rDp
rESCW0CkSY+tN41RM/8yFYx+0onDLu4NAy/bhkyVYOQgesOjLp4wH0K7WLBnGWgE
+b6/yz/oYwd9Zut5hv60uHg4ZkIFW/bPRU/eTZXcaovrg5lKIDEvitLED3HGkdxH
GFgHh9y3JPFomynTRG/dAdu/8ldIxX0zBrFduufUtYnWTeouEaUX+TMFtVzf30D5
U4BgATy92ysCswGdA32Ti00kjaobxKt+L8iVPQEBdcSV0HVp4q2IlLdOj7WpHgTv
phG0GeN3CXQH16UfiX2JQVv+Zxw3akmy2adzq7UI4mKR4D9wIgc32nYMWebuvAkA
DpiUSxnit6XM2YiIHBKMTqaohF20CWgdDOhx9ZhWUF0UDOWjUiCEIQKDH2UfL2Rt
7pebFpH9k/na860p2+XUNRP3PsR2Nbc7O2pkwOi8OJBy49HSw1vqDMkXkNA0lPRf
cAPUf9TeBg8ZRzhideO1GsCG/7t9al2kx193tulcMLZGbWbZHgJbeeQMFB8V3vQh
nDLpUnbB4Ydp8mEdyhXyQJjsn3jya4LrRx01BaxRnLqXfLnVGKSbFEcxryq6L/RX
5irgUerdOmstAd2YYcSa7Y5Dh0pq7tNQ8nLLHGrCMiiIp96iS2Q1fMoMRAzr+p2g
QIGcR5Arl7v1C5CNzkynruT740ZXLNjfllc9oRPiUKD1IoPp+WQwkWk15b2YGMQf
gEFHcgZn6wvFzmsd/SMvLXpMa7C+7XL1bGTl9smr8aUcnrNJySP9U5154cTB0Jna
UyL9vApqnx1zn02tsBC+53vW04hYLTMkQTXyMTLbFdIVNDw89c0YBrBKyq7H6L9J
kpeSG/m98c04GSyIZm2QiSaLkRISH3/tiG59tHzrGTdZ+hoLMLlwFecRcQ+r8tjn
xnRizlpmHZuotkfLOs5D56okj31nfbLrX+oyMVdv0MiLH07zQ2Qi/dsb8VdK+5j9
KHWrPcqAnuRIYujJ42BU6oMMovNNUNX6/C+sz5snyZbxbd5DtV5D3F4wIhi2vMdf
oWd6PKfa5Ry2Fcs93ahNB1iQm2bskpKY8klbRyHH6CEKeYifyKyNLONfuCGzeWzp
OjrqkJD2dqwSmB6GrTXotAiH/St4NmQ2ehI8S7lFKLuzZRyhOyOsT6k1zVkdP2fr
yWobakYgBXZWBK/FsEhbvmHoHdRjHCa8JNSAahHM+QANgtlDOA6J+oRTq/zo4u37
7fARs7z2kE2jXBbiOynQX5L/uUBzQ8vZkAkECKg2s12XIn54jqWEO5v81IqmVFvo
JCMVnDLB8xWwoQKDRW2eZDjQaZ7DLm3WSFjbDoiu2lvYvnk94IC/FZSfobJyN2FW
k8LWO6Vsb9iXHm0P+2ScaF3tS8x5IGRxbrufbiWn7EJbDkzbwd0ej0nsyY1b280+
2QXwvG+NCnpw5NpXRHfsaNjMpfHHoEJjY5K6SZGHaYY1PW5+4f4djNsUqdKByv7e
2h5OVGdVCBoFtLjItQjzNg9+ET3FFporUOuDPcPw1EA66bhzc4+CNprF80l+q4dX
IiZdXAlN4+2FxyUhPpphw4ZwpFIfuNvHoFDsSaRjpyUmCqyylCxDSonBsnKboRZT
AO1+WxnIDiFgmsWoJCBMvHcaGgKmnfH8BstIVw3/toWHgFOk4v0cr6GzeXB9t83v
az4xRJ/IQAIReXk7QAHIQ7hnEuRYBh6k9sTXIjgPiSLXAl6M1233JgVPzY8L4Xxo
k4Kv22Y6e92+RPJGElO8LWHBQotOodT4sICB4nHtTYcMHw3uZr9RO3zhEh7vXY3l
BDt2ZxSOnGXhijhLKwBVXx0l53Atf5i4NhANwVY4FAE1LZydJD84hTu3oMYb3JOr
fZNUGbbc1IJ91z4b50ESnGLlDQkLvlfDQ7REd33M04AZJYGuTDfAefhncs/j/TVa
XpWRrU4bzVl5VIrZWCr+0FUmaWKCMoYeBbadNR3/FiO9JZPqeFAJcPc0wOVdxQNO
eRdngvlsSh4LSuaZOcfkz9XA3TBOjmynAgQd09MBdTQN3Rl2zYi0HlS9XzApB87N
MOLi9Yet9x8y1Xw6pX3qkwD7GLbqM2zrkZAzbgTR/ctNp27iGDMHJRnUu6SBNhaL
KqztiB+vCgyqD9G3nid1ZxORiP8gwHp6g7Ba8jhipy1FJnsKUuo8q1vTu6UIrdxB
1Jz0q3pQA7h54DFxoYaU+ED/ea6BfpwhgkZENY+4eflcK1KIWVtIhlPWIRUNzsbU
ar0fVGLhwxCcbOq4HvM41+2qgQQV0CUk5idWik1MWfA8CKvxf+ce7IEMWeeEaE38
mG3cQXx7TV6EHDR5BDQ/50mYrDdwpo9m8lbZszZAN31Dx1KOnQ4tH9KjEJKH2LAZ
oKs35C+pkjGn0CyJyuv1+thct451MKlCD4oLVG5wHriqwMMw0nR6/OkAFaMJpGh7
DKMabj0ul9TFl1WdluQo969Evvo/nOVr+EeyeYbWCVMbWxtUwoABwwHc5AiI2Or7
dDSwRLrKeSIGbpMHZ8Yg9UOB6H2cu1EoXg8m1Cg0YBXs7entuqS93q4yRSPNozj8
e+iNnIRRw7JCHRMN6JuxRwKWCrtDQ4gR/asVAkzyIxQuyEDWH08RcMIQKBYyvOY1
ASmhBZlTQjAGLwvKT/JXBc5MOhtC/PG7vPpX8sNROH7irrAKKkUDU/8pRQzdpl32
IAX09N9pDfv0aCSI3KIv0gNrAp9KyGqqNYGh+DBvpLlBOQg3SNawUGv3dN+ZAhmC
ovR9g8nuZHQyN7/KCBz1nK6uIlS9ucxzlyoQgTKL3ZF1d816uB/yb3cDCB+V46lj
TCv8FbYEmT4mDN/BqeSZY9EhZ8JCXuRShTp8Q8+dfEvcgWJt/SZsdMGRT/awtmnA
ERdW3HS+SnUUEneJ/ChUFZ63CXAeHvrVsELPZGDYc/feYBSk7kS0dfms3tlmD2ic
+Q6sr90+Hc4FKL1IvuinVkXQF5T0JhEdUiikqXQI0h2GcNrfpiLmtFzY9IaoWLk0
69kKyzbazXaWk34BeNpNqtLrbN+KUDGigv0DGiWHQLsqcjxH1ZWKvBdALJO3QYsO
a4/GHmca8DP4baT0wHVQ8LCPT14tTPJgK2I+q96cavJ649m13FI2n41XA8eEgP0G
rBOEBqtcqn0VibtDaXYdRGreaVCPuEMEWJ13MLpHrKXRwdizYdI4jM70hJd2mP6F
ZMOAa5NdqbhCioQeLBIZe/KegS2LPynxzePWfxKW1aU99J/46hhVz5XqWp17s4o6
l0CUT7rBFIudNqWLRkp4YY5E73Vv7/LCk72wX1xIt2/wSdpLrErelJeUnpjdYwxS
xHH4YLTEr/an25Wq5odlTmZf2NqZlk0FOmQk+f/k/BGId1N6bwF3Zuo9n+AEQIQs
Lw2kB8hcN7eGKoFDybQKzaMuYTsyNl0rjOnY61VkDwTlu2Dc8OVJSrUpRXY/3WLo
GTngT+IqhpCjZR0njsSzD78mqx8S6i2lMHwT3PiZc13+sAXvKAOYsPoMLXavmlpq
5+x/kyQ5oiO7K3AWIVAPnRr7DUqw8BZARMFW8CxcTVQqTiy87Qwhvnb1uiwSEOFe
VMZnRglg9HAdFvvxBEOXXFRVYcY7F2/bihGsVj2mg6wT2oXexOiiRy1EucKobQyI
BWNmO90VOQ3UaGEXzANtETCbbE61/HYapduBhpISnq8yu3JBlWo9r4lK/KthwFsO
6FzzxX7UfxIy96m435j/b/eksLn1Hi+8jU5tODxgBxV6XH3AHFBbjkH8pp7/m/mW
K/DzWqwP/ecJId1kc65cDkn07UWgSwgmyzh1pFccTieoKNvN02IZBsViZ9mkDkGw
MWxsK4HlNcAcu9R+v9amX22Nyq7IvERs1sI4BzZtlIux721aCNNwAjvfEDOmqOIi
hEoZSHXUgcqBziWWpxoaWuCYr1jkIx+QVQ7mDsGCfoNfMzicNLJ5dWuajydOu23T
4yFygF67eYtjB2A/lmU6xJ22dvOdrRVnXdbQbtv2kQiL/8XberR+9WO/mgZvudyz
cApyO9aG334aw+uqCXnC2AJcXSNQCvtTlvLu4aIhFMSkxW14kpoVKdwn5Og9QZCU
7YOHUEp/E92cGapalqWKkjdBnb/ha5jB2IxtLJgbIij58cyPOVwT35kv5yf82gCd
7g3aI3SXDuDPKJPPX4GppnUqMLa6GBO33xmLufxlWlQ1CCzF+nJz/6jazutUuPqn
vtJ/kvTMO1he5nAVZrw5mu26ZMA5LzlA72oQDpdL1bOO20+zuSj5GBkquvPGwnG0
8VgAdsF08ANnRIxao812rkdG3JIglxaF8oJFrBul1P+S1HaR8t/txdeP0/P0x6iM
zLbPYgVVATctklRf4lvqkHQFjArsBcmE7jGop+mxEEa7eIFAT6Edwt5HvupY9GsY
cOTVp2f6q8kWt0X/G2mfhb5jYWylndKLCOXl+MM1R/9wmBNEO9vqwIsOAdQl/27h
8OyDq2tMFf+4znApiebFXJfKsRmz/EtgiUy41Iuh9k6JVxu9959SwxFfSi86lzc0
cUwYaJ4tCivJGSC44lU9zz0XTQlQDbLCPVSPppn7VRZ2J1G01ODI8AEWZ5HXn0It
HMLnMd6qNLXN8vj/xI4aTFbUwD3fWRqJeEV+WXHRLaaqlGgWWAY9Mb+wpcUUpAJj
mrfbJUEHnmrWyWAOymWTaRDLOnlrSj/XJv0UWDXnA3IeGsrXJ8DI11btnGnM5hdj
V0s0WgXRkm+fbM3LeaGuoW8eCZsp1iPTtnAKMPpOfcquAHUH7/Z+4RzPjkXbtj8a
8bxhDQw4nsTZLhwgSBDZMPi/dlsCnKToPhRzuq0o7ZFxNT8kaMCMOlkrcllti0rZ
j4D5jBLm6cNt4usYCvFiUP64v0rAUkpVV7+HPnk4WRFNC0En1F6frngthQpXjUOa
w074dxTDjMxa5K/DysaonsqcZWSIoQg/tKi6lIXBEvpvUxajbXTvI5qTjuQaUyJQ
4UPC900LL9WCS8qy1Y9OmgtiZLSHfhx4AZs9UseU7Z9crsrmiqHsHE013dsMohHA
jMZzq7nhVerveisCDVXTUD1obgkEWC9VSpInyrux90oNawr+pIt1F37n/+MFIFlz
pJNJDzcMiRlZZsKU3cBotTDKi91F7fLGA4uyhJ8wHpXhwTtC4ZvI+L4bFCuTibQY
w6C2oXIEEx7OIacxEELj9Wgwez0okXXzIY/5pH8lUwPFGEPbSGPaPeb96ThEl2XZ
ztJG53sAmp9sgZOGYMKevLvBi8IJMZFuLJ7TUUnD+401EjHjobSYL7xCBRmVfIIW
bNJJpJJ+6DA9g/lEKXoRJQs1tQL/iWUEM8d2I5odUt5w+8CTuUaUiamVkiKLXVX2
tb57j5DjHamLswovOCW02uIpyNFM70f+XBCeFoIGqTaZZ1msS9ToW5i5XRtFzRa4
PDfeXwXhOji+Q2HnpNQA3sU68Phqo4GaYd6NB6q88W8Z4Bi0HwSgO7rZUQlg/7rc
/341GbxmVDkh8QNlSrJ0MXwFVNrOe+/AZ1Y/QSzhY96+RnSrqz1uCjV5J8FSnzXC
SKMSHBbxGevU9y1D9tdLBrqPQwBBsAYo5v5q5cfXjbYctQb+dtrXWKNtaQVMhhtH
0f0Gu174W1IVSBliu7PW49ffUuXFCln6YCYLhmHvgcdS8j6rNp1P9Ie8lh3JVgpI
DeWNeXTleJPMJfa9dyYRlAsOUUM0MVsm85JjORhBg2Jct0NK5LYi9qx2VnvX/I2q
lD6PqBmNtadnbPzMWicJTmQ0Tsu6KjD+B6LXalmZjogwN7gNBWC9LP09pBQ7pQO8
IPyuHywv5l9m23jO5HqlElNuHDho2jbuVk4rwgHd6ol6EM4kjHCDgfsNBRsgWfjG
/3rR9UvSAdU/QAYJ0NsxcnCr/1w8/J9D7PcAqMUo2s6e/Ju2hdNrzX/+zg42RqSI
HVkdVTeag8dwKx19g3axqFd/RYPew6jL2VLiNuSeZqCMjXeyG6RapN3ridgePM/u
VHXR3e1kSCBddNj+qIgGj4A3O6kEWx2XsEntGxiO+wBZFsHAEUxN4Vc73rEaCtDK
UrZcX0ZLMYpoyBny586C031FFjuXUA/THPKnTbxxSC0qXOsZ0lv17ekC0/CEz8x1
tqXmG0DMmokG/u5wZA4UQD6CN/sCTlsnfPT3bxl7u2sDVnxAkuzmNJ7QSBe1n3N9
HuHuc1aREqGh01hgKtKqOYbsgEqhE895+0OeDFpYR4TH9B5LOtbN6Kn6UuCLRZzE
0p5stMa0p0kWEbxLsF5Ikf1wXRK/S12X/vcizJUzEKMFKBerRk57d79YQbDT8sLd
wLY4qYGf5CCidS2wAz0Cc4MDhJRmnIshNlVSs5MtYCTpR6z4iGZyDkianMvQvtje
r3mJPKgzGdSmuD9yF1FWm4Jz9V6ERcFTtHtWfWpS4AMbVinsn2Sp18Y5me3qcttY
R/Q78AruU6ksiwiWg4Nsj6Q3manZnRNM4TynjvfcFGWzUwbU57yA+91ENpqYlYNF
ZXwWnXXqDAr3qqnWM6TD4xuExI/s8MWdZ8Q9yZAmvXPDoaN2rUibaADK9O081j7V
3VMNFbosrxKElL62691hKi4MpadBIL2jVx5Jnuf+6EWchYVmODS2+fgKKIMJAJlk
01Rp088/bdqh4SvygPHwW1SPGUrzz+aECgdiQwhSct+Xla+rAd7V1EY6Op6p4n2r
KSN2RQLh8Ed1KtAzCWz8jtEktq7C9qiurv0OzG8dVK51GVPDHy5wopZpoUP3uuZg
QKWOyh8krkH+G6wtKFHFXdb1Ouz2vPx6rC1HbDB0oef3KoObHOfComKq+6ti1QR1
RCaRS/xT3gdvXi/H4FTzwQAmqndsLz8pT8ktYWm22RwDwyCSE3BI/ViOMkYkUMkY
5aeP+EJUx8iuPEaRhfpMY9nLn8JE+LgM5NzAPBoiW5U0jTiF3qhZz/TOJeg8aeeL
x+8MEhFRSOpIZKJErmGNDuoC/BZCBmgwM4npVrOtQrpHG/InjkIpPQYc2KQMnLhv
UttTIX6T7i5TdKtHMCWA77QTBsknQr9918nusLRcB6Npy4zXf0DTElwh/kjCd7wl
fRDeSvdplKbhfLn6Lwd36GbImSIWSjOJvluSdOdz7RqhyDV/STCuq2apk/s/DLGP
FbWVEce8QbaSpVy7FufqoCqQNrFsdJLQjQcWx/vi7kXb/Z/pLYAqNdAjJ+zgksOo
Bk020/TtIZyMhINtKOPhQoo/UoeXWW+aQ6CAbZPbzVBI8AjCr+OAr6FT/3Va9djM
BAXV4u5NQ779T2P+xRHcokRLz8b7RmTBA3LBoU8tE/MqX4b9HSpC84pDG97tknue
fLYDBpalqv4SjZ1O/AYFFNxLyMcEEQ0I1hthe5ca1/Vu+ciDkXQAQTETgcnsg8B3
wFGx+DnERSpnXncx5s8x3jnMJURPlOUp/TLvOv/dkqSud8JQWPClJEpV3+MjFvVl
pkSSwUvBQGVZPfsoWA6L5/GHiiRHCDy5CFkTXnD+hWviZaZgNzKC1BjwtjBuHqNZ
rVAmbXeBJLklsiN2d//UiIB13S5Qhkdm9bWXkS5c21r1Y0SgcjFSMks6rBMvAjXb
zsekPFv/V1TeSj6c5He81efRsVVz8ISn8N5CRBKuM/ijBTf7zJa9uvLo6pzMWSpY
4wNsAz3B7fFxqYYJGhbPSWtk9bVhw6Ugr0NtV195QETue/T2P9JtSjoZrsB/mKX1
o0wYb6lyPu+gEvR8Ua4AiA7CfDgV7a4/ywHyoHqXHLdnmVsEZ5JpNq7qFPkiZHst
uPQ0am6m9QR34bRVD5JZq5lkPzZb8ymIG9Vow75hNhlSl26Z8KQafsovsPphEh5+
aKnQDVMOUm8IlFkM9Npezel+ebyt9CZXqUfhJVgq/CYxi7qAtUPDEgFzqOl0EB5r
171ySppcR26fAdP8AWhoAqr/0d1ntO/6Ke14K1uU+onZJsyFVwAnb0VumsunIqFe
ti+usTBRZb7AHJo17by++6jxAu8uBK+Mo5j+1HECFns+Z9e/cEOHHE5uMTMK/apk
n8WmhOwOxLpvCGjvR9tj/txK7SwNtum1jvmZQ8e5Sxo6o1ygcEtvA8myM27FV1mF
toOnFAYTxJR51VZAPHEqoAUaq0lTPHO7virF1i0gKC2Ju1b4zbURUjUkLreQy/RA
XrA/itvc3zJ3tTqZI9XlCDk7X/mMGKflLY054NJtTr2l+ew3JWXb6vq3O2eSsSu9
T3eI9V93Xcbi6DkaZGcbLTrher5bxak5uBLBEZ/7UOTL54M+/8Dd0Y5LWYPWlyDz
dBY6y/B08jc6d/45x3xLgvVyosUq/3lhI7RER+HnrJa4GC5flmFLY5BJ+uL2S+oK
6PBfJHY1X02g/XUY4zqLm6yC3ZM15aSom+/EPOnPQbwyrK5t2+3ij69POFu6SDS+
wY0Hm3D8zQ9+3d0wsPTEqSk6ejYT3g0KJvnJqIELsXCcsy4XkZ8YNSZep3TwznP+
Heqi0Ls72+I+X72csLuXj7BielWtSYZ0ak5wuTvyd76O75pOM3nPxSbYUPQhO2U1
6KlzuznE7DznVVtHiqn1kdbciFE9yTgwowfE6DCabD18PJr5tcTogd9xabJsd/iu
ual4X4e9SXUESocndzppxauYRjPjPOgbXi/qlp9Cy9PKoX5TZVfyLNuKt/vTxfde
ywaCQnJnyQd4dr5YG8EPF6Zn5lO+n3PVR+ypq01waDt5ea1OIKvpTtF7/lR3+yJ+
nfcgncdrWQ3O05a/OW0ojD5anbt8Pc83OcQfZL7X4O2BWVzj9khLaaA6MpRN7kOh
/rQC+ZF259CD0tPn+MPmqSL+hiMp4J/XVG9WY30eI2KDwlqWQwQEPkkBA1ZkCF/t
qH8LcKpnezPXWArd7FIigUjWFp8ZbiafRd8JbjdzRuv9NPzdncB/z1JnwX1zf0zj
fv9W8mpcpvqqXbhp8wAn+Pq7Hd2EqqmQyrdVb5bSP2nr0EGYiWinM11OAcwT8wR4
PWcntj2xZF4RGogqVucoQLduz6EZ49u2QuW3lEc5ZQhFjmhRP610nSxR1MgXAboy
d+djHdFYpUh4MXQYN/7AF9C9/jGfNVk1cmFkq2MHWLCkVUJbTUqXAnW2cJcy+2iJ
tjLxsDdm3/mV/H+sS08rqIIgbQkewWUNy4hIeSg4OTdGHmSfC/FKIEWiXLQ611H1
pcSZSg4AQ8RDtlbu2KdOsTL7fvuHEEi68/2NxshrHmm3Bbg/OL0QtXe0neuPW9By
D/BdeXpswxR702xtSwyQ2Q5dglRyc8vGf9yW6vJd10lugHYGA3XmHXnnbt7xLtol
QAsXEmJ1APCEdrDSo2DJdrGdYMwkJ88avNwnDUqKg3OIuzPfbBvAO2oKMSUJQRQr
Nl08mmmZmxUmaDTGtWNlf7lnnRdVYcpIiiuysLeKuKlHPE4qgUSZjydBLUleQCvv
USn/zt9Vq00yXIzYDb9ZMmS1FzGvzrxdMk+E6qMaAkJt/9EAuuIEeRwe4AEkAeMk
02GzsyMJBVKgfdRnkQOpTbVu1CBqSzMiSmaMUZFPNqWllSNa09ZXjV0lem0gY8SU
iXm3aVMBv0msOTplbF+Tbrdz6oHWTcNOemjAXkTv2an6PGvRZmO2kePN034KY/bi
YXQGypCQqCLcogG4pm4B/FDwJ8GlHi4WDGlfhnwQYk01mvZava5eW5i/ZnEQWljl
AG1TBmmyBq1hIiw57zeo+u2ammEYDrK1sluNe6n+SfyeQq5J0hQji1Bjp8Gk3OKy
quaYN21AArhcpPPXtwHGjmwoBRa/jPN92gVsLBTc740/noWBxCKeP657aexdTIip
pUJPHyROv8QIutf8k07RNQWstG/D2oVod2KHb6OnHBaKoGZgGl4l3S/OafBQ8c7Z
C5wTTX+Js7Ob9+clMWF9d4OWlgiUhac86E3fKEb4fsiFGXCf4kzRl55XjOj/Fb2D
7grfTU1rXkxcaEm/F/bhwP1pZHaOc8v7yyyNsyAheyMKk6HBXejAXWikSkEG1LtW
LlLTcR6jYc4v5EwvaoPupmrZCRAkB9pJtdoba3OrdO7xel7abhACsz0bg3Fj20Tx
yegEeZ1hRBGvlli+8zXUsSrE/4A5rdLRfRPXhu9w3b2IMVTmg7W0RI0ZJ1P6VEil
o6WlUXh64DTqoGK5WHrgFwQ21Hvjjo8M85sNWraVxfYvurnkI8X/fbSMFgIYchVJ
zI/MAynR3aPPLVa4DTreGFIUw+jPz2VgT6cqwddkuRbI5k90exAZ7Nu2RieOwi7f
U8Zg54lsBp9rtb3wZWz6y5rE1AXbGC/82tXbgbXUxdvez2u5J7XmVaAujJ6R/uwF
fx1fuMLVkiC6yovFoTqWWcssE5/c8H+4I+qtsUESC/JVLFR13WUERoCxbMyhXLks
5MbAUjUmak1+jhkr45knikuzBz0LqzMRHUXGWjCs5fWLERlkzJArWKPASQkU+SZo
EhhlsMItNAJOgItMeQSLqiAqCROmRSsd3mOzx0Yn2JDys/Uvwskn42tEHcoSjGMm
+RekEKD6zeIEJJg8AJIeC0GNQ3h652uIs25GPwLEW9iAlZYB92bLIKQqozQFvGjL
Wx6kWb+UO6Jl+HOx5rdSgKOA18xjdjDe8s3E8tH2zItzHv0uf6WNc8QUWqwDAWrB
8wtDehbrD/agRHnCdWWrYTnwaIWAJEMiGybfUqG4dZh8mwTv8xvoUVjZ7mgLXk39
kaeGAv3LFndApCk0DAATZyS6SQZMqPLkjBcUeVr2KEBLVIHW4LU2HiH9g9Hpw396
NguCvNywdfTdZxr+ppblL0UJ9Ntrergr3aE9FOY7CXouAn8B3yXDdbiqIKEVMVHV
OUL29bMFWDo8PpbScORLdDPZ1OUE0vO/zTz6aIcoRon4Bbkmd+Qxj2qCGH3x6Gio
Re/dLFS8GjHPORhCtm33Q0NMK6zl0nPVhkKNR1ACERyTIzhBui+bVB+2nyaC+ba7
U8/ni99K3j+XgieIiCGZD2230hV8e8a/bqq1n7gEka4MK+IU6Yp30uroNmeHA+gK
DfnpvbUPCkQhHhrf5mDWUDWO8Ag0EQ5Hl0+t7aH4KEhlLgbgLidXFRm37R1lZa6S
5/ozQy9y926mc1+xDf0/lEh28jsJkcklOEn+kplMcV7vWKkgudvO53ur4vLV0KO8
wIe1SVF7yimuwIKXwN9zlrUkbiiTt09AT3651NW+BHeeZoLWo7iRSZb7u96toact
6joHoUysE55LtI19xdOU5nO7/DfPGAp2U7gal90WsXwRI+yn6Ofss9iFJfrANT6m
Tk7wvc9ur8fVTJXMLxwEbQLEh0h6IyFbIADHSEc23hudEeG6wQ/SEeAIK1flgtwD
74RkYAZU5auAIn2cqumnUu6LO0CBfCXv3aZf8v5LFWH5nVqnuzhnTS5z6zjhpcqR
0f4Uo0WDtvwpiS9Mes5tj8WFJjyvPzPw16tb5JUnrE7bwg1RtSJyBf248Gq+4SP6
gdeKnzUW0S1Byx/CReHUCNbgi5X9P19sOgBNXavNLwOiWMEXOgLRjEakPiaZo3G5
Jj7X3th50VjaHcHC9xoH+5hbhXzNEcDD5jVT9qR1t4kWqYM27RC/I6Z9grvvhuB6
8cwJo73rqribOfZ1l+YhVS9j0efcYLNHHdB9NCCubhV4d7SQzPmytzNOmLM/wvJe
eaDxyOo8yo69s/0nBcyR4FeghCuT+uAYl+CN/huo2sCfhh9R9nSooaJ00VZj3hpq
cHYxowsWt1CpIpxkuat0+kd1xraQ5NE7KyUKjRdfHDfDRt/dq+KFtvR6cY1eERFx
W3ZKlzFLDhIIMoW5IVR6NJnmkoHjK2cFpmM2T5xkI4UG00hMO0qnQ9wqG/BZKoHL
VVc543loq/UoLI2XXyuwYoDsoWY/jWYsdllI+Yc+D+ZGXoe54yjz6AjIZ0fuBAHF
HLUGNiX8eZASq7cMKEuwn9ZHVpw5sDEbbMxDCTFqRLK9BlPhLwV8rSeGD8p85txa
hD9PhcrHa+YRdLT3B1U70IQCKKP3ppW9WZRo/FQvgFFJRAsMxTgB2a0szZw5LkLx
QqfuXQ4XlGWtxsW/50321/g8ybdiBnxRcNCDx3nPPIElDC8xWRNe4V/sXsXTD7/W
Zftfl0jBt3lglVDtLbEPA4B6It7yndjAssf7EPb13+Km6qeENY59OwTvaOkM2q34
EGJOY4w26bbnegrIjLTSVYwhv/DoiAjSkVmRE7XjO6vQnOOy57mKxtT0VS6QkqfP
AKPYczdQ0wqJYCti5KblkgtbQVcQ200+DsTMFAOpDFvmodDOVVcbCZEfc970ytvF
3F5NLm1XUZnxUXvh/vBjVObFeHUfHx8pjop+cO9VYCTnepSccRjqxrASWhkA0Bsn
8Z1dxGKHuUfXq11+dGXA7tbDXB4Ss5wC9vfF/2EDH7W5fTbCYDTGLUiGV0Fg6ysk
UHyw2HZUmct0L6Ld6nBzI8bhbHWH3NXEYgPecYvgCwB/iKzXKAAyFZB/SuFkVlwI
DT7XMKS2AEHc02vowd27127j2oZQlYleT9TUif4n6ISqbZ/JfBXWDysIDdivlP0A
EA53qwWeRKuiEgUJA06KKy6gotdCGrtHHJ8ZqORXRvINsrKCffaGMXkzNEnJc39g
/BEkBQgCfyKAq8+Hkh8IG44tY932tYzg0YgXWLm5YnYZtE0mO8H60iDM+Rbs4RIN
a69FGxWri3fWqYuJ9CPXQNfCj8+iY9wIqw/MvXCIMnp+JR/g3fZb4grpZQEK3tJD
WvoL2GyJC/uq3JlOJI8kfx7zCvO8zOETRPVnIuzLsdDCga6N84ywFYqH6iGptZA2
Zm6ePuqfY5ZwQBBTo+mB+RmoMjtyooCsDs+sU8UAv9thKRjS+DsUaNotmsEuWHYk
Q9GnRSABxkVajCTfEoP64EZ6mUzAfAaOOgSpLAzYmTlxM+w4Yze667D9o8dl2EnV
IdPS73dxV2bF4GKNYfqE0laCzAJtYGDCFiiILC9+UQKCVeIDCwnoR2mi6I0ymC9o
CallRAsqGFrg86KekQfTZISbMhfKDalEBji2eB2SdflYprREL45PHzXFhA7Apych
WViTMGjSI5PW7vr8S/FQia8Si6alv68cpkBWV9kURMn1PTkEMfnTP2jUWeoSQ5KN
y8QX08f48teN8rHt7/qj0e3n9nZ+inH56iSN/cm/kro8TRzXxFEBddrBU6oMmkI8
b2UU5QIbQHk2WSWDl7HRkH1LusWHpSQ2cfXpHthK82hbC7bnFx9c1ICnEK4DzB5X
xE6kBJcvLZkpXgt6jF6qOKzyV1Xm5I8dk0jHZsweh2n3Ke1BavQj1vo3yQFLeL5O
deTpkraahxHIUIqStEoIvaDjguy4HtTo1X67AtIK3Hz+z9Ozgr0XSsX1k2nXQ7h1
124NpzlMNEX4s49ay7MriTEa82KFCnAI7GzDRA8z6iu0Lm+bZeuFvSDmZk8eWo4R
4esbJ2wz8FOGD5qOlOGvpJjfQjsY61sBYUN4sPAkKDLa/X8bPOTrIDpBA92f6zul
56RsFOnDORn0ayX4fscIFAV8AIYLUtnkFjU+k4k+2mLwJksp2T3FXRpzotGcm/c1
OgGqsPpkJUa0IoUoOHyaEfhRItpBWxJTe4BckCWF4LiUqmdoS9rvvUSVHcHfQWX6
nkfzVjyebuwwhZP/HjtmnEenNbzxpMMjWldK8C5Oxt6pNNaKBGQWUDC4xc+X2i62
638qgoy+uhOcr4wSvWBCv3WllyD2w0rtVaexsLde/RflGJHVDh2DXAyq5DEkaMbg
9up+vfAZ3bJZlKjV/qk5hrnaL1qgjOvWVaY/nYY3KKR1lMCWhltDk5W5tPtyj/kD
8dXcASWdEIdiPcGakLKclm+UXUUeCTa+aIefctT6vbv2o25fKcolqfazvbX5Wv3B
aENFzFulDmV+iw09OO5Cpqhq8HFmAqodjFvGEOJ2LFEmYLh+nyr3KWNDIAy2pqZe
whsXBF1UCIFFnfmCSAlv+8HhwAf00GhAoJ2+70o98yC8lmfw13mpNNUwdIGZT/VK
VZS0PPruFB5IGSMKxYATUMWA3dQ/2jO/3+pwaXKrkZHzKQQHPELWh5tujM2zlyrz
rLdN4lGriHP04ReXpxr/iS+qwOFd2wuIdyBE9tcY+yPUSvFNmwD3qMDlX63qWhg6
P42exTltCoomgnL7OILZKMQwC0IRWEO2OwfhqnIKGqEwDanmFkaTm5D7Th4Uku00
hwhCDBWx2H0TzWVECtPXRIZ2PkXRYxrkEUgTbYGkn/PDkvdulMuKC+OaI94fqZcL
M3HUpm/xvLQgd/NG+lW291cMyiQXq02I21tVwCFwzhy7y9Kj3iWjNKly9r0tw+do
pu9aKbsXqVWL5yZwf7XmlwXtjUbhf5sE9WmZKzpT6yRkjKxnykIRz/IAXKuE7dSP
ACfYWPJqfZRsl44IWBIcN3PgJajXrS2fy1NzHguuANuyXOduc3v+AgwsU9whZeNi
72WN2KDH5HPuo3mGJQ10T+rvM19WZReoMU2dilfXA7j2+F+HTlyHkjowi0XpklXK
cT01zCbvhseNAYIr1CGZ2mn44n1LHYfztfQ20qhk9MYbY/hD6S1BNGmGM5PcDKmI
P1CwoMXgpR0EFh1ekPWW74tdcdAnx0A4ljd+i2z6cGyfK8/qPXK/Sx+FsoFM2MYb
Ws5jnyALWidbFWeRB0eMJWutkMIOUz6GNj9aeXjBnrXB2W5mU2zKjcRkaSY7DjHs
wPRkacm4jLndjoxMPnXe4RT4Lw2TsBABbWzO0889JLqZ6rnYm/Kz8OCnCnkAtkgH
f7JuybdRCGVbjg0UY4bTVHTJketjcibCp3IeMeyuJiXf90zHcyZrCODPzE5J4qiQ
uQX1jnRFh+BJk3FkikRQf89/Nk7z4PumJ2nI1NLp8u8puQ/Le5Ulnxurs/AXkahb
I3Xr43Ijp4YFmaL3zAqySQ3yyybEQHt2I6WR+ZQJgFKOiouUCkytiAaFIbj6IGGW
CRZv1RlRRi0G+FyAhHEB6ZUwzQ++YcE1KNNKTqp9W/lPvFd+D19OuHZnsEWrByOn
kZewUZNU0LRNQg8PZs8menjgZw2Jezq2JDspuGEO9HjxueDMOcETBcxMxc720IDp
cDy8yz0Nwo2kLIXCl2daCDxaJmHd3GA5sV4aQCE7ZOYrknsdW4zjn+dqoOQ9OC10
Duos7UB+Rxh0puS170KvWVCm4DCou11KZ38NeoKLuMEV9Y77jAQUmOUDU5DCgPh2
R64L7o5alqtYqCKX2uj4sUljxJq8v2CXF7Kjy/bwT9kam1L7H55h6wxEXnsFSmaQ
o7uYQLuSyCsN6RgmUNKf/LVmMajaEqjQN/2J3IuYp1hZF2yHNc/CREuCsNwV2wMq
vcgElRusGMK3HjmCjFnw4aGcFNZs12IT+p0B/iezpOrrc+hXU3ow98VIZaNenuOV
Cs+HGL8is9jEjpZRbBJ7hDFUob5RWAC/kodKCHEnQW49ZlFft2S5PZ6KDMtvvHeB
zrr2Xcn15q8Ebarz0x1TTzsUv8cPXiN6llhNxXRh/lRVMmGSuD7GoTic49KbaJ+W
UNbklTKvt/heF36MmeBpMnpuG3HiswUC7GUhDeYH7oRqF4SEH8yqF3HQGoRQICZ1
pNNLgIWncKF5Y1qs+gyWMNvRpaHIXk/RrgN2yjXjtC+7eJngjEEldPEh9ZkulTGP
FuWVREl6kiWiyhf4bmdpkCTuvsRDRZF5w/4kMmWXF73+eoiOFm6f0LKC/iOqD6Yo
VASpQxJ0QAbsBTiZX/1e82bmIwwmPCUVd4APWFCWfaIp4xdk9nQgzCV6zzWsIRR6
je/HZRO1KjJGho6Nx6B34+oQXbdN8z5q302mfgvb8iLVzb7R5mP8D7BCSwW5Nm/p
XEpqhbMKhrL2SFj4weePtcMsymsOmjfUtpauy02tgIIVOMNAFinqNgoviftM8Air
39F1k6bsZaXF9MNGyRRNJXVRLuv2kBH+50aLnbcRLPnPVWkTiMWcacl7/ijfpKQe
FbdG6bwZzJ5PTCeEtbAkMNa2z5PEQk+OwbOPF5GsAkHGBCU/pX8bkmgPWSr21NkI
3MPI494L/j7UlqLQksnFrrNX77slN7ZvxjSj7HfHwjjoBkmTlUqF2gP/Brpzi6qq
0+sD6+5Oau/3Qf9dwmM5NwNcJCRBfw7Mxo1+sCWziHODid6VqQaEUXziasg3YM6Y
gWv3QemNNyRvrClFKCYWqLY32sD6278SLez+M0FF5Eu8oj3pw+3mym91w2+PWi7w
Waod7Oeb8c8VLV1B6IvriK9eFH5/omF9tJhFJEIpC64538tO14eUsEn6xWmEcSl7
h8o3NM49RFcW1PJc20m+C9Rgc9nARVKTWxnhn1Cm9xBA4I8BES9xSgoZxMn4MNBi
KNDIu9WUMbGZwSuKExtgP/9L6zhJOojTu1oyIsnBovPG447EEYNXvATce5vV34TW
HaejSfadyp0AREaRasdu6pBBMr5IB2RWiHaQSaU+YE0kTl2Jv+K/wLaEfhIpUl3D
xxrszjdzj6M2595Lij97ObWNzb0g9T4xbbKUIW1XRO2/a2wle8PDzFzI6zxMsszb
JEHmPiLNatoNUSDtz+mQdlTvD1/38EKoj4r90CeQ3sv4rkcCFxS4bgBReau9b5Kk
hnEVjePoA8EdEeGZDzf0H8I+j91y/gISgOSBqo4IBIPbawB5+eFzF0TIy2Ddl+Vs
8pnmP3hsWihiW/n/b5JKhRHeC5F5yGtsdN6AzoS3VEdNqbw/pmdkocGsXNAIEG/J
G+Jy8BmChunqdvbJ/nyIOKRH9ueZ52pwbe/5qu4dYx0tte8JaYY8qDoqwtsko3bw
29sxsZC3Sdh+yppZnHJZve3L3kK/MsSg+MRhEyPBCFn+2TKSmeYeEf+aY8HKaum1
Fw8VKpYeZMgDsFq4XV47tR1/Ys680eQ45gMMWGdCmPwEaURIrpcGUivV0BNfiYdS
vckwQe7FFfXrzEPxIUpzD21U1REQVPnPDFn2gXZQ3fuFoInLkP+gSosja2UaEWgn
ZTkBvIAt5TrdX7txeASt+C7xrhjseSmgdcWmUL7bSJbt2WK5ooLwZ1aWzrbg5AdC
vNtmyQWYnBMOF3MHMJXLQfFPZZnhw3NpfJQ3ezG/6OTZ+J+4ie4Q4yHK2WLwjmWO
XcX2306qefqxW7NtiCyHsVRA3fVva3pHLJdrZHO+9ti4bvklI3J1PosCTpJTWBYk
UcE6r6nDeA7oJ0e79ByoyYTSSHhCK/L7h3ATJetAXbMQg2742mNLDaCvc7fYmEjO
wmMn8q5gyfFOh/diVLOZxp1z2/3usyvGIfHWudSMTC+euzsw0S5A+WvirqVui8bZ
OOKE+Su1Q+Lhg8LN9UMo9qDFHtSyMl/6rJkN8ELLyo9Q9XnVqGn25Uk8AWV1doHM
zCTvoiyohpeN2PQvInGDTPO/jup/AwZZvXdn1vpdVV3NMzFlV05KD4Fb16tXK9nh
q5Y4s2bedMFcjM9I/9m1CYSNTZyelT+5yllYNkdV8YwfbsaPpsAATM6dm8HcQQZj
i37hwsqHrg/wV+Y6Fhc9uUo32nNMYyC+aHu24kvwKB8QzPRCRNIDP/HHvQntR5vT
qQltShzliVqH3Zbld78yEjfQvHlxOKCfQwhXTVqKfg343KAS76NB8BvY9IEHNU3g
zhpKgyqIm9ZpAqaTB+kOawBMvvS+hc7OyjvQa7cdCQFbsSzS+lroyPSlCU1vvXA8
0A84gHKE8a16PNZOwqyoOJJ5J7KSP4/k4klTkNAA+kqQMME1U/cyOoHfBxOw26Ml
+TaWbh65i1pAnLNg+vM9ESsbOHQNAMARQtK/YgS3kE5poevNr7skjMSrKk1pALAG
mn/Z/G4/e4ux68M0WngkefJHEnn0W4BQhQsTvfM9AQwpCRvq+GpGOoWu91/6+rkv
Q0aBfkapL2xSC+S/jvIf9JpQHMBmtSa0mmSzzib/f4OXyPabmoEU1JJIyUd9l8M0
2gNHPwD2Zcmp+gWJhQeWa7nDeu3KS2oLO8X5p7STdPda59GmlRH/8IPrDcPBLbTV
l/aD45Qo8bBfGN6DT8fbEoYit2I3NFXQ4B7qsJLv5GeMstUc2ErBEahWT/12nbTX
kUbH2n7Yb4yUEDMsQVJkzmX0ZdoGqVtP09WMDGh6GpHxYs/AijaRwtZaxlujJ2SS
jHvYbPhMw6sYjJ1S3y+DoEYfcAXRD/zzB1MrlSa/C0EWUWjQcBNFLmJp2V30t3vi
6DxNV1PhBhDjc27lMShPtT1mirRq4Y0qCMFr2KnLhWPtIbPqwg88R1X7DunrJOAn
NTCDvwHgOX5HbZARrbQpYIUY3UsV1nivVhpWLFutVOcJruXIR2gkuX05aCPCKg30
C4/jqfdzEEgB2oAg3+CTxPAkRruKp2wytOT0wk9LUEP9oKVpW3R2gfXsqCJS/uih
ZtpzNcE7vfSmJvwQsK2uUbAg0IvVm9GlNS1uuXhKsbtE4HktOtgkxjGxLeFaLCam
JPXgUgiEKFKSrGGLMM1yglemgua5HphAZwOGKiLllGfAHyPjxX89boW+mgGn0qni
d/lGKTSknUbDY6KvQWt2wRO/8C7orDov9Pkxz1sAi+i+B4k3R/C5JVGhVQ+589Wg
09BQ71dckizpMlu/lzSg/kX6pbSOZszesGAEJkDazJcaLxQ+sUsWaJELMBcMLTHi
irxT6qYz9k10xJ21JqK8a9G1+rDAEhestC26Y9V4kLDQV96PKrWrrzZX9tT8jUH1
VbEJ4fAAKHQPCdYPcRXQP3wSFPwco+1icgnJBAR3Af28gIkztfhgbBEMT5qz3CQe
6GezwYiQHN0c3IztAbKN0JZqM2BbY8QMrmjzfm6jloUh4iqM2ae2lj8JxryPonMe
hkoQKD2m6ISvFjDyNM/QLaQZT8/B8ryjmOJP7ZQ+6TpAuMlA2uH2fueUxqSIkcA/
LniDUAkl76FYkhD+wUvZ+xPIUq6d+TCr6l1lfnhi/3IxB9rEtfy66y4YbLdN2dbr
B1xwrqJ/MgadksT2cxBihY/Qyr+dbfzZy5vNL5Zs5XiTW7Rwl+8n+BY/yEWixeuK
KHxaLFeQtvspspZbzgfRwspw1j5CWhqPoWyXQ0MEAaSX0Du1Hd7zLizbaUTd9QvZ
1FV89Fop27iSXyrRxCcafueTqNWDMkTZTcENLHEPqgRolxX3zJhC5Otb9KigLRZm
1TcpJVtYOHgndGqll0aSEeWeShGjNSbGyNSok1pIOLk/5d9cBJesg/rLnOTaBJMf
6CB1THb4GJzzbiZeiC6bnTFzveLCv6jXRBluAKRaD4Q7eh7FzS2mRDEZ7weUX3Hd
hVuj+jFgp7c/QLPIjh3Fw4ICfeFntzJpPVPYFty7hYv2gIjMi/WLEL3tW5Gh5qBx
OB+VUIEBwgxCFTJkPp0e7SL4nEUwZPTE/SfnhGF8J9TIVi54SjJrub23OZeA24Of
XBVO59nLgxvhQvh6W0IH0Cyl94sGHhwoGn93zzxDJna1lad23nQbkX45BP2SP4GL
Z9kkWgkhfGpAUQp2R5TzylsoSnfOO4IctBEIkQDoQhOCAHTU44QwTBNLnAInw/mJ
nimjMJG+sZyGxklTeYD+AGDX5l2A7XprDRUEM6WYQzLJNZ3u/AbZvLpBaXAHwfId
p03AuLU9NdlK0cgL1GNfZuQrCWIkK4dFeeHq11RUpHpQQ940SqnIDFFSz4z/Lrm4
jQZ9TYpRQL0zuXP1PrefbW1eqeduxKoCIlyt/2gv3hpI+6iPN3xIJbe8sH6Pm/tC
nxq6GeZcEH281qF47K6s0AvhaUzpJkiFGX+4wdjiPKyupq9W5TpAjJF0h+S3qlL2
Gd2vXDnGtyLs/4s8sTbYb+aoiLzt0zYNhskMbCbwxH/4azun24a3QuFlJYKLEyYv
qAjsBGtG95jF9lX5mZRGltQCcXAaBLPIW5yg0PUipsPGSdCxpKJSWP6i+89aDoeg
+jni28PV8S2ys+oyr5ljeAf+NuXDh+4s3bNgwatHhFJRF2ejVzgRCevqYQqUxrjt
haaDMeSDZTTeOwDwgXM+aOaq0T2lV/Dmo7Pl0g75c6DGFwno+B5W2U6QjZ/YdPzw
/HNj4UvxkL+LAoDrq/Ood6QZFqoxKf5rzei7z6Gc9EttiXjDJxlIvNX94mVs38Ro
aYpzE3UvVIoDuM104fo0HqVK4LGpVLXtkId9x7ikUFrwItRBEJrBe0xovcarKTbr
qO4qNnqRyIXuKlQ8tk3wuq1cSUacbdDRSEuH0WErjAdR+1bBjgN/sCeh8+wcGFPq
/sp5oMD0Z8wufIa1WXRmy99vxgI/J5vJfR4iBcrFBdNS9zKBI5ZTTa75TcqpNWtx
5LmkkVCMaOwDhZx6lGg4wRjOrKyzFjHP4QCnrywVF3aBofKCEqqpWP/wFeR8Qqgq
O/+RCuxG2aPhWL+Uo9mu/edAX+HHx5SLI1nrhXVgDmwUiwHi0ZT2UjLGlG0HXX2X
elUveCgAEZvAKcdJzsv6tDMr2m0cza8a6RH6yuLVo0RGq1fRFqVaFJYRyWmLDT54
sDRzZUOXPMqK3j7VWk5OyJqnSJVSIFWgmXhMh0L7U2KTOj9yXpZFtk9vq7YJvauN
I6jWY5k06TszkOZQBKWE7PKLcxumMlvUNxZV5aRhoG0yQpWV/WtcBY8MwjHtirGB
D0CoMBnPpL1GDmKKY2cUBHZrFfSeGyrXimamw17XQqCGvyTg70dIg05/OWwoEE6e
7KkC96fWrbrn50Rrcu0QsPFL7U5wevY6lRQRKnwyXZxFqX4EvFoky/tlf5A+qXck
IUz5Okq/rEG27P+qYTjB3mJjs7Yhbd7XgmSsSTUjVYzIHhgOnEazXt+uQkMHDZWn
Ror57zBQVhW1V7M5vZ4O167M6Hvcp/ODIrF8PDZhDwu6R3vr7MsTIpS348j6blCU
RnJdmeJ6AjXumsiJkjqWIGCuxyA+bmnBAMFgpv7rXIyfiKFIqkynATDhp4JiBSzS
Z4BBzWxLzpf+cPhXUEaF+mHW0Bd1cfyjirELgoOjKTUY7mp5qyov9JZ41wPWOY9f
kHU5W2vvHZNWQfKNqZMp7dupnZKE3Gw3QfAe5NVoPL5nZnPx5PYhrjrRUKEjuXw6
BF6BzejVwIQbY2iD6NRpIsB6vZAs64sUR/Yl268cd7qzL5MdA+U2B1P34enFEjjd
rcl8Tt0dx+ActClcv6/PtSos3/Nr5y9XmS8Zb06q3NzwVLQ7VKVCYxmdG7bgLI4q
P/xOEs0j3Y/jcvxXl+HtsstIGmu4n8hOUDnD5rQgQRn6hZw0HM+yyEjultfBrp1I
cNFiqsWnj0vJeHfjjgTM/6k/qb2OVfmzu2HQ1X0FjjEfiRYIacfHBSMrOBuo4fTU
zZdf1CDXVfe80zuB+s5QxWf2phEnF1bfR0kuI8O1pI/U+OjUXWIVPbTHJ+EdRnV0
Pw9nDsuQPetRmVHQgfeSmfA1erZKtxZcbz7cBpHkIjOzIsDk+mDA7RQlihX6vsWB
5GsMfSac4YcQ/VtNgOsXRD8Yy5QtwrgTDVPQUtymNKKnQwAad69+vGo/44FWKgGO
l7qZjCfiOFTNEvSjr02dv1o1lYYUXN6F0xgvwHSw318G3j964/C86F+wUx2Rsls/
zqgQ8MzpPohZ89p06pOnoxDnJvmbJTlSi01iO0pxtO+35r7tcfMBE8c9uj+MVP9z
im5dmKQuw9/d7d2mW1Hk6PNcRke9oUXE7V7Wtuar3W4VGIAozG2/RAjMz0CBfPIo
DdlAoCpRasSmbsrKrCwvKgyU5QezMe2qDI3pmO27oIOYY9lNJmFCPk7PkD58dtx2
UElKlNgRtbd8T2c6rc9HHxzeDC9BNeZiHpFzALgiWKdcVehvmXO5WuP7szGocIxg
+ywFFGS21XTBqgczoxkT61Wk33diRJ0tqq3+hqdXdA6t8IUWnW5vt3fQpPYgKMfC
h4r/qW/psG1GYgEurou55kk0BZdJtuGTuxmZqHLPtmDCBV7MuqX0J/md2nQeqf+p
DWB9L3rD1Rmw/3PfnsEiKZolTr0W4xtzgovqL0oCmirQgtohujXFTT56qdsEAM9z
UnwA6Omdho1xa+d8g3UeS9DJGK9zmjSGIDwl4h0uYm81koghkerTEB97JkYW21Z5
YPkWqKbZkUvru4IRJNMW8izK0mzmT8mFlQz8k472PthJWrdizxXYsfFTeKu0bXBj
T4dShugJcHJxNLzRFUV/41giexWlrLsLZ2nYUnO9hC+CAlYHVLPlg4syoz7aoMuQ
to6Xx/VAJfBbcY/1m7qv33hgd/SJXY7z5Q/nF4QztNFniUzcVoMWX9386tLlAl85
lClydFWJa9ZWxPIQjbx5fdkzZEmwuyz1DQwSl5FKuDsaLbRyoHa0T24Ved0d8anb
hNduHHFup8wowW7yCZsXONTDO01Fz8JC+EEovTGvlgl89g+H958/Lp6cp+KEVOJO
Yq0uJI1pfwA8L9OQDGdJEDExgiiPWadj+E2y4kCa0IQqxcvazi2ts/iMnsj/flI5
lNQ2AwXXN/SYu++u6ri3KETqVfvn1tS6nI5IZv9aV/jITDMQ3iw0yRwQbQYe3+w3
BIMw41hwemZc3zaFlNQoTmqj50ZqOLe8uLg8qt9ojZYzdd1KJBo+qqeuEIiLqy3m
gvnzW/euoR0mSYeIi5eP4z2Javo8doaV3g9W/UfkucbFtfF25amUZ4ADpn1NgH97
Fy+/HlfYrVp0fwIDnOuQhgFNKJOFzTzwk0JZrZkayjmNeHAjzCgsHXoRP63/l+R1
3eooIxXinPxD2dfRU3fPPZ9GTXGzLJOo1ZYUaXU30KJCCcRT0K1mnhMRxhFHuLPA
3V4Tc0mQ4wt9JjhNzWdz27jnWsiH3Td1kGYr0gAgWYvT6uzXlbANtGVixkJKjP84
5RI5EPH8NaIWG8DlO/aRVvP+OVALCjS46LsDDVYd0p8bA8eR8ah/jc+x5Fyo1/NR
k7XikiMHdDLrfrUWrV4P2b4412n5QJOQxkNAlcx3lNvKlXwZRfulPdoOsq1YT0jG
3nNSg1y/WF+Y0ynBYCMOAYexsu+DKs9cuidWw6pNOSKMAZVr9hS3g3Z4MwhNmOJ4
HNncFTIzMnCjkRqrgCDO1YFO965EhKBqmZuw49Swezgcm1CbXps11R5ZzYcfpd1C
fd/MtVYIX35ybpg3daKatmygbQxs8nGfuu6WmcDUgGBxPDEHn5cBXxHOkDqZ7vz5
mkkfDJY1QrBL0JVzazZPRAy4bmzvEUHDlssp3E5soT7WuymM2bvF1q96QxWdgNF2
2YnPRj90UBL4KJRRWfb4jbo0XeNjhl0hw3SDCmnRhb14cAzkuk0lQEmAOvyySlxF
q5GAv4B4cI1eHBS6Re955zgyyYKWjx/mehkl/rMzkxVU3pUrFjdyFzOg4Usgle7H
1ygMMW49HO9vmnYuD1OT+5Dy20uUKEAPho5kOYS/bfpbVdId2ukcoIJl1D9cLoLZ
F3A/qNPAAkIK6OFhq01I+jX9bJxxiC624UUfUfo8J7/AiHb/6KRSfalX1pIFWuyy
UfKNmfw2IcW10jwwFYl+8XKTFHHDQbG5uq9KgQ08dS6BHUtCXePvYbzKAvbHeb2/
oYlXnN05mYwba2smE7WIeWcU0poMETF72lXnake1fItH6WVHMJK1sEORMdM0r3uf
K1WSRnShuDr0S9bl9OgO5O4QJTUkCexwGNEAM8H5Dcw5G+n9NctwYSVDKo9ExkOM
j6Yu4w9RHaK7JcMT/PQ+EC5AFMsIr2KouZOJV2elH4luW+0etFLKQ83FmzTkhPuG
M6lLubcqHnSxWVIQ4MdOD6EqZI5DdTbQXao1Tt9/mVzjx+AociTatXYsR7dFpuln
GuTVEewWPfW1gy5iWiX+NJn0YaiOIOQzoo0FeGuYypuX3xMsSBNn2e55J6j6+BsY
IkXlAkxDhAd+4BDLNPWFoZg8hd6MxSMgUQ2Fmy3M6ka+luYxrKs5NGMrlQzhWzE3
nWu7uvJK82W4WVKpCt7HS0CN0y5M2cYAocmwYKNCJResiwRYC8pPBlPCeEhGGBED
hJiIIZK8ir3EWEXkkh6zqhyKYS4sQ6pkP03czkPYhudkCDwgkLG8gOhpTSMnLPhl
v8O5+5mZsJhPL/CtC34J8xp9x773P8CvKAVe8cuUXZWfeiqjUQ0nmQARjWJG2QJN
/L6pGYTwuEcY09H2HOwOGXqZ4HWFhKRyDXuKJfRwc5phSSAh5cnb04UAcZ/j/zuo
Z9pDEbDlJte/1JsQkxGufT/CCDHBXHwzofzesqEJJADUR4AdyehwvIeKfvn9DmV8
n2TrxsmW/Hs3YoFRFaVhUQxIRg0OXvY+RgK9Q+iAd3LA687xdbTEI+gT/etgHfYR
Eqqy3RB87tokRbLTSh8nepq6WQmEGZ3AdoAaAC2F5opH6oJ4cWoe7H2owBkYP6tu
W2lMG33hsb5G/NzmUpzQMD99BPIvFaCXXnKujllYZroWNFtbzoCusuKReXtUK93W
xGHkuHMSZtvlS7ZkJKHIjo5GkQ2ugGiGeFS+FI8bsiitEdJiuFzbGfvZ8HI7QTx2
9qc3HAxQN68JeOnsVwxYwlTicgog/XL/Gf5tRNuCpsXD+hNGdCf07Qd0pu/mab2Y
yfNnnl1ao8TtkR3O403CZx3GQ75K5OlRnjf7Oh6jlsiH/2H7dN92UxrlBNG0fCoc
N9tLK7wU1Rp5uePY5Pl+SFLs0QbgxzKUUrsgEkG8mhbAvaXbGo49Tws/76aeNOHb
irOoRyC7jVz2TohnUftAyQKiDx2fq4By+pAKjmU8lwRxernsseehrkWGAp6hK/Kv
mk7jjN9r6Yv0ZK3ScnMssLJTtbIcXCjfKoLmtAtrY/Kl2OIFCuFUHsGO5Lzd8amb
3q6qaQhwsNNVvpaBPJB/K7IawFEz/wPyJ4cWBz+5YJjNbbcbPrt7Y+ct3vRttA1I
P/XjZzDsUyaZGFh7zOLXxlbDsZLVmOAX+uqn0+D2OA+nmLodh80KYYyfhCdsgWbM
A8/QROyq+q6YipBNAYHmDEqTR2QHIE9nzfbO2Jg1WH2BaJhzFNDO7HPaWPEiqsHR
VYtF//8bfPNr00824HV3Q/5ln5PL7iPGusyE3jkOii/zv0ZE1JUsiY+7PPs5PKnn
Z3DJdo7nzIQqKKT85sf79S9e6WpEEsw4p7HtVyoPC2RnYL0ZPQhLgRnT4ojghjSo
IAKiv/NXuKXdg8WBVZ2wlYmOuXh0MQV4VccEPWk9wdpMveHv4nzpvPSToSKRwGxf
itI7z0rviF2LOivJ2LBIkG2cmw9PUYHRsjCi1nBgOs9G6Um6TLOK9+rR7u+zOFWV
46HMUgk6HTZDAPFwZZywi/iH0Loy2G3Y9+FCLltzCmx/znc20aZFFdyCX997CGvE
++vRCGpFKhujlAjHyZLieJ6Lap7Ma1jUnUlbzdXstbaZTBCov4KNwaH/13udOXOE
I87OELbd7sPstwY6tiL9YbpSzfnGsqKuX9bUkreCf9epGgdsdTufI4vvLpTbeVH8
R0VUg2tQN38C1GIov+ZuzwzgNwHH7S9Se9bcfC6k992A+dasiSGleoUp9IU89Zhs
5DmyKLDrrtJq5b0EkDz0WnszXcV0HMaHwKqFmgnA79E1sA7B4G5cw8cjmOBofgst
S0efwnxSSbrv8fLj7kQXA3fnN5guHE/aSW61A9oPqYoaUTSs8jXUJqqSbijianKQ
SSJ3gQnIEgVB+PRUccEtD2NwCptxpoHHKSBeh0KZj7BxA81dkdSNt0R/wipqaXvD
pfNaJuWX9fcFch5dFm7fDU2bo9qBKpE9XXjrlzWfYva8s2ARGJpkqh9e6+AAfErP
ga0P8AKD9Fm8Y/ynf4xEQCbslixEliiANrriqVJMoyI12R6k80peEXB/MQenRpnq
Gzpl/hQ2gTsnC8eyLpJTfXpLx2CrBFlD52vh9PnmTby/2xKbB5phMnPcu/qS0Kjc
6/s1X5jqs/vEvB0IDJXQsUkLcvyRq9aFbzi+g8/xGXg3uG0S+tEFLTzCPY575fql
0k5okUe1tKcUG7B7qu4ijXpojQrsTuiY1x6OBA3KdtA3AgOokgpxqwVUxZs4/13+
XRN+2u4k7B4DVfQ29Ard8PAngoED7UxFO4WbMfTPejAAlxmZUCjG69DyV3c03A2w
+ZgUVVAPUpFCs2CB4NVtNOzBiAEqZebKdnLTqOAFrn0UxRVfr23qiufLzQD7Tfth
QPjhRKqp7IZS1bPsrrlaDkkBwlSuYbmz+C6qiI9LmeT43gJufJ0+/PsLABI2aeYG
3UO8eocKIy1nLCdWYDszyaGpOaTa87iwZn9KcCGSCsBv9pNXq+153uiTm8rzT2vz
/+XDNgrgIx3EDV9X6ASAa9yPM0IFOBw9Tq1KQ2FcQ9Jw7q/cZ1eQSNMAEpr6vLxU
wxe5zBm2bk8OplYRBQhJDkBjlWHoPRw4t0sob/+qdkLcOEbNEyrvEBduQ/YTtXvd
47Q+/yin7BKca9t8YChzk5Ktu0QOKSCBPsAoHymfj5t3xtIuJoKmnt1gu+v1XYt4
n8QEpNfVIzmizWb6ap/O0GnsOTtkc+gr/girtaBK8P70+pkINDIsepVYyGO7YIWT
05/K7duO8ZDTMV5tzi7VGCP/UZoQMZLL+I6GjYTioQE3A1MHHQzR0bLAssJ+pvvZ
giHQE/H/o+M03dIFOPVeSfy98uqzUce83xoVm++OZpo4Xq3anBrknGAETARPxXzR
VRnM50OtiY6uRc3edCOzfjiQUkNYgnd4lQ++szjZAr2l5vXlmQO/cylLEV5wUBw1
HIkVORa6BoL+th/EY0OGEPVkO5afX+kp1cBSJ8BHcsD1ChijKgW98lMdnQmqpgDp
RxSan/xWuaIxqggXjgbI7CZVJgHyBoYHmj2l9ODvDxk2g7Z5qE7NpC/FVXo/qWf+
evCuDFlUIXw0zpEpf+0rUrbisYk6G5w9e8fUT21beTmqF9QlrGKAm2eMGaxewtxg
/n21Adsu6+N4XdAjV4bdlS88JjYula5m62Ij7DAjpzBkNGCCGFAh59yFyAlavJn9
KCTOlurO8IPUdZLZ2ngVxLWKfkxgt9iu+tUahrcfy2U0FLEwPavL46WambEclRrf
3rD6XCCWW6Rw6O1sx4mWqd5OtUmXCppc3sBa1UcN+VBu3Ac9aImQ8FfEnyXl1ihw
el+po8xctGt8Vj27fgC21v3CIJTK52GwUc6P7ZcB6B3a+OJHLHf7ljVJnEvAT3QG
LdI0r4Kc/wtreNEjMfQwgmsdGphPHho8rCpyoimEtSycpV9ZXdQka9CzvIeMzAsm
NJ4N1O4alORdeR5ZYOS0NyD0AYJuCpPnyGJFSNFR1mm/1YLFMqsYMUJL6AppN1/X
5xDq1735Zr5IinjF/5w9QhL0/zkE0CfNfQMWgDQQWu2XXLZNljtzAFECQWeWulm0
eOKHQhwpPg74f+BzZDL5UZyvOWyLtj9zceRvkmyZ784Fzdi/1GUfr1r0SzDjwg6x
S9n0NC+jhs6awO3iOW9pDp/gOIt+MQtPDdzsjdszywdqtjr+SkdnZzpVGCHftG7G
SPMZqJ1TTu8kxHvSvq6iuQz8lhil8gE9UGcvkpoj+92G6mYwMLPdpqIte1Mw3lhY
KRaDij+YKekfxobO7ZsWACq1HMCQJ9XLbKNrt+/4SD3EduGnVEAm+PcxA+aWPugp
YXYmDNMoV67SrWdeG0vxgD52gfKbnWh43wm/4E6YRlOLW+e2xjWsywhkqNap++/S
6/xri/tzV4qeJXzz504qfs2gywyW9jYS753Sf5siTVrNdKtHiyLMrqnl9+a6gNIJ
A/UT+6MvPx7CPtu/DVFxS5xdTaT3RHScvrqgRrutoivuvoJ3SqlYtmJN/AgRnoiN
Fmvd0T17JfyxegMr/99O7NpcDLx170MgR6EK4KCmOeHXtQ7MSJBdUi4rlhPwv/gl
5euFIiJUGAbAL//HDqBwQ3dRy90LX7wFWNsYzT3nMToERWdpWS8Uqx23DgJ6eQrj
CfdAPiZirQNMk28gPDC379L3rtiTbpdnExTxE9aNgODQquXDLyqBN+NphgVXew+m
Cg2f0BLJQI2tjcpB8kkirHONCQ2SzZwTjj7r4oMa7dejVXtAMjVQ9+DUFL6i/Z0K
AtGEuyOhvgaTQPUwuOw2yNW7eVBBVsyUTFel5e8MED0YU3dfR3jhDnVP6wVydC9d
+cHi78TorV9oWvSsl1Fh/ENJZuh2y5pBZXcmhWUXx+uU57wxUYVyjmLFrsxmJWnX
AXLHFgED+58KW2G6g6XlurwtLauBcK0AR1u/Pl6md5A2HNiUY7KWxcJR0gEcuVy+
u/badYXcco9D0hyYSkvueoWV1DmE3Bxc2KtRyOB85TRjL2Hhik/wgoaydFWUwubq
9aAmBKOW56zKlcY3rn6Ouk291X3FdGGq/1jhlEhHJEzKWKLYe28HXv8diXOm/Vpv
a6F3WuZyPB7wYlahL/feTQIx5GW41kpnjZn9iK4ShEZ2ILmAh5V8SF6YP6abLsBv
WDoj6mpiOsKSDmg5SAlYQn591e8fosthEux+ZrfwzYbwmR+hHRw4XxAFPo9ZcSau
GQifvWDAJTFNaWbXcp3UkKxliR2JoICbtSqgkDIq9fW9YqzExSIqXDgx/okh06wc
PzOT2mFwYsUqiCu+qEIWO0zZXYkZQ6sxZak6DxXIqpCvpotAwDDGTXiQIfWy3MVn
Z+uT0C6dd1sQaZEfkNcFr57JBAkn6B33hnVZpYOPcBDOjREGeyq+nXq/5HNe3li+
ZBzZUAPoaTV2KfhaLZv2VWlh70PjtxmZT1/h4TpYYc9NEuwej1/X4oaksYe+8jqb
4Y1NjWiQS5aDyiLRz2QbLtrSIsxdH0GkjkSB8AWqJMlN/Sb2IFpreZ4I5vpjNYwu
CKGn7RpWTLjZ1b6soHHFbCJQAgbwGdnsNLsIsJQHJAUsER3odTcm8yWAMzL39EvB
EYszYke716lexbQEh3lipOWfpIKUCe4LGa46LeLpb958FuA/kq9djPvndFZszR/n
RDPDFs1RQ/HkLZrPApknHJGzipPAvEZjQrEQJEG3ig87jgz/cO3BMb4AVdi6rnLG
45/EmfCnsb4ZqexzEsU0mH5oT2KDAHRfjkS2eTirb0J2iVU+y2EVGalddK3vRwNE
4Ek4LS1ujQ2I7YoXpvtrFv45DjKNlGc0wM4AgJuL+o2P2CV7Rp3FtuUgCW45E3e9
FzUwvnC+kQv7ayi12KFzDPIKxkTFBy6dHk6BF0dUNlxCi+URyD84hSuJlaHS3TaJ
D2VF/Hgr3hAXb4HZCtzxqiud7B+AIzy+gCrQmURG9e9SrKRlRa+Qm9lVEt+RV1qo
3FspGgfG5xdeic8K6tN+EjZDVPk+0sfp0Gojm/eBeJtArP0AyC5Wfo4ecgU/Kc2r
MCbFAE8mG39nkuyYQE9XYc5ZdUAT8xdznNY6mJ+l8/JOqXKgybtZ3Yr3GdYrL4Ou
6Sce9Pu7KoyZq3KqnNN16vlrR8VjbuA/11ZqI0LNBWnqVqzfVoxoyVP/pNhvfUvC
1tBGi0XA+Ic8q5et5UBk2/EAYuFP6UQVoKYGcfWeRTYpstQqOl+h7wArjRbV326f
QJv5tJxfFJ8BiWRNQuEdqJYTGx8zFzs7755w1GoaIYasdQIFDqSZNs7hbJt+1uv2
am1y6i3IPPsSnDgbJ+UWgH6bFYVKwOZVDCq4jrz6JsKabK3718kxVtlbwsw3DyYS
1/c3bUjFuBcAYX/DkakeYsSbaWjcgG14ENr54ApdaXjIGXqVb6aPgVW/bhZ7tTkL
tBds+Zawuk97cxYF1SS+9Za+BdfPL7NZBFi2UH2BK29xskZFpfQ1eQiHnTO6pwtY
89ecjvFkm67+VrPVL4hVrmvXEZL43oWnQfhoQbntSHvhXA2MZneCVGVQxR4fevTt
k5mqF2XdcbkB2qIBxhFbvkxmZcqks99M1hpR++Lz5WcpmhN5RfZZokCQBTgM/NVi
D/r9gmnzHavZHPiipabkyHUqkxp1h9QqmHx+SbdnXliRlkW5jAXc1+Fmx5w8xDly
OT8w/zGpEGUTIKFdsPbY2cDrIsywg3vRuC7tgDKZ7AwK0xZ5usrGipH1S/VaIUB4
IAxm1TZhVpK5uFnFKNZjJvgupyFAhyfCngvsTwaEAYgnBLbWkr6GPIWCy5uF5tJn
dIxMus3yPz4KGe2vJI9yBqD6jCcGZ89gP4mKS8OPC6eh+mjpZeMkKRluC7RooujF
6h45I+IynzcazxdGBCTJddyLINj34dKUninAMgjKP07PQoLcTn33SnAg//G8nJop
Q49X7WFft9/RKiv5LNNOQ+dPFmSEWGsTblICp135VLgs8phlaF3JlKAhho2X2uOQ
EQ7kdLznX1jgxZ6iRGcBAfNqa+eJNcme9SNvY2vXUuy66SufvjaM/tVTgZn6M6SV
4TpfXFLaxB0HcrdLwhig1021nLo+y6vjpZyCc3NcJhwvWZLru7NlyFCijSJvUh0g
kOqhtRrnu4g2rHRjR2wln9ug1Obv3KlcSKBnR22gASP/H506CqhZ7TUU8xMh3fZx
RwmU7acO5Bnt6YO0g5vU49RJ041dKQIZLWsBc+cG8xguuQ6eXptmPVY8by5+RBS5
e+jnuxvK3Dk7wZrQh1c9E8w60dDn7AkmOAq1SEAPc3glS09aPJ49FqcydtqGZ2ow
UwS3OOxX63ozePnR8z9ZbPHGMvARxlDcLN3VommaZ1Gkb942dByGF2zgr84Z8sGs
BhF87LppFc5ik67uygxWruMX/RNwCeFlP8R5warLpwBpQw2pgRrRQv+2Nl1Pij+V
9Ms6ULZGG4DdzvS6gtFHFO/sXxwU9BwbIsM02qBrvBnpeV5MGS+WD/cC5IQLWwh5
zoFj7w4sFWOz1FBD7UbNrjmOWMxvawy9xjYwKHBwbrLMq19VbQ9txteaVJbLC2jq
8AOfV63IKEamsdj5e6s6Q5wwxwO5EMvwH5mGiCSfS+kiZeubSdUFkNzAbHeW0qbE
VHnk7D85il7qK1Vn6bDzp4LNbGGod/4Edq/Dy9Z3K3qos9nrQT9bAd5pbgG3JdKh
mvi9Ixof8kZ2MuEQ9eT+dIAi2GipzfXeTy9SGv5ZHXvEw2Bn38TTHy9V8X2taczS
CQpSJke8WlbPFmvP0B51WYrruBJeOARVZtDceRzup8Qxv1KFDFH6f1BHHT1fZXK6
1FMzCW9J8rmVH9SxFHaV9AWwsEU3+MJ/r1/VMoeF7tFs3B3Dsxhd/Da0ovZYIiBQ
IzHdMfQns2JR3lWNGUo+4kTH8lTDTUp4eVJ+OGdvRJogBngVTcLJJFWzg3LSEE6f
ZYKtcumOJNCDWynbLRdRoX4RULW47WUnr/+Ytml4d1WL0hlaxCQHTkc5YbdyDVGd
6FBi3n1PHGVTM+AunUlXGs+l4fSxPIIvpilA1hjTkOZPuOJg1oC7F6zmAeFj5FF1
284qRpZAqwy6UpV/Wx1/tVNGqgT2jOoY23Lgfoio8nwjB+yf5rFF0RFl5GxC0HdM
2fw7HyYJhskjmbIcrYhvTPitb6GeeQ1iyazP4SeRXxiM29x7un2LaywdFg0L/23R
vP9fG7cpnU8paMOBB1QBVYJ1FV0cmjd6idY4SUZM18NILeeuoUnZkQeQVKnPKaoA
5XFT+TnRPd1hQtodpK4eyZqXjXLYrY0WGPyFUklUl035ScvHiSkG1w7XdRQG8P3J
r0pwHY+wMYIOTq26xCpHW7vTYNMcWwDRSQ3Mau6OTsVWjSjOz3ZYURAk9GswO1QJ
XzIeywENYfh20whTrH553T64k92WFTcTsmoZfPRNlhMawOFLxMTVphpjlIh/p4D4
3TBbGisamaF6F4j1AthG66RYBWNSkwTZygir/HNcRQoRSHmkj3Se/XqFJrXQOXda
Yp2XOItDL7ghMpa5D7X+nYklCekgYLyLkYxGE/abHrjGxTP+VSdOHdlhtwxGjChD
YPOPTb7tQuESVrG0PipATxN2RvlgT62ThS24VT6F/clfgRC9RjXdKsNJa9bwL44G
UqsOyH/xOcF2dqY2wWJhsfGRW/uNhzEkcbnigwzhaegzkDeJlQBRFI4euIBu2xQL
TBDLm6QQgJHWx/c9aV6R3ewtkBrLlaqqnuqt1GsLWYuEZxJppw1JM3hO27JhzBlI
IHLYc1vnri0iLNVvas655jU10zDxXiE9JqCu4yrvyJ8Bl0OrbHAAJyYWmKRoScMC
vUV5nUSqTqNrLC2FQkI3Bu+BDTW4XaHsIGDfi+1xQ1RskYw0qfszXA22zJEHFp0A
gddd58SCR8pAq/7Io8U1vcRcPqWJZ/knz4frkg+iA2aBngT7qOfF+6mLzsJyiwPW
JMoZIaBz/b/agFek02/MZKPooOd7lie14Y13e8MTbukxHVQINhMgPrXWpX16OXJk
jZ7ManU3252w+EXsHCWJ9xJ27Wyp9v8fUwdrzyBqKTGfuSdTIo2NncLqSayTwCPz
EG7oJF/GUmdzUjrS/Hc0TPLBEy9/RhVRhJa5obFc4kn4n2UcLWQxifMCZL5RGIpc
+w7vnlgnI7Cs2O6ts1jY1+lqNzmhgBQGsZTk2QKQKiiGLZqASMooqCQaVwM8N1dh
xzLjGQFcGO2M0t5AOUwgVvRgex9wJVDb0UB6uZ6S+TRVBWgTgan93RIce6qLvHQx
9eAHJpqz/uzPeYe1TR9bL0zvCfItcFQNiWMp4nDgAOGGuX2VhMs92sXNK4SVmsTr
DetQ5oQJUB5nNIraR2m2AsusDVE2llnc8lXPt5sD4WA54JaL93FsuhlPCnor1ZWN
CGw9y0DXGkDwwlCeqBJ90LTS+ALaS/PrPsDaV5Zt62q15qVy3SCGbPOFCUPyUoGH
ysDdZWochdNLCBeQor8om019lwhiBmlhTanVwn3DCnOL+vmxigT2nQa52tGL+Ey2
WxYvSXJmtK3Mku5MepPMXLHQgKHt9Y5SRzkCayhULl53NPw2af8+ulie4CuCV7Ox
TmA00ADYp3f1OO9GYJUmFxaH+YHqCziFxCgEMUzKzJ8OmcvzMh5surGtCmC55tIH
brVhWYvPKNnR/b08CIlwMPhaahMCigcc1sTbktsNSlSlMbLRqJT2is0W1KbjhUnW
qD8y225LD3I9dLe9X9RYpYpfiAXN1CHoKuSyIEyyj5ByW/yGg/8oy6pnVxvfuip2
r2lYOzGgLhWQlrnt/rVYbYux4rxS1p4avqPBiAlM0ZOCVVzyhM+kkBGvAXXfcMdo
3t7w4NusAtBf83zgKHKuEG7QNmyMGdCCtDWtJvNEkMp7OEhfPOeiDy532WyBfJdy
CHJgv2TA0E4PCsFiAPABFxg7ghr94YgTKhoeyr1iwYna6jTkNfMkJ+jatZhZOBzo
NSP3+M0BJmDcCdZupAQLv+lWIrIhObKUPeuvwrn4jsgS4+CJOLACQautVfxr+LvB
uu4vUMhoVtC/eH4PMM8urXVsRSvHmAC1qvoH5+tcrKmWGg/W889ceCTMvrZxju6b
aYpx36xnlUBLg/8wMagK/LBohBxDJMUk98CzLXQaG7tLrPsjGtmRlOwPY4sfKe5a
932wtSCPHFSTh4tNLi39Ib5NMAwns4tDqmwZyID92yEfb9ENzMbVRicvuWxnw/hY
/AKiN3oE8SRHw9FK4CithHGdfWyqW8SxxLg0tL24sdvYwHMihKuR8UqXvZBO3q4k
jCPAzUbqgHBW3fdWF2gN3MZE7FAmYaB5BpVvK3h/gmwA+3Bj/utPaOujgg04U/Cx
/CakXXsHh5W4U3i40Iz/R8SXk1xH/63M7mL0EpWTmw1cZ2/MI1m/mHj7fi5WRA6U
j7HTM7ATPuiHWqzE40EwpsjynxDuiB7BxbXRL0Q645EdOdYQ4Z9pZgOoJFSze8Xo
nZbrLmDlJdoYuzcLsn3Ura6qu4ymI5hbC3TB1ObMSeQ33cFEh2NHeUO+AIk+8lEX
+tlq7omb/yPUqGD3BeVhmCXHxX8Palv1gwYZDQhv38DvSKC9XxOqpevihMJIgtkX
M5KHWGm6SQ8ieJjzqeA1hIgCRjh8Ke+KUkOCLYrsyzXXCyzWWtnwyfWDm8jgWq1q
TQKScFOYWawpLTsQ8MCSUlMCA/rIyYtXe/LApuFvnK8VE45yROla9/MYwWRCSLqk
bi8sPN+AZBqYfN+sj2wolfyUPJ82zsB037sBMIdjKr32RcB5D52QW5UXElxoBy6k
sPVeqqI1bb4dKwa+/2gvNiLHcE7FIQdw99JUwdhdFp1PyRaCS7jRzfFiLBUD49Z0
k6tzad2SpY8hLFg5takspxFcBqmHkxHMx2k7i2ZKZExUw/BIr2lr6zIhfvM045EJ
aEEDomcyIqrsWFzuXRDEALQdu7w81U7OLu1SHq6mQwjzMZ4x2SniFz4CMxTHuckt
3VrPtrR0E59+5QEF0NbGkiMOmJvJjMdImUI0NXhTY0PVErXmZitIMjc8VyyuBVII
Zzn99UcElV0rKTTnnfuiUa2BJKP7ZwU5LtYIOsCpTAAgLlpKrQz8F2Q7XJWmFCQU
DcXj5PShS7g2jxY9RDzDD9+U3vrRyGH1AkWewFNiGtwvlf8NSrt/xrhpVXHtQPKn
/DcsHMcIcxittJtFTKCZj3UPs6UT0S/LZF9PIqX/BQ0G9Fpjiv4HjHi2tawskRbD
KIC96e/VmDuPsUXx7pPYS+ZZcIqVBw82UZPrOJmGtS+TgsjR+Ul0bJiZ+BhFL0mG
US2OUltTzQtt5yuWl5HOqcvVb86/HUwhgEUvQ8CBc9CsXKVlhGMw6YxTNHvdM5Zi
dxgUvHOIoBjt5mg5Iop3fkK1qlOsuZKFj6KAVCvIJ0C7/zkk9gzfNP+Z5a77koDp
jpa9icCaul5wI9FnCTIl9RAHkPWWcYf1JoxTjQlzFAfvG1FRMYUKcOIsa7fb/YKD
8Kyl2QJhr7mzZ43/VVjaJxuCfi6v6TzIJY49unHvglmad8IJGFai/SYsTFVkNk1R
BzXfcUeJfHyl74+YmRTbAIThOIhWSQMMEsQzeNHI3G7kDRS8jWZ8qYuKnKEK3VOy
gu2fNcBNAr2kqtTB+438f6uEpLBd9KXLeDm6yGBqb2w+m85sXw9aCFwbaWb0JDiC
oPuKhvOdfYDvGnyWAqCgHMW8bGAQdDVljLegW//kf3Q5UMh8nH8gR9RM6mj4uemo
azd+N6LzO9I98XJsakYBImwA5/fobNrbKR1lHwqgM6uZR/OotI1SVtFK+IwBZJeF
knd2ptNIWexdw66Hmh2ewwQcCVjgLVXXofyRtRbAZPgW0TJtsPhcZAsNI97z8hxS
AAHcmL5RymYVs4QUS0Du5N7ccKqdO1JGl8B57gil/ChZ+6D7ciBMFRx6gZDobKqZ
OIrdyt2OZ7PRY3TIVrEBFubrd46xRzbe/UbIAt/pZ8C75nABkRN/A3W6SSYQ2/MY
VbPLGvh+DN3JrRtP1vfw+KMlkI9lW+lpjRVoF21vWMgn0UfR9EbuIZmxfDlYrmcO
j3yDR7Ods3ivhT+IAsHQPm//MPXl0B31/7E4v8eqHjhmpUlmc5TfecNLc8cINajx
/CiAgbaiLp62riofTiOU2lp3qy0uMwfMCQLmEOc/JGXdSNiCzTUH+nGCO4oxtqrc
C25nzdG2VjFyK4rq6F/B/ZAV+W+BOHw1/CeTnoj0+I0ApYOMpIhmyAsohK57BRVZ
wB8quyNVCLvCdOTMoAn5RhO9yfjvh9e4ck3CXOgFTmonyk1f7hZWt92N1FY7vEZp
IGATCQTEkp05phXJ+LIAnwvAm6x8l22D/a4YK63rFfvU2rx4BHQu3CBi2RG/Lnx1
rFtp/hqLLkfwbd42RpRpj3wxPcozu4225rjImAG0YU7TWZ3bTOdYf/sS5dfqGmEX
fbquYxVI/qYVTaHLQjLrSmrVZ41j5D8DjWke0PeWCYQlpIbeSTZ0FvQ5xPMQ+mZ8
/5v0dw09FhRYEiGxV92hFUWzCqXW3falnmfeOquG1SN5A/vEJTnDn5kTriHKh05Q
wvEXWtY6djDz7Fuz3yMHqgNbTDiyNKgnyG97HHqJxaotQSDSt5Qnb7kWHNWfpODF
fAVwkwq0YDbTl7N3aB/UVyc6wcw5eCe8Tv3KHgQ7+0vd7m2kIWOo28kRBjzpN1oK
UdPPJ5xiQL8QXGQ6/No5jexDbdNRfuVjg/sCXI+vwO++zJ3xErp99jH4+BbDLM+9
4DFiDRYaBCVk84Zd053CasCIACkgAX5f89lR51b9SashI3EHvs8BCtsYZ3uRSEWv
EYpR5PQvlsIQR6xnNN1hnXXtVkPC89uulLMS4vca+Br+u+gsobMi4eMAPEE742eW
6Cy9EdjAzcZ7rKOvrzGlRMsx7Dpezs6wDWK7NDQUzA9obcsOU2KhkOrbBx89LzVL
5mHE707hk/oYDokkpvm78KCICIT2jOX1hgAnTpennBq7iNOjXQb3/FTHjIarPLYl
7VbRVYw/4sorA6AquDV07P++nYuGaaSzcGa/xQ58wOc+JmtJ0vLreVhPGCDFf37l
VSUGUoCckGr5xeQYCcn99m0KoNl1/gfxgOl26wMNHRTa4F4sssrB9bJliwhc3yPd
oE8ct2LmCuz4taTR+kJz5aN2CbJwCNxiLT3LJNd9o/9JQp/iB9khf5SHNfx0m8+k
Dn68koISwqpfTUZwfEq7lzFTic6nmxJLoDTPiT457TDL1A639YZsNjbi99lyfLI0
5nMiakA5NjJjT5GVNRJ2CdN4zh4SV0yEYstW2P0tg3FC/8NSC5LOQ0kJOP9VoOvC
Yt4c0q5v+8YLyZppkISOAUuJDc9hfCH/vQyztwwG4tQeRYD8POC+y0TDYNXWV5qr
XVd/JSMHPqxJf1a30YZ/IPXrP5Upo96jrL4+/3kp5Ejj9qYuYA9jP8WLxjBYhYKY
5juAP7Z7r553rTirobS3cM86XdqGmszSr4bw6B8UAU8kJP5MjTXyZBfUH6MNVzJY
RY18TQJTgefrBH+868aBKQkbww83QMDhhCguL5930EywPI1Nm1gd1X/AyXgmuzSA
0XQoxH+q4WyosMvisaewtOvhwN/HPlOo2xv97NsCI7rFQKfBqHYwKWqBJw3vmPiX
xjIz7Jkh7THTN56TKd2IwHczD/oiIM3EuQVCmlLL8JgpN5H9gZyZqyrr9l4kZfwG
T7GS8eQ0flA94ySdGwaRORY8l3dC+ReZVbi20jgPltbmjrJkqFtcqadG37haoNz4
RPja3KoLQvQY5UauQBhrFrXrEtPhIFp0GOiDVooAwqelIIaTreBth1jqzv2ej+/l
uArCh9SZHjPRp1jB/jv8c5xzhcMqlEQ4LqxbLx3OhitiaqWvn1XRxHuiN2Dkub1g
aJr+r30DBYEzb5xdFlwUllH72izLdZZ9GRA6Zljeydb4pCNCMcxhDaNQ9qF2qH7c
AFfF839PnQZoC76JOlFnkqNgB02g4qCVK4FsB3uZBCjjkaKcCVFxHBB/3s+a1EL+
qJi7EKDj9rr0mM3Jj5GtG7KN3Z879zqTDsVd6GdybpwH8aONYxjmXfzP1o/b+mQo
hjLK7pMevSz6ynsXe32eR3CAd6Xmm35xvySUQPq8I2zoBJv7xp0VvzymkInO2eon
Z1lICRjIvXh7y6IgDSfwT9SANSUqmBIPQpU1gACEwR32v18IWo6GfLc4NpDjSchc
YBI+86AAABGBl0/lh9VCSFR6CLjyzqQOBBwswmNR/lp2ENf3Q3n1zdRgBU3vn8XM
aERLCSy0CII10UMZQMrzJWKSOtaG1FdFBNwabSLx1tXvXDrDwIc5HIxy1ALRPM16
1oKj9smSI8TT4TMMAwjGZCpHMY42Z4a0Hmhv+c1abybIyQeJQzoYmDyYSrIc8Aom
eKMV4YUNRgkXjDMdkj6eeNxdka0hrmb9u2eWxkfZicKsvOZM3sAJTez3RMsN/9fz
YsNgqMjAj/uyDLon480hGasvdXlQ24rxvEdGPxPGUGsVRDCjgioO+HVOp68Wpyy7
3lny3PCtynVc0VnQdAIUtAJ7JmE9PNZfBhxhs8Fm+BB2FDdW+ldCE0uG/0PQcJHl
bgflaC4eea5IUMinXSFm58f3QYwlqNswKJO6Ce/80ieGiS/8G+KT3lPA17aJMnpG
H+ks+za+rrPoxgQ0ZMXfk0SXT8TdW7Z2O2BwguJFsUEq4shL8MyMkOUy0o+9vHON
ZuY+CDjjhPnwyo+SFIRuli1pCcau5YxwrfNXD7/3Wg70Rgln5TrJh6/jvYEZbk/U
dfOy8A9jN2ctQJE8tjnoZZ/nnCoOkdNBMY8Pyl1ZXuhrZ33LjAn/f571lH0sJX3k
VdhwNNx5jpacrArTypaEoQwONp1C41tegsUzAGNHmGDFINrFgkrfV4+j4Hzf7zYx
pb6rMFTpcjIXn23K/vOb7jCOpbXawCdy9753zQ4sQjcw8xt5EtTBfSQC8H+14LqZ
o+7UbkswwUGuPLDHllekYTE0sg9K1O9vKTqspeDCQmUcZDzUddiimF3Pz6ks3fj/
4FeGNCPDsdn/XDFIgEp4+4GpZtzku7SxKxMjAgoBB0G4KtvIzamN8tLTlazMguRY
pSBNkuWb2jCASKemCHcsnZFDMMwraHnjAwFiqyjXCB6ra9aJOxOgEOfxEFlatBkR
6X2NrCci7d138DhpHcpE4NVR84GOtLZS19poo8O70aptR/uSfc5sEM1Kno29UA9/
fgUtp9tEHrKVPC96hEgV4l/KukbGkDLRHshGCmtTq72Ou3QSIMKnlZMupMN2z+UL
oC4IeE/SspGbYUb7Dk08oIr5MVkLgGttOBXXVMRMHX2PTzEPyCxfqmts7Yiy9lDU
A4QXO4cQP1ozfb+5AcB/hOOFzGRXzwt7LjxNPXLohmanJJZCuc0mg13Q4kStIGC6
7DVTTvP17+DgQrsbHZ2S2h74NzbXqsD2R43zqHisZDJ6RiEoquyfMIu7Pg+vyBVx
a7EXIrqZ3P5zwzbMTv5qKx1TQMrnTsgcCP0OBHz7OCrO9dw4FBgFlTTWrhlEofPE
UuCqZgjXfpsXPVdW8HoDfgeMEIU4VS6qnYPM+eujx/U22w++xom4fJn9jAvJDw8N
Eymn9rNPYvQFMOu5AxEzwKpgWrIFUB2WRCg5dHifuAFGgt9eBe714HTs35n5Tv9j
Ehi6AYZacAW8N2HNQOq0UY8+bvXvId64ql2cXDGMT/GekxX4T97yYC6I4te5D07n
0Z1vuoy/MixFTqO+hcLAGOKNCPwriC4MqpnwIKiX5fOATOwA8k1jsnAcvUJdacGl
2QMnynjzLrJzdJnOQjQY1F2A0uB9HMp1+XqO14Q1H32MkI2rmM6jL3Y/YYnUnxd5
1w0DbGSMzUZbidL9VAgB0op0izV4lBrcpAwqOuiO+SpOuL3RaPrskWzghjcisYxX
G08mDKk4aYlFnfDy3ouvrpR15XKqkvAEqZit6HQl8TGZgzbxQZIQQywtt8No/oUS
oWWbwV8WFZsLri8C5RIP6fGxg/OkDi4KKYCdwAaW0wGOIPRiP2+DX5OnCcHBPzsI
IlXq3cJ8aT4ydRWihYjGhzVcVGqfGVJQ8iyaRoUkXiVlCTnddA4BKXvBcKwIMMKA
rRRXRv62GoLvNrtliWNkGv8uURP5D4nufsOo7AtIbgNB42voAe9bzUXqRYLOfBcf
uIlwhjQ9BsQYCg+3jHtuaRt9VcPs+9ygpiguAp+Dlq8L+d63yiul2LjrUvoaGmId
IFzgNcoKao2nYr3x8mCwFn2Kc3L7CX+Zuf5Izj9D7B1F0fex8UYDCRWAElCn1UI7
FDYzGxGIWVlzZOrQjfKhShZMLrNufuXs22O5OZU4qO6cgVxZ+9Ea3SOkiC4OVPQQ
Ph9lNBtBGT5RwTb1DJV95MFgAih9lXSTA9gP8HUQjs/oU0FdM3mBfc/3RVvdHl60
dRfABC61aU/twOuLdkCWfbrDY/CUtOQeEl3BxDfonvlZNROyzD4ltV2y7ebAj9S8
Yv4aTk2Wbnjmxy3HDW6qHGt+3UbrflRmNhcx4Ckf7ZCzH9K2B/A4CGCy9FUHEv/A
1UdUIYPr4IAJbkVaN2Q2+nZ7pPv6HdRFhbLETy5kpgRCjRKSyQwAPQTSM9DTm482
z5medKeyxpIQoXtEyT82lTM5y1vR/yqFvfuI3uRCUi6UrSToP6dqEQu5qXk3ov73
5im2DNIEGO7l5Lx76jrvuOR2fC8zO6ndWkDtqRHLpNWOX0YSZvfmMemOa2P9I5CA
1SZqymRmqdVrx+vONgt4y3zjodlTXiIYZqWbLOpFU6Fkqhx6Lp9xsCaW0bruZUJm
lhAy4w534UlrgaJdI88Q9aeCbbJ1dOXqEXTaIaIjckXBNWP60aw38Ig5v9oSsDH2
6hfLHS8KbUdXG1mqyrtw/mpg3iaqvf8ZR2ZvGSlksmma/iFoXcAl30IqNI1YKNGu
s61J5r2sKxlJ7Pg363QZebBWMToKnfaZCMFE6cPi8A6OjIbVj/l+gfmPNWQ4cZNF
WM8pGMrqS19C7OAxE2RkVeGT8qzCcghYuEVr0FdGxJRrKm0NjXLSwY/5eSlh4ZF/
6bCJz3yli3BBhnPEAUFRpbH7rHPkV4jGUlWpH0xbcdE4iLY3I2QnQUCvmFB7Y977
3f5Z0vuKnP88LFqno1ibmxWSG49+nu+uF4XUoX/sQMRtVWN1tqEC6zcSUnsSlfRK
ssAlMjEAN211sIzyj8VeESTcaeCLzUCTYVjAN2LczdhqVgKCtlQFAu+hz46JIbTT
kyt+o/wUCGh3eNa2+Wilvm7Ts5aJtVU3WssUw4fUto6oziS88gcZe9Z4yBTkowPm
SZBvlHwREyaQIL4DsJFCvBcYWZP3LN6p02l5oP5ALzNG97takw6krDHhaLCpI+JF
ay9D+W5nDtlosFpssisnGXNDPpqHSnPY6dDvzcssEbL5M1S6ql0Vhqc4aJQdn9G8
4ZLVG2fZG/WAZ2uDzIeIutX8oMbJzxN8g6FZFJiMjOlpj9MLIjYDOe4RJ2By8kWP
ijn0qaCwmT4jG977vKfRDQhrNK30qMSjo3AEU9l/U8Qj7R8/8d8+uFFfRGkg5vo1
b5TjVov7ADKwvh64ly4i5+itoiRofYk+Ap84MQmoD2yPbq8mE64I31N3txHx3yOq
Mq2AM/XV6D5SE13MxMeFrnRsCVZci0+gWJ6jiUBIfTYx5zg+XfRstgkdXedTSeYf
c2YGqUp1IQydSPphoZVzlfObu0nfNIQxnexpWv++zZd9XVYHU6flUPsflCo0Jotk
iXIDchj67AE2Gd9mJOWgsnP7t9QxxwuVSBJVlUC9nbFi0ikteopmNCTJgiGiq09x
Y9lGmTWldwsmHlg5br59SWtwDY8CSOe8Ib6ZV0uYBOFaUA9qB6B+SviHueIJfRY0
qSwcqMxtrtk0PVEWV3dBF5zATbpmTNzpjWioHi+t9KXp8RxUJbjHW5eSyudcqZ8J
pbixwGwrny9iE7RW88YM7MgNdF1DBd/TjOj8pEKYDfLtgIadZTMIE/d0+0duvWmo
rbzFRpBpjuXnpixdBtsa/KDt7zdz1xys2hAi6VfNrECRw3iiblll76/hbIRggA+F
mi0TdBujeVzmroQWnBMKB7xsPXQvXADCWU/UYPWpUpwGkvA/Pv+dL8Bd2KAGVzMp
R/veK5NCL0QdyZgot/mp0pC37PzMytDqikXgCUBq7hZskrWfnwqfza7KGsGOs+rf
+sN0ScfqfaencW+cL46d39XpQ+VR1s65qtIOWZRerBvNq+il0hxHqFIrkiSN9QSi
PIrX4aDGWSV1mJIEP4L476M3ylN7OaDTjCfclHAmn4oJAdqmZMP/jXpcQp4SX7iM
I4pSUFxMQw/Cllz12KxY7JNJ44KEgtxr+PeCNw94VfrRf7CZBoAhB7LPrrV2RB2g
zADbzmys4BaohjBwzCijqQvgeMZserYXAUQAgwqqzRiE1K1v44kCeXQZei8Bqerz
GXzXLyelnpRbGH6JHeBW2WTqdxyngU2deGk/n5f0LvBaS9sb/XG6CucH1imN4JAq
6nTH331eyIQsma5ndJZWhKpGwI6ZxjZuF3b9oS+RKYBHsyQ51YOgAe9eRlq7UZhL
rhp/yRk26L/BbVVS5wrWS3FzGONI4ER7fIHhafNH1DMPCbXdX1GvU05giVYUXPhE
5uxXCRcAyUEGm5OOYKICtI888ZoaAmMSRirAI/x2Q6AhBUbtsGB1yytJ5FrnD7+y
Wy49em/2HeeZtfOW4z4qzNjaxvu5MvTNPJ2reWR4AFqrxzIHK6q+jmwSJfp519T3
8tBfaCnhy6hJIUevq3gUf51gvoApXtkAWeIqCT+I5slcsvjh6EH/oM1WGRx0btgy
ln5djuQfXUCNn7exPIXXS50iaAlzIdxP4S5i9mMNmQ4ChBr7Rtn3PnXLe7gG80Um
+YykpatO1u54Fbcd+fK8UZ8WVHzPIksnfuRxtRLeUFx+sLsKLeFVvuI6eguMLCWo
92Ud0VFWJDWhzVIXhow98MwCbq1S4zclmpm39DK2BZn6C1xRaPaVWiDpHzL5mV2b
pFVqcTIhZYbrLM5vpcOZANX/5w9PI0tBKnpsjh7mL8ubu75URvu/3eOFPvEHCCBs
MP1Kl2AUAgXgQUONBPM0WkIboquN6Gm560YVKRvdBHUfcWv0dzgDJ6v+aXiES/Rm
pCzQTYcQzpA/9fGKp6zleUpKXW3ho6bbVhcPd6y5XqQ6vTDMYLHeueJauUQCYdea
ZoGHuW5aPcp30JIGXaAANuzmNqhblzxyG+Uc3PkSi6rKGXYFJEpqsWe2JPtiRUqQ
Uw1CF16nyAQISamHdHThka5sVZYo4XLN3N7YjwUi+LvYOsECxUV2wH5Xy2xZheJ1
qdPuXtwfXh1RGhwNaCXXzU+Iv7ZG7MM13x7E0OxNngBFGclJ+TyvhZJTTj0gcWPR
E7aX3bl26TUS5Abulu3f1Jwi5KN9vpDO/rLAk/VJsYCfyFxW8OEL/ffUwC+GDEjm
nTHywT+VBxqTFk8QbBW37/pRskQF3wykKWiz8uiUTEvCuRzdq3h7E8RZ9COQuNsK
mkPvFSWGki+JKWsvvwbuKTfBSkjQ+mOA9OyqMan+nt/NcLjG+erLCnqMW9IeHSDH
gAx0qYi+80g48cA2hxuNjQhpzrLP6AmDcIIRHd1alAc0ubeOMpfdN6xUWX6CIQL6
i934iXqdX8dPkfXkGREX8xrgJ0Zty8hkKBNDb7XA1BoWLEFF6GTTLp7b9mQ0ntMY
QlodNRfqGDiMxEN8IGsIG8kG7ZIPO0sDU7wQq9qSgZnhpc9KKU2L4routhvA0mEY
NxVDdiQJYml3xH3jo6UNBIX4zUo/WPnKjLn2gxOc3sbq4APB3ZTqRa05DGWDGXJy
SLgGotzs8JNZmRJUszAcIptrWrmogDzr54vIG7Pf6sOhHiLPSRrthn39yO0ezUNq
pYMXPfS3Sxxho+hSZiKdsLuy5lcBnTvwwBOhriJ5J4Qd7MMXJ8JcZjbpU3qkgrlx
8yQh9ke3s5+G7eOB2A+dr2N7a17ITkHxat7frd33AcWBDnLZZM3yOXwYmd+RQ8ax
BHYyM3FDoO6yeInhrbJdfTq0/cJ4XVP32tS+Z6Ny75dsRZb82Qx7LLbNfla0bLWh
i+llQysHmdCTLuGZ8YSNIPEj0RW+qk65OQOj90g5HB2IZ8yT4QtVBTFXOJ5hiWfO
9jHpyL+2VqmfiYDOrKxk3JCB5+hLSURkHTbJLqzDVJNJVVzvOe0xZLeYedse5kYm
k6z08TpUYRqsWnpRmzSyfdjga0BYk8itWIm092MdF1Td6TQ4O5txi4/+2oSXUzB7
jgV9QUz8HQ5NdhramzVEFV3jzZJmGsNjG8+JO50hWYEqEh09O1w5YTQWacyjbmy3
rXRKqKPwagb2nGobyh73R7x+kCeTGSIZxYlQUqG9OJT2vfPXJRCj4mZ3X1AGEV8t
iBfbwDrKHlWdAtokuJms0T3Gi3l+8o9QNcMKgD/U7Cdt1AUBoY9vh0j638gLcFZu
zaTdamI6GDiDKFuKq2gtV1de838tQuPBjls6tMTf4dModvNigvjWQhTDxvaVrm40
7n8iMElR+v9/Nkc92j+sBjPLKSFo7IE0l/kmqDvg6Ce5d59eSDiL8TZxei1JoD9j
V8XgnZnGr7ilQWj+f3ygN/NSyVH2yPN9/qDuKQWCdBVWP6/Oc7nqwfalsh3F3R1E
KHwbpqUtjcTcWjQiZMyRYYxDapNfenIo0hdHjRKsw0mC6JOOJC/WEY5iI/Dt51z9
CrUMBP/bN8z6D+k9vr5rAJ2Iw1IcM5+uMGPoNMVMAjmzPBQeqTIw20L2hs94gyYG
dkBvWCILQlkvpIMuqiO2y6draW+Q3sk1o/4sL8Zi3g2wIqAejz+veSOeTB+BN/hT
6wRJFnflUE9ADalYzl729zFcgQY6giJE2upahjhaGrVYp9y9TkC/tvAxLeajYp+S
xIhhD4De5pdjKQSGyb11MC3pm3oQ2GD+ss7jHxUghyHtMOPg5bO1vQ3D/73n2lO3
NLXPLm83eI4GSv3rD+qd9ayAHQP3CymYCdTmF40GAljn3B9/cFG8XUI806FoQzG5
eQi2t4Yz8pxV42lrMHfYNlFtMBjGJvINkY53W2g+DEAsV514XCTXQpWXn1FI91xq
/vAmVIwyUM7rFzsWDIccVSHGErhT0aCTPC2uis1JKoh2e7UD0f8wmxRsVKyEMFb6
wHnl/fomTpVWjDPB3BiMeCZ/GnSgtR+c0glGEkviKqUqtTztGUv5SASXdmBh6qAp
QPAyoAGmLO76KjA3Drif7RTxceKUsTvJFlFwopM/zXWlRY0qPPhEH0V7CkXo1dKk
VXf1CMJ6yUnmb7iBvYjr0eVo5BcExsp9IxtQ0CsMVk63GOWuoylnGvD0ZWBWTQDL
plcXbd8Mrr4rqwonPbZL8H5QG1Rkv/gb5wbyAXL2ZlzLy1++U8OAyVuIwewigWEH
1uAfX85xK0HWfa8a3Ea2rdhOD1FRM7Pwqc/3nW4OyMOGKsgx26l1Z+DhDGHkRrvC
/V9tSJDFXFpjX/wtdTFBABhE6CrIwUtBOvpoU1PRi6tHM1t9TMlhwMMX7kTOqLw7
w8T7ErG23lUCujkhqCDx2NPfSPlOgpvGlOhVrvwztv0EkOvY3Xoz/cuJEygnBmWn
qGR9lkuv16xVjiKAZ4z4oezfiP2izR1h1j+Gj+EeWXxG3fsQco9XLiFwwKaB06Pa
yPESNOBxGVaJ1VwgnrDC0Sso7sJWHRc/G25a9ORCzEy7fxoYtOuIcoQ3JmUqY/8F
ci2Lm6fE+CcpoCO0LIQ82uN5dpsGBYklKL2v3J8g559SrettCzrs3RarEuZ+TgvC
J+kx5qMgUJbRcclRiyRHbcDwyuWNtyaFFB6dud9+GS0q6rjpcAbrb4gI0sUOPpVM
EEBzQq3Dmn4JgrIARPFcw4T1srLUJW1aqIFK6eF/EzCKp4r2jLzkxivJrqW9YvgI
gD/bdXoBX3NVhvHeUg/Hr5GHUpNReuc916ohvPJZT9H2Z0+oeFCpF2OPDqr0d7ft
QHbQ2GUyZ614l5YlJxcmnH9R1nFfAOYnM9kzq9eTa+CAAPvTewJVPUNVRDBeRxhk
v5yM+2CmPYIetn+yjFos87e0w/YFnnZq6gVbaAN8knBg5f7W2+gihhUX3lf/dV2K
j11rnga4ccRG9McKRCn949jOaY1WwXCzDThiwKyocZRwfsz9qHvXOmsEZy4SIR1a
5dYi5JtYrP+nzVI6N2NzXuXuaYDc4W0SzLsDFAa+QcOaQ6iigj+egqZ76wxvorTi
yA5UIEVswvUChQaOUysZXVlvI4tfjpmShA5ga4g3z/n/Y8vAS+97dhcMm3TZbhy8
zBlx7lSmu5evJCWc5ebzM4n2/eSGEM14NfTlxeYQZ58TvFkHMW3X8WDMgtInEyaT
wqnfYZTMkkkse22sAhYBZ0oFYQqmhpAdgca2Fnf/ONDMnhrqnubu8sAlB18l7M+u
ofQgCYNSD3j/ZQN/33m1owNwKj9ykW0xdCxS5OPT8NXjpe06DFOiyAFdL3ickWIX
grAZymzd6Tk+AEZ+nQanKAo7lsUJ3jVu8GV77vlYlUyobefO2khju1DLjZl2Mf5T
rcUVb8iLCeWSlLVoTcpSSaay2xvO+JBXIU6m1qMt2Emx4DahIkA8T6c38ba4uT5U
2WHDAt7PnsqPtdkyOHhZrjBPKOXpNJf8dDFBmOypo+R0ROathy/s3trNjGXLgQT0
KWSARak14Db9ByDKLsJ8uo0d6VUmRvIXMaVQPCOUmOKO2qM4eeHG4in2gNK1aN4c
WUlbecCAGvoEl0xGL1TIAaBMP7Kohj2672Z3StxxQItNHCO7GPX6sBweiHvwmqDK
BJ2THaUWRLlhD/niYcozluM0jtiQkENpDUPugGukRdDeOpqcba3ORMmdZ2tHYEiM
D0tTJOzKKEtqTlHqLwCT16LwL/4zpwnmH1Db77JXGZxbk/u/Y+HakNP8R6LDL6Mm
ET8v4jXhIOYa45VvfJjNT/DWSPxYENJ5eQvYghrGmQ7PAb8AnHIpAETs+4fUzQWd
S8dahmZsjYMPAP+2z81JjaKNMDxauYuUvab04ymCYDUaYkp3tPOLf9UXBGtbca+0
9z8+2xpv1zUNiS9b+J23B7TMD6I7nA/5riJ4b+LGUfDAfZFn+Yk43XGcDKiBWvS8
3+5rgmqn/zh6dfkgzGQyGP0zfyJ3JF3htJE2KBoKQWaTM6yZV/jRPGW3mvXRZu8d
2kKJnzVTPSRuCLuiBkbI2fgmbTJBEOoOM7K0ttui90DmoXI94bt4eP7YMrR4Tv4l
nSfnfy+MwBChkzx7kIVizwTjSP9wjyUNT7ZKOMrqtsLlTETBWWEZA4IZ6RCmM7GF
mPwGcTjKWAaoa2nrHXHe1AGuFAHbTyplbOb9CD/Lxcr0ZRuX0He98chREUz57P2t
hNSXc+5lt1GDz7vqK0lMF77cQU4crKD3sjFqDBv9Qu72XeIj/LzWrTYaa+JeXOZg
iTU9Wm6EXE4aBwVPytgvoSmpl8GxBRaImdMEbDMKVU4Z4Qqn5naKTjB78ZDBaQJL
7/lr7BQ3H9IjKOPZ5RiIHB5LyN3OMAwmKbobpsu7DxsthPQi/UcXuwLZEw75k7EI
B9xPXAVrSzbcAwQUOxEkJqn4DCTKOCQbfPdnvx7dZ1D3xEOU7q7FPPmtG8SdV92D
JPFcI4zzEhuNKBPkM6cKFdYzOWtRmdecx5QB/dsTA3J4jmsRtZxzz8rh3RyHZpYF
kOzf4ZOWdTkhxOZA/HgaCOnheWxY0E2J2foUtMIa/OxPOF98VICT21EuNaDSqUY8
gpzDBkmN/qGXSxUAenS4CB7RCAiC7h2N96ew3rKYFlZdCzNkhB3ioW0VBUH5S8NO
YWTwly8weRuv24xxOwg2uxOhWj09pWCTI0Dw0zhQn8JpIyuI6/bryYdylZLkzaTp
ePtwcl2ZVAJBqvuXw71H9hh4dfSjs/Og9o7+GphYG5beNiZmai54QWw8cbodY8Y0
boG6aa+EddaRGnHgN3pXs8tXAIIL4YfA6QNqG/4hMFHEmkvDKLRykwdel43bxHhP
Z0WPYRCSMrUJgorvSX7N9I0pBmMUnXKXvVHNkzL9zop0pjnJ1J43ylvOJOa8N6J5
QCJw6EfNy8yl2R1XB5AKgASOh7d2Pbggb+SUDN0OaUlNzA4IDgIGfqaUHwVOEXtL
PtPrCBIxg30fZ7oHRQ7r3ackLLjGr/VKQB0d2Wa58993eDgkvsomoI7sHfxj5yoj
AnZufg9wqm6USCU240SmLloazX8CMRbLGrMkhPqmc3U8YmtZmnrd5LKbB6XTaOeX
KorkGqGpLnXXJyV0Fos61iKyxNKIm6PwGhnKOfOzHEZfa4BoDtLGRDyrp6Lo5904
y9lD9ZxwUoJQ3nTiqIUkWOkC+7u3VlPcbojzWXMmAqJ2XJnse6hVlXya3kbo5LSM
0aHTfa4C0R0ZSNxF1JprdwdH4xgHuJDKxNS71sYIkAubIrxxT5s0+hIN5OmFre5w
dT2cA3wzqIDza3AzmsAdW+C2BZ3FBHKtkORZA/VxWQrLzn+hLS/JGdKm4I8D3xcz
2KQvFC+9bd6mnz+gDfj1GR9c4RvNy7mTLhNArN509lWefw06MdjW7F12WRXAjqFC
ml5EjvTNvLmBS60RqTHmQZDkGhWfknPdz5DIYsSOgkwkEUVlT/5RbB/Kw8EWWeA/
JwUsm1syfPi5cLJT7C9dmoB9ACZGRkVzqJ8OXOQaPNYkMZVWdB53KMoZf2SHH4v6
JpJOjOD4KmGg67v/vYgKBrAF3fFGivrz3jQnBv2+vI+nJ6CPvCKt10vO2lOlMw6N
+pYWST5vJ+ZbWYlNkcChu+lwOeo9pNKNY40SfpcvmAkm6uOC+aZOiR+ZfxDMCxxw
uBwu99sCUgu1/b1ihwH2W/Ysu1JT0bWcXZALAGMfTYKSOcIpk63SIaRJCbZQZL2D
fBa5PALNV6jNjt4swf/w9MjsnK2aHCJhQEMwO27chwr3OUzM99eNmCjYZjqk+/gi
k89a8zYs8ZCCjnJ+uQ+FAygYr3nuvtyXNOGIF+HL2D7otQqvAxsVhmXlk8k+nVR+
EHC5jsbXiOhrnAbuGM0D9+sTe2zZF1UINecpZwhHWh8Ju5GgrdDSisjp5ycDeHno
DVvAKpXaJPODM2a9i5YowdrM75jSsYiVZevOj8mN8IjvLy+sa/HwhhhxwSNzOBY2
PACq4wO+OzhRzYryRMQAbt9yBTFKgeh+rXhMBvPKMiTW0kvfDKLWuWtxYs8o3sZz
paPma2+NdOfZDYvKz51/U8CvpBmcnlzONXnBYbFKvgyH0f9OJaTgRhcb9Z8ctHl7
JngxL8FOX52eapDFUM6gMq8/mi7ueyFO+54kO256hKWP9RhdTjp8odgb45qg3qAI
cy0+ERRdqt15C2hafS9Hgz1o2rIchFJksiajf458QyOU+lFGO+gPKgMGExyd2Mjc
tyfHvAl32YkDLV/g6yQLmoS1TCMBybJy4KWxGXxbobxPGOESnX6AP6ioMj3IZHAN
TmK/cIYCQXds28+/wFQbpXXzNq0khOtERAptFoMVqyxMqoyVmfy+Gtcnjd1YfISu
skhq+3kTI+kqFVUaOECtyZPwL8/tmXe08ZU6gHp1vXKemD5vFL3a5+F1kXOCnE2A
ByP/MEXCqhrPCZwMAf1ocWaKCwy0U9ls9MFossYfCstYXy2EWqOl0XbD+ovhYd8H
V1jxEKRKDvMeMIpdkFS3Mb+xaGV5Jm7vwzuHxsQqb2mVTB7lfCkEry/C5z4GqDzV
EyYhI/ETzmXMO+Ayjl/AWdm8lpGVApPMefRoWPnEMV8AbHQsQlBmdLee4PTMaUPH
JJJLOASlrLJoW3JO32WZ3dBycBT6cdc53E5uZ3icQiiRYcUkWi7ih/F+YpF+4koi
fCa2s1WaXMMXFoko8+SQftvfByKFldUywejEcNSScDqBJcCol3v1PKKlRVhii5vV
GW6068iv1NJtl9c7T+jD/nKnQBB4hfDw7H3T7fhNx0YdDh+OKc0pvqqLzoJMRptl
ijDz64hczqOIcj3tDvj43YUqBrfBHqG1n71bNCCBnK5vrI8Elh5Km/HGuzN0VMFs
+9+LG0HTXJxN0rmDv2I30o48WPAFh0GViX/z5wt2bpiyo10h5uipNHLemLPuc4z3
PzMk68ZjPul5A1sTH7BxCu5JAbDlCEY4xs0PNL0PaGpIoiLY1zsPzoa+6UD/dfdh
K7DCMB0/IafS8B5cydblWAarLsgXxRURE7l4nynmfWQOqhZkxgo1xPCtMSrWUX5d
wi8ZXZDRvhQ6vFqY9kfWSUj7pkvhToHXnrMeGZbWwaJC6+cylaVaODe0TSseuEq0
cpD8/cwSn6NG2NogpyiNLaUGXjey4zRHwnyBjRAGY2H+2aJ361q7CbROwPPaSh6t
Kzonos43orj6K8vyIyjurwFGQU1Xhp3SnsM3bP67TZP7835KGcM1gY/fhHXXrKZI
MCCHWcEymyRUW24GC5bJ7fpU1JSBVLq46zTJ6P+ESpKPRu1hEYhW0AvMqjdI6RBw
UmwFIXM8WSoQ8m5m+pjrw+0+4TbjCa8lG2MkoIEiYxCJTM0c+E7sD476yGQCgb24
fjc7Tz5Uj9YTwm48jQoADLWpZSelUwUfTZDSw0NC0AfFaqJ0wg+WKd6BlqEN273t
7tsBuVBYU6ihOYMGkA18jCDjnTSpyVLXoUgdC+rlIceHZh3b0MODrjMgYObJT6hz
LWGbViEXc/2txVE4h4IgGXMr8tTSX4HjAqitUmc6cPwvGH8eq7pQerETPIFZewDD
efT4odKeJsgyZChSHdmLYlCSdByl8SQRLZifKJSRvtfDV/Ej6YvQOWx3ERHh3Mah
CkRoD4/qZAFo3mFkuR8zDuIarjzKmlcjcDMmLq794COqk+4N9tU7egsz7UBv3Nbu
9W8zreOUNwnKEB3hdNzsFq1i2Gbe+jUAjdkTwd+ddkWuJrhgdxaTouCfrebRPlqu
JZ7mW39C046667mX5hG+TH5632UV7z9YeRoHx6MXud+7gAEU90t79MlHLEqmJ6O4
Bl+q45xwQt3lv+IBIAfCFjdLpV4XcjtoI58MMfHkxDzDiF7igu3Gn9i6uxUuTVva
D71Dl6+KS52x7NSfGGLoLUDoGwDOu7Yf+cNfGDI/9S1cczyPXD3EBYpDx8V7SQeE
2v5wIVT/KUYRdSYfcITSM0yWfagCLbf03wrttE6xMO9DkQn5FQFGeS94vtUNkYbf
1PFtBNDKFcmXSpUPQnQXhjnsizFisdrLWXG6RLuN2YGxmxIX3W+OGMkY762yfqp8
chYyF+TaDpS+TE16BUpIGVyMtjqh57ffY0Ji3Es7I2vth8HSROjrZZ9JUtU2/kMK
ldnxMo5FD8HMSDl/yVwmCFgfUJziQpMMhJfgU3B9fRtTpqrBm/GlEwDy9W5k6qjp
V9GaIzFg6iIEHpMBXImV2Bh0ocjgSwwY8GXiTa4wyP2bzFTALxuQ5vG401NXlB4J
kqecKrvkeQaRXTUCfQKFgQyMRRQaGpdGIsD6fsBHSfksYrnM2ITs5EP04FwT6kwi
HUlNZaNAHb3b7M6wXP3DnVLD0Kithol02mQnn23laBqE0BLzL6LRiOFnISLktjC9
glPmkZQC0UWhZqJQuDve0+7U/euteiWs7nxDAsKgKaD/IzPjkekYwp5ppJbLvJV+
dDqFHFP5cT91P/26VwuJjAdF17SdMe4G1poVJT49NFV2K4peq1Igmp/D3dAhHoSO
fU2h3mPu9Y/ZLxpJwJAlT6TK/e+I5EZ0Xl5nEdj2/IQvxNs4SltpmpEGwJNIMCS5
SJpjVl8RFQS3gLfmvqwgLRlX90TaSJoT0vpxtPAttJWRzc75AplyWuVMNosEbLxc
b77cnT/jMhis51IZ8EVQvmciyXitqY9MOihv2epLIt7pzNw9wPlo0jSWn15wT3KQ
DnYxIHAVewK1gdbz5rlWZ5px969pqntvvkw8rgHnt4WMBoZ6iLQiOhJcrr5js1ut
LZp9TgcrVvo5ltFpYxs4EoEZ0wO/VzmjTbJJzZe1HpZTP9Pd3+spxoANpyWh85Av
9Mg3YL8sVRndkLeeP6UazBL9Lb5IoI+mN7R8c7w/XKfOeYN85e88uIKd7v1vrZ6p
ZeXOS2fRTUFO17BhoCiS+kBttH2s/ZYMjvQkigjUI8iTl1i5FLRyyqA1dP/+toTM
GMA7Sx2Q2J2ldvdrTf7JyStg5YWXyNhRXdZ96KfsQ3j2e2UB/lL8lxpq2U6FARZY
U+VT5Hj3WuKU6Msz2AZc4fK6wyPBhRH/vTLIhJeru9mWalm0ZuI+4sywYkZEQOAy
Fv4emrz26QpL258nxartJRoobDbU/Fq/dXxFxvWYEIOClj9oZ6cvyUP7faAY1xQn
JrJHwho02P3oUG9NZvjwrWk3e0RJLCVN2/DW7JwTeHs+6wAIb+5dlM+MpYqLx/3d
YYJjCyLDreDlJeWS5ckgoTDlCcqO3chnkm6wodhwAIdtMrWfyYAVJgbMslhzbOQl
pQg0eF0RLE1nDTFkouUhU3fnj7iXfNq5D6eQQVuaQIwhW/FG4QFG6Kg6SQsx/T4a
/KXaWF2sotrFExHJtpOkBlF35NcXeZAx7F2YDxm2kjqw6bQ38hH43ueCUMlKE4LH
80qcYV9Su7uQJn173Kt360e13th8it4TjUPHJRe0UneX2kR3crlaNdWh7N9KJ78O
TTQ2DBbGYk4H9hH4u9KOpL2CHDfN+tq+28q5efD5gB6JiYiGdDDF7PBnilHA9qcY
Z+UTtfqe4kNBvG1duFbHWFol+aAEDT/DgJcqEojkAxsZ+Ww0VbbL93g/vFjZP15t
zZPqnQgIgECaaCBkD0izeLFlk+CpGcjKF1olZuifsfJU8BLx4Ycc6rlYvIeqYSoy
O0aY/q2LixGs3YuTqJUvfnKz8SYkJIDgwMXLxtKYTknACIQzsCBW06NrLjOjX3lz
QFuEY/U+w/w3aSA8xz3osGSbZwjF0zGVOAHXwXpnDabJC8QcsdjQHsJeHtRFJrjV
ykYqboZN38AqfjZX1jEyvhzv1EQMDqtYuE53HdmsW4DOKWNaQjHFKVLvKM9ccsbs
u7zQujlU8MCqcSYXPT7F2bsYG/Y3sl3u3xM0+wL9vxv7dOEO4gb574FOE3GuRxzO
ERY2gXDn2Dx5S+0NUKOql5bfTKpQVS4o4v8C/lKc7tK+BwnxjU65poxbjwonxjIG
zXzJjA9apMSh882bPj3AzKHEvL2K31BRH5XtIlt2Xm+7Lb6bAHt5sQ1LO5npd6sW
l0OowcGjBU3uWkwR3VTsS3i0EEqC7F7pJ22MepAIK2V2Afxab4GwjLoGYi9W8z3i
19e4nXXjDV4d896OU0aNIpVlZzqC6teYXqA0iBF+BzoVrXzzBQ2xFlzTwcOHPd8M
+OUewGsivx4HQISozcgiDDtXeZcBwNTmqDAfmcTSVd2cWRJw1wMtZnFF5uj5TJQX
jZ/qXN1UKJvTs5f5mmXPqzWTmdrEBTDtW3UIXJxapiZr6FnZMCtQahwV+WxdD6CE
o2Jl0/s+46eJk/Ji17V9kPEIx6fl7DMuo1VC8CBVaZpgemza96odStiOmwY1FBfE
I73oqeHkbWfAbMKHTfNsxNI/lEs5KkZnk+yxIyukcP0pDCn4I58Z80x4FwqptTuS
+It+68XusP7q1Jk+TRqwnh771goiwY4cHS4KOBGjj4JdwsgUtcMQr/XVdftFcbZt
C9I+ZkjdZNnF7qLH93B37ObDMduoSGMbibmluBOgwQrB4AayA8gRNOZAX8duaTZL
BbNiAa6/em1kB52dCxBhyL0t324Df57B5b41BgQiYXIxLN5waPd+Q6k+gvnf+G99
w1qs5SYG2r4x6HP0lCgkLxb6yQWo67HyBlRggijtSE3d1sFLdwIZpUyhas8/GJW2
XXmcbIPfEffmJcN062gQyY93S1CJKMF6xTuErkvOkFodEITJ5YBwnDZglyFST7m1
Eu4zIwwQehEgOm7hQWT/n4OIb8Ac0dXrbncxq5KyB/fAs6J8oFK4DDNLxrr+P6Yq
767MSPjd4zJS0ngr6/9r7csfP8tTVuPHwQcr1yLv4Md9yh6aTJwEXh2N3fHUVsM5
qRKO8eewp0oeLtuEj7L2jlhxFwWL1RRDwHv9bE3JlXx4x+KBHcBcsR4Zgg+6EogO
f6LaMEpOR6BXm85+1WQCGaCzpE7r2eQrpWY0nnAcwea7K9Ah0gal9x0EoB65zTzD
Xs0FxDSYbd5Pxdm49gFZpKstd/D+WsmBJQcuhlDPWu//QHV55HwdN25qiEOpqPhH
nn33DSGHJ8jK6VJtyIw5fEy/i/HO3qx6idwR346I73L0L2PLCdYPkLplWXyIOQ7Z
WsqRBPFxi5wK6ARV0/eYYucy1RbSxdw5WYniDpxiRoRrBJldpqXKe7B2ImWEp9Kg
5y3rRU6LVpj7yjgwHmf+oZlYkWjsu5Nn5EeH+/rPGnXEwafOwlN8lKa1BjYKSgsi
nw2PdWHxKyQnnGA1v35Mn71Jd7nLFhRgVtKqfl9hBKIbRvAJCs8/BMQ2AcuOGhqi
4MZVN6mDnWRra1Ro8nnEZ/hbLYdqLPFqVULckY8hmvUqR+XaiBgG6L1EIsDZ/jli
k2pZWuhcpNdndTsLDFKV5IQxdZXsSAvpMf5wrGohbmyOnjqX43PEzPK9I6yzMCfV
yivLkz4C2MBczx/SPQy1POKe7NC1XDPYQIWbMpC0LKOG2mIbcFQBuPxl4zXBAk+S
v4oYvNCZ3m6NlOJC1iXmPhlrhivy4X0zbhEMHz1HigQxgYGkOyqAOU51y82b+Q5t
Kn31/AA8HtsiOFapMIix4/4LQkht0PqEbrA8gkG4IzEHmoFmeeYswZ2SHmkru2Jh
VhTVDDIyTSbjkPwKJnWiBjzZidTqBj/9sdlpS5g7nKKlNEmEXvE0R6ZqqwZ2+Qwc
DK4K+vpkGJsIo0Kp9xR+Ofrr5fwBB7aFAKso/r7/0xAHVlFSLiDxsKhMcuXf0LFG
bk98NT1OsJP1tknUj6ZFn/8KLgqoRQRT+y6E21dsCqxNYt140NQYEzf78lo55ixG
Ec0WmTntoEK1pWi5vRXimNkZNJers6KP3GYKuiORPw3l35MU4GUBFtyhHl2b1Fmd
xN/jZ/3iK904u6xPAfZ+iYD93S/MCB5n32KQDU4aqB1SdNJEVHEIUirPysLM6kEH
JvNAmfDIwYVD/vESOY2xB8CeyXpVN/B8bjHBi/LvfG/mmXZ1rR4FoG6Hx8qBuLUA
IK7z8BBFhMjoPdS7KM/B6vBLjTr+UqwN4GpF1Ye9sHLhDqMuK+tk2ynyhBXyQmya
39AbtvPNO8yMdPhqMP8HP/vArp4jayxl/Hw6MmcPU23L1uv4Ms92jTPjgqIqs7Jh
AKdTNkXsw6fi+tMwL4h6KlX+gJbJTMR5rgHe34trjiXTfMNHlem4aGhNv+r7oFu5
PehSvKW90Ryb4B9BS9fh77DrSKZDakvmHsR7leds90ahNgDtLNBhH6kQ+7h2k7fO
D2S+911cHwKzc6/Gv/TvWBCA8mGLoOi5DFa0LBppLFNS+iHMY56pVRgFv7l2Ehli
BrrR8DzTlPp4hQafszPYHX2CQn4VniEQRhRZn3oeZCJ5RyJfJHnhlzNC12vr7+37
EtK4DJYUe14TSmf5JfKNTWHLzLR+uY1eyXV7TPdKQVaXcTNy2KshDz8PIxyKaQMD
WJX1qmdJq+J3/kkFDmzrVDLnT1udd/S3iS1gITqOtlD83xr4XZrWbfqLRzSYlUWk
odCJSdq6QlferCnN0pA+62KPy5LaLsFq2hQu0q6PdW+5OgDKCvnx2PEzttkEXNOQ
5kawr3IIhNtCb4KzyQa3OH3iQ7BgGXa5Xa5DZUPhZt0Te+kcyNh/Ds0M87Th0jta
P+nGuiX5hxIjcAwsRaVt+XOgjxiiwU9mP0zh0fnP1xLh8Zs0Ltd+oXP5D9iKnV8a
e+0jcsjrbfOGQQd/ES2hdqQBOUZCY67C4Rm0GD0WTd1oKYjReg9iNJVEOkfOR/fA
9E0SUb1QYNLePZ+dIpzTuCPXmqr8UHvl0rO7gPU+Hm3BCI1n6zSpesJX7rVmWKhg
8de4+eFxFi/njmSD4JvYIOx7yht+sDWV6BfLJaxABjeZ7o+ghYNug2iXLwusgOjI
zSVvAr3jV08JUQiDaw6CklIryoGZf+L0z4O39CE95IDYiYvCrTv2QVbK9GzyuhyZ
/FjvyhoU9EctqecUwyLdaknwwBadgZjx8dOh03MHQg2s9K9kt+IBh460RpSUZFPw
IbOm3iF6RxbjBhBE27wAwsq+BLdB9tEs5m9f6yKSfxBoB1g3ZjFOUkCKccdXFbWI
J5Ho993rWwSafE4SxmGIJvv5idWLUs519fQhm9rg5mr2lb3qX3JwOTQCkVTngi7i
0wSMLLCrY49J9ktqBnVsthkbU9AkUtt+qrN0rAIZwFg0hxXv5A76Vp4B9NFj+R4U
GRZfDTHQCCDJpdhDPc4/A9OMZecePVnJu6dOJbrCOORpTugygGrUBhcmq+R+y5Dd
BcUxtPCHt+IMiWND6db5sq2/+A3KAQfdv1Xw3IK6J7X5ytYQTkjtgqD8QIRmp2BF
EDlNnXTxXbpsd6i7XPhHr3ZvGR0yOSGdij0i6tYQzEKdcqnDP6ZAeJUkM+7kYah7
4wr9fWG5oIKzUMkypKiipFEzv6+UsgB1zsd6YweDv7zx4kK6yyj+wXzuOmZVbGtu
ZGs6eLw2xjDulwiHLQsakAPcXGBd1DNEs4Ujy2f58hwhVmuH/wABRxdmLW/T7RT/
nfafoVSXJpSgPclT/cruoJ5yKKWu+3cbyHDXlCbZyWbzhQRMF0LvCyKBIiLCM6Ma
mamc7eP+zCe9uE8E2Xe7rzpZLIKblk/UW1LNG4t3qLy1PF8E5gwfoND2GB3nfYsn
mYD4QZ7PMfVZZglRHvhyo8KXAujpEHkSdTtgh1ke6EuZjprFvxqO7DlsTOWa/JYi
cpMG8dVXsQDNrN1/q1w4snG2T+rJEVTpKyMP/fCXXuYQP8sb6x584BWp4CGJgMNC
6dqa1+hoGHB4bYV1rPEu4nNHqwNLlaaY4Gac+vGnYGPWsVyPiNXj6ttNggZoxKJT
2oWFhLU4IAsxxgWi+5cUPsikX3B5FeF2bHDCHgw8Gwtnw6lZbg4t1/tLLKW8U2+K
CzY+xISlo5Ysn8MeYMSNU4QwHxbl0Zbgow41iauMX8J1pdv8LKAix3aOBCjtj3ER
ajfnXD4EGn0NTj1Cvk9SBvqu0KoEw+GZAK/o/uU4kvA//cRPEsHfzPRgKCYq+zDq
z+jbtZFNtIRmtODY7FJuHHQBWDnvPRa7E349JEkBGscfV/m1DVa4BVM2R4Zk6szq
pdAoPr/7gMiXuUmM8ha4Vu2NTKMOxguf899/J+p/7Dc3dPDZF2YJu8mRx7teNYmL
GsI0sFuBwbTDPW9e+nQFbVrmpNY2vv+f8DKcJAf3TxzP4pAS8GXV7hx0iKEjUO4m
6j6n2BFECtcDlHZnlrteXOXI2m371QRwI/1WgSCHRyNjjM1mKEGZp7SqZPGaARaX
pttqHbMWoS9N/RkeaB1qYddbuHj7wJDF4gXTuP+IN7d1s97Hzy4M2yfOo3wHjpr2
dhG8s46+AHeXq+/TcS4rqi/XPtK+orDg264Pkahg9MmhrqKcpHmiCEhCs/ZwKFdW
kMtgUcN1UbdUs3Q4Z8yX1InSJxn9qTAVrlclpoJfEgCxY4WNTKosyAP/CGFxJOC9
f5rJUjtf9ZuzpHv85RebqAKeRkkTyZSa+QSvef4TMNkdw94VnYdtoC/ulCk7dHGo
ve10DDysSOkb3eyH5kGtNW0KJSO8dfvp5cYTaUtgGJ5rF0Yz7MaP3bbRbkBxuWAD
0XHi/UN50XScPJ4dnKKn2sIK0qIlT/EQ1QfKq9D2dAdHP0kUDVeDcalMKeMwW+mq
jDBhKapSw0Neo9sF+QOOCXQbAigGSR7BZ4TBygMOisJJ5z2EX872ixpN+wSblyPw
Fj59Oak8VUs6g1dcNKmFKYxopsQtjlMS394HgkQtjr7hgbofuQiBIOLWYg9zzEUH
y9qd2snpNX7w4sCM2jifuIsPuaOdqQZIp3Rnn89A0rMwu8u8173ufgzf+GeezYV8
zDcNDui8V2/q4OUCE8Ynyc7LvBSefxm3Fi9IlAdts0C3rr5Erp+cXmTwiCFWGhiJ
Yj8FcSfiXoqUOhm/+Rzitferrqj/pYcSQ4Xj5Y9FbnUqSHRYPloUtP5cIzj5RyzA
/9jw/8zqRGNwHRzabn31PJNnYpUOySlWLbRsq3+NbmRS7XL7IVwWFBIhMxxbqN8M
yFyuw/pluNVD0lHxTP/423GQ9h/q0Z2uB6ylS9eBi2MspZrxlAfmtTlvta/yAagU
5Hc3tt6sH9LSrQhC0C3rcgKae/bG9jjnW6V2ThnuddIK3Q4dBnZKq4YJE6doxOrZ
/AORDStkfqrX1Rk7c+QwpRlzojYyDbTU3nxqa8sVA4U7HqDRvfLLOKu7V4WtfxQ1
+lmVSW38fyJlyDvM5E+PSDZqDuJpEOnPca1J7CgWVKrn755S5efhns9O5k6rMGZG
KTK3YN1Ytbf1E6S+Vit92h4I/Ae4GrD/mX/PnBFEEfstLV5SU9pWIiKpt1WuWmSe
f97k64mrSHPUNoy1AMFhKxhceIrQfKjJvKHqc//sJCu6F7DRqO9MLIIirfRE4da4
GftMaoTjrB+FyuFj43783mMb5cRZAK4gBlD5A6L406KXZZtM9ZjIBCS7cyfSP1LR
7o7zA3cyhaTLeCizrp0MeB4URbSecAPOQxvssCpaAjJvxfH1rslXGFtUrPuKcQdD
F43Ed9c7m0/kDD2DT30P9RmtSI+PbIdTEsO5GDdAViq64ivzVzAwF7+W/JM9YpBU
e9tP/3gToyb6++q5Gm3/4u8FX0S1A30DtQj9YePSfXb/h+01G5F+Lc1GGoi1wEdU
+aJEC2HHT/8vDuWo+8HzpOyVfo1SNMmSr/XveY19Wyg6WS6XRtTj2sYZ2MDX45Zh
1IAcEOtLMIJDfLH4spiQIQsw2IAIzao6LT8SOdBTe9aolgYlQCO6y219HOKKKZ/Q
nG5LjGVtsitrJXmIzzshaKrfiSvK3jZ26XK0v2VNxhWhzVThysuR3ggpvw3BuQna
iTSG0Do0VVcs8O6pEP2tleIY27eLgiHU0iFnVaHk95exOjdJ0epdCaByKCel4A8e
kxJof/MzZiasb0JnLnWFsKATJZVa0m90uiMqep3ZffDcH0p7rJP+Hb8fLc0rR8l+
AsPUTNRJpCUTFnw/qnC065wCfsdrUV5vz9jTEcvw+XqPEoCwM+zPeNIIftlHbCWy
bU6fRvi+5N25/F1JA3LiWuO/qpGmU5t/Ad43zvq5E+Ql5acLqBGK6vrFyrCZDO3S
OeE8YM6TzF4SyojHlWqRp9jcfHuTkLKvXFd7/FUBVG26IvK6Fl5qwMNxEkbM0tut
DOwCimTQ8PP6p77VHVvuLTqYg5GK6ma82jvwspMrL2O5JS/Ue6qTrPa2Se5M1Hzx
jy8wNEp7BTsZvwAbKvqWjKbkre2FmjUAIK/3T7aFnbkhrBZlcQ6X/KgR508CPWuK
94uU0tEO+V8PkM8YmKVTl1iTH/F8ni2C0uRUZo43RmfJx9Up0ri+QV0M/PR9nVzp
JfGSRmUTApyzKX6M2VWn2pNMKJvORqxh1j6v2XOerKpgxhXszGR/ZHWsRzeK9eO8
S1Svh9exBNjgVb8KFRTcW45pl7ERO+DjrirtFw6uE6UeR6feKdOIt60v16BckO+y
umca9iBDEJq63fcImgBh0ImOaHlg8kn0a2/uwXnuKBOE/GVyWr6CDlUncftx2yIi
hpSFglC4EU5piVDV1LUYseEHtcHHyjm/4P7Tqz20yTcBdR0VbGwpkm6cJD6w81+Y
N78wmElUVeU8GMwXBIp0FMCgkVqob77st+0J+2C2u3qPMv5UZhfFEWzw/6hdfVZ6
21TXzjYiyOghCqw/P4r49qdDQM2bcbG8XFf9TQqRjW0jfxYqS0I2CMeeCw35KR8s
aJcuuiwTe585rEDcvFTc6ghwHd2BI4Ne0ynF3dI3ccSdMTCzznW9AoqsNeQrN6g+
53KhAQM+B09sfRU/OkbWV4ZZrYhagdht6BNfpihHNajNm4ADJmhJeBT14NYmFl0t
cTq/7meRqXDo/H6CMeMTr8+3DMt/t2Jags8RSQpDIDoAjJLTGN4rm65LgbMf9r0d
wdklejTNUTUOpVHNOJ+YPV2WBqAF7VJU0qPaCFkX//rhvlYh9qUdtzLGDN/pr7Wj
BZBquXBYDITc1AMaMJTbx3TuZgpJNFzyyx9nc1OExlNNiMJ0rFTgC3uM2rdHTCjL
iDruGt4wDs+dTaQsNUFoKYHabZbTEeIAuct0kM+LY1h44IFJVu4IqWh8h+RL3eRa
CA8zGRlKBwLD3IDFQ9JDve7NRtrqVlYBQgGQcdYDrs6xSzWUBzXEjmMyP4uXEw+t
lk2DHL9oGRSh1o2iaCixO+UYVS8una6HotuuNHnDBDrMTuUO27A3+Ct4s/h+ekwj
zvmp1eieAMhAU3cfAh4IixD+dF6U78RbKq30YOkXZM0p6r4rL9/lvyu4k9ywBD8t
ydRV4Qdd32xUFsxMyt4YBHeuC6PdUzhjh+B36IS5JEGkpOAYHzKk4pbAbPbxVMTE
TJlvIk8pRb9/FqpXvD06mvfRD361A5UyDNQWad3QQTQHIHN0C3n6m80q3fwLYAIk
YjTB4yUbCKOBUN/IFu0OEOBL0nxyfTydffwcu0SDwZPiqVxQl8xEqfiFZuZjOLsS
/9PNvHnBnHvZPVtjJ0Idm3liC49QFPxCy1LM9Z0EXbGqhW3HvNWkWvMVBxhtsrDP
nXOGSs43+dA5zMxfFnnAmsjeCNvjHfUMWn3GW4qtGRs4cxPHTzNqLzyp0LzJAd1j
MOkPXneIQw7D/JjtSo6cOykX0neStx/wuL5hwoaoXjk5rkSIhoSPSaK7cLXTQP0K
WjTIe6sEKGvuQJ1fTyGutCyoAzzo5GuDJQk9UdY+UVTfenTPXZTlQ6fK/QKlB/ar
kygokcni44DhffeJ0WCeT8FWQ37X6fYFpW+BC0WbBzkkiWlShF21EmtrzFoHavZv
oUaJtA5Pz8wt4WjC6gxyW1oWRHxpKbtvHzkehV97aobvzABZJlZQicHImOmoQG9f
uggvxyhhvZPG6O+kBtnoreCdwSR3AbXHV8fEzXLjFCtmTbBPlzcIsp7PVrGJlCqn
1K+a996jr/KVYLmYYMbQMuJj6rkXHPvis5tYr5HA8zhliiepr5rc+4oplP81+EYM
S/j2LnPCOcZEf1ky7drzVWRJd65oatXJt8MvRcvOJKukk2zfwzuoTU3ei0suX5i1
eSBi1CnA7CO+kNvOphvlbOwJw6GY84wcRAcVikGjSBnkUI/F5k/BFf7KmseqRPmK
vX5dQuJ0zQkhIInQOSaRHdgpqGMBSKJjpDrV4cWdJVUAwh1V+ttpnX8bcTIB2mQn
AViDQMFG22gPnUsYJVQ1RfEwYI0Pkwh6RRv59SzzBRvBlW6/FpCZXvopGA+e46Zn
ewESW9P46OWxbpVPT+dAOSQXE8XYcX0RLb4qXZj+NL0qZRsf0zPEreoirxmIF/mN
NiCuRnESjnfvJZylW8Gnatzwx6kY0VuXS7eiNqWSo0/eBP7lTdgzJ9PovHxmnjzI
9IBaSDa67HOlpSzMuzf9hGzwPzdtBw5JN+Gb381RZaSDrWDUW5DyaOd13Jr0PbzG
ic1xSVDC6fAOfI2tATcPg4zd/fJcY8ZQw5fcneePTOHQvm3nh+0YJsSD3hUXg1wH
SJc3J+REqkP/a0bmwy3k+Pj/fro8xxbiYgMl17TFkVWvWdIaVyA1s62Ug+RNeoLJ
6sTSMc5PKpyLLFqc7pveCaomGWPo3uzMdfqRppL+js9MQ0GzFhwXfiw+SzBdCEeJ
DTeE/n7Go5NI/awnNPBG5wG9yIZW9lIgpJD9fwd0n74C675eVuCPOblp+opkRJHv
1CVm0vb5eehdhdE1JL8iuIJQ293s+V00FB+5sH5VMZdZyH24YlvJK1YtlmLJUcqL
7rs86AusDmTm1fa7uV9keli1SPY/OMmGei3e22d6UQrRC69AkpIjXTxPjqPCQOoh
mO7cSRnBphgoAe1XhWB5qZtWN3kaUpGECK4Jbwl3TCgRHHoNdvMokAUoAxPqffa5
Jy6HP9xlno+x/uddD0ZyyX/Jm8Q20FSTsSx9xv/IEyI/kxgYPZUFNQWGsaSTkWau
b9PCxl0jE3jCEnbJXY3HhQiSNlTtqWvn8vBgdz6bZWvPs64HkjzUAxW8oYRfwauD
M2NwQ/3M8rA3StzVr/5doVrRBugt0vC7YZXtJEgNp+3dlrYuBsiwad4THY0sCJ/i
f9zQxN/L6h6pK6TX8i6XYAYDqUHeQLatG3/JOsHoNfIUw1AEUxD88WKL1n8YDqyX
zYXtQoUQryPHHx6mbwj2S2o2l34lqbpd37ubvmm7J1t8T1SA1SNMkAhV6E4EbRrw
78CaoEGo5U+qv9U3ok9ieM+mjWRf+ZAxX6e8cdGkLJZvcW7TB9BVLcCvH/iqr65U
SAYItQVCom07VvTC2rxrLOu8cQact7oPP/3//r6KhUl47ATsujeGY45UoQhEdBqu
mt3iqJ9l8UHxXR110Z1J9V8AOgZDchO4G+LucS4Dqf7JDc1rdeOe/QxEwY8uNXYb
jsAVUbyGu0N52q0kS83S54RR+v5JtzkLHCCs1JyU27L2n3BqjbdNvk7Bsvoyt7TK
WEYPxsreweiNLaNsaho9KAd7Ze4T/+tUuAxFI+Rj1ODDhqS1Eg+ijA77d0knn8Im
YjNdeO0ut7YNykxFpMTAgMyOIQmI7Gw/wFWfKoxfwiFOx13/ZBUWQxEKlwE6ckHE
8xPsUFeRuR0URchgSE7vmHlZUW4V/6YRXtDmRfUGBrdDpELcYW/l81+6EX1bbN47
Kg1jvtY8QjP0UL1z25y5fnJX5lyn9emBJ3OuW2qKMvf7sRZd+7SQY/jZe58gg0/1
wXV+uRfJIlv4BKrMl12v+XvmM6LGSaAH94wPFyfRaV1kx5mRDndcjUzJNHUnpTCw
iaGu/JHKPoISxkvPwRN+N8kb9chgyqN4Q5YNFCTdObN72Jggx4yp4X6Amm1otT/S
XAeyHnh8AGf7ALa3qHsnYMVmDpKrpd+R2N/HGUYyRHMN8yxQ7tmGE0k3bFXqYLWt
G6uzR8pZkScfHOVti3naKhpab9btzqn2TKf8I8LwCqThScSlzR2SIe3O3ALrbqY6
BpXGwZvktt2AffemTpBjdsK1o0wwnDk7Djl4TGN3fZSQruKdCNJ/m9FQSnwdPrRH
J36p2bYt8UoV75euQzIMSn1tPoZDAMJRl0yKFui5Cn9V54q2vx+XBeJkcCzrhJuH
O+Ar+xvhi/IARONVmNw/i5+tN9640uX+trhIfyjbmxeDa/ywbevxNV8MrwGJ+X6f
OkAioQM5nXmqrJ1KGiYHtgeqad5n3dE0Cp+KknRObO9qQiKMQDxBA1L40RvPFXM7
DiviRWRyWPyDOPjcdvr7IALK+fkjhnBAPCWeF3qYnCuwrSEpBGBYyZEZofZtIM6V
7Ww8u0pRySxGU/eGyAClJ593h9runmPg58GTaBSmknpGwSEh8NSDvOxPjyGzQIXo
tWbBfH2BX9YFD1q9wOf6nqPUiJIvFDqEwuZkEd2yIwZ3b9eqpNTisI7rZWyCs7Oq
qzIXr7cL/LhqbbModJHPEmwOvLGdR3CgNSMa6THi1mXqHfch5Ap4qIoRFZfEOU0U
jKmBD0OdqLOSMut+AEzUTeOHPBeypLEOaf+wd/my00qZ8KIMb5M3tgvgnLG7jsEE
s6rcF2ZgGM02ul4DqstNLY8vSZCP+wiYAovM6BhIXLOCt94c9LgCquZ+Nb1RNfSJ
idDSZ1vzZMNEf4TgQZCKy519KPLxuKcLS06BLImlkhhXkjCeCnckhVTJ2+WOPepx
yc8VpYtu67mj7VLPmY1mh7U4Sxo3+Tog9ZGfYOvnHSewaufen1x/RneSlM7eklay
vK+aiwXm1TVylcNYbWkbyinx3xYtcYGMtNWdoclBJ/l6tKQoPxLJVD4VgFXOsqmF
ulgDDYnqcydhCWKnzAIG4L01erWVuxI6yq4A2K/Od9Qyh6rHMNCFkuJ86fSbyx6n
z6HrMHOrtiTbty8+8JYfw46ofSw4Ur4Dhejoo3dl9a6ErZ/Ys1Siu8+xVlEroE6K
jt5SLzZA3gW/i/PcXtWtmTV+5A/L25a03RuXJwt+fbvBUDDI4hN8E8SU+BWaAjLQ
bWTGiQpltJbEM3Ll9oOks71A54Td/GyWUMKyoDRqkfBGn32UhzJDNiZOARO/c2P+
h/kvIzzfBRz3bNGxB4gg1s3+EAxIiyO/u83bmeqwuGsLQpviMPoUAqcnZGt44+xK
V2bzLSDM7J22Plfk0JDafBXGDpzKZQ5D9QjjLNlw/pOqqWHLfJkk4e7pna5zKD4v
cj6FP3uB1kGys/+uouhckDr24r2lbx/yYicugj1lqQ3QvmIuq3VLDF7tlG0r/tRa
8kCQ7hrNUga9KOFtuehe8fxNRP6MM0RIxh/WVa9/5E7zOqe0B6kIuOeJS0T6Duwh
+qZ+CWh7PlmjcvVVjQqwfhuDkJl+BVrMg5zNCtSjndq3IGzdy/4wUJCmfhawxIG8
rz54mcQIQZVoZocWmLbF0OHtwzBo8vUK/1cHxh6lCwaTy+VMqX4wBXWkrp489aAw
FvyRjjYnVTi9yVC255Vn5oL0gzYSWc8X1D6ySd7JppLy1vLZRLP+EUOowz/0G9oZ
jox0phj+TM/SCth8tW80RPqycHgW8bD8tG5pQQcxorV0Z65fQGluAaDIVQBx7DGj
iTR87zq72mRDOe8QjArsiqkgHv8YP4kBRZlZ1hewO+ZGW7mlxmnUCWe9FQIoKzUF
R04nwAglZl92+0ojahcjPSkN8LuPC+sa8cPwd+MuCNtzPLyHtTsCj/MO7eTQM1yl
9+ds9fS22TajV7pcf/oki/ctxPzhbBdn/h3Y+f8SowRGKO1D6sPG+r5JHveTopkA
PmiTGEnT34LbRNGz4CFA0SdSW02S6kl946ckKevOdg4iEL5RWahVCXT+g88OCBwu
MPkspGMixXREOWpcrQpaFav7p+L9SjCbEdrk3gKKmYeQlnqangjncUxi0EJ6b5ix
oQcNZgP948GwLg97ORsiRJldZqLHJesnxIZ24INuZHVwRXre7qfV4kMxa/c4+FD/
49dSiYUJjb6r2yBA8jzfI6BeZeQZUkClrh4v4ISHD6QTAXA0FEMkdPgytObfB6Dx
7Urw/ID0SbIsBPM2aW7Kvt1J4x7qAJ2FvhClW+fCkaKA73NowXSHNXtligEpxWL9
XPZ1HV/Pq2MZFz66A7qoirPnkbNROoVUzzk71QVqflEaESBW6MsYG7jjCi7Py62Z
MCY2tzx5ON/uqwrayKkFSeMvZBZYdlCSSPADd5SyHjGnUQ/oIukxgUPkE7XdGyl7
AjJkwlXBmZx9YtKJMEiCbMXbmw9YsWmXDWHB/urSogznZBnyGQj+2OFykhyY3mNx
0yRB7/F7Gc6NPKbQA35Rd61dKcHZYrpq8wIkIw+WzYVmZ++9h6qcAVb7idku8w3L
gbnuHoFWI4XE8jM5hpcio6zPxfwjaXivMv270eUT64JW53Myw1ZUaYZApsQ2rrNO
jcCZXa7NAgsJdJGyRd/x8v1A5IbsILiZD5Yew3bIrH1F1P6te7EaKQHjKgyqng/+
2S7cVJ4lkWIS/YEEF8RmDRxUhFz95VMlhKZ/KjjQxcvd83UlOVUwm/kJjdS5njWg
lLSIZsFoYgUEu7Gmu9Sww186G5iu10gQhDp2JXRmJQQ4rFEKKxgQX4a0xbqZCyFI
PwpvgOXFPMjVDhLhNpG3AiuGRBfptYXLiTTj/nRaC5Pht63qCCnkZ/n8K4z97FZ8
Riry1nrlAJru2sFL8wTtdmJpHJ8GuYzXRuzpy/meev/P0pqY+2Pq8xvJl7JBTcNp
YusUpl4diep7Bqt1AQ/CD8CAVNijLlRoF7UaooiLessquvS2L9L0npq1aGHFNq1M
RCD1ZreI1AQvm0hDO/rmiY/GFG/WhdShdnPToakadPDksi4wD0fQ18uyd83mQjLP
+dDdp3t9+wzAS8CCdKpQ6tbr5JCFvss2fnFxIyJKkDpMG0mQjP1+Ns3lzepPVDd4
vi8m7ABwWv4Llp2WrA47inYpwSVmYzRJGIpXQDgtpusC+uhuarn2KFUs+tTrRWgI
NYu0c74/d+V6M4MBsyNgC8T8vRPfHkbEXavgUBbXg5QD0o+NKEbkc7GmXKqsXb4E
Q86f+8jViiOEi0w8n4n9r9M1hB0U6PkPaUs6KulBZDfiGqD+VgbQlMQ8HkyLK2uX
ElAUtdBApUy9SJEK8MPRE6meMSGUVG4cCQhFN/vfDwtR0qkeiUFo6PffOBIF8Mf1
m8hSKQAGEihUZhrwjm3v9nUP8qIsmTPIeYndirhUQyPHy7qkqXdTaOZIhEwwEO1v
3cMjQpjOYaDWQqQuqhRNy9QfjkZ9ozDpm7k0nEPEsxfqIGCsmkBV8Ax0soUssXKY
egbm/5MmXYettxY3BCJQKzfyTCnSf8Ltgt1I/QLz72bKlZ0FMmelKoyWfRoCxcMf
h3z2MbrDoXhgfljc54unE+8Z4E14LNfOcR2vhGlJg75UT1ZYpY6j5C6lw9+f6e4w
Hlx9MT57fqTpdnYcH6Blwn1OsR55W4d8dUBKuEwFF4T25TFaXXkrwy3a+qSyOStY
oCYXyRo8ifY4YhCkI6C85hKKblOWoiFLGwLeLOs3p1p9uUdEtTt6c+eKgOUOPT84
oY7wsY2/sJCReyX44xkfzD4+Ug1GehmhrQG3pADS5BcVKoMQOzKaBvwty8+F2eq5
Y4XvN/rahYr18Za7Ad2ZLb5zuQ/5R+i+RaDQ2y/2UI3r/29dIwuQBcsMOogU6SRR
4gwpnsgkQJWM5l1D0SbV83ZsmT4pAe/LLWlkVf51MMoK/84Tf7c43GOnM7+e8+Ts
e6g7N4VkRJKxa2s0y2Lkkn3aCg30NjXJIHBCjJArE8kcvLBo+DLzdhn3yK0K2Q0R
v6NeXeFHvs3TvHPyNxo67YGSuQExDifnveUP699GwmdT+sTdkbuSVC/U8IlboQxk
kV12GPnCbN3Wv1Dfcun2thdsRpqILMXd+4kjcOIFxPyP67goJ/slxDaHH+LYKsrB
8sozupLphS/Nvt+Oot79BKaCJJ7N4YcFaxG0jGBsbCRteS32AGFl2S8SkW2vsARP
BpsjhceNvCNJ+7x0zQJ1LvqOqxGPhIC6ci1+wrGhjG8d2cyzAf22NcTWFkE6RvJa
/gf0rZOOU2yGUkWjMlgvTu1bvChSPI16a8Dr3yfBjb/VG4wjOP72LitCUAby5aRJ
9kFux6rBjuPd2XAYEwhbwAPD0C33OqZQ/M4kdgn5q7OSjCd+KAltMWUk4UE95dXU
/QN4uxUKMyPXiJwt5j8btvuUj5bz1kKHwBA+GNIeazq6u3hd0VbnY5OBKqGF9tpz
3dQbjk3+qo4WaJgIQQalISG9JV0kbOcuPctHElXdZmQrvPiBT84h0uWKHCj46cDd
y+57yRDgIp+su0FrIaxr4eENZYmDmZhbSvH0Q6Vi/dlvDh2PNdUCFa8C68HRURJ9
DidhdVcc4tuia/zaRvHxf/urkGU2uUSEw6D44f7fqxrynZi8BWuEsud/jTXVbjQi
2JxuZIT1wcCUGBPwSsDOfxgzibL3hKV027Gvn0IXkLQklbVDRhoyKh7DdoTpFKKC
DeBxXP3tfgfH7khw9vk4x3zXgsuoiSIEvKMe8+CfD2wfF1b3+w6KD0QagqEzFto1
QLGw8Ki0nzx2B/HEySWrQvIfXNMKi9avEg5LNf2vKS98amqKBKB+5VtAlMSqeumX
ybbKg06QVTH3EgAoUZj9KauGD03YPMnh8QKNbbfZ2KVLOzntrh1Lx4FdaEs1kH5A
khMhMiOOZnFKx697jof83SkzT1DTuPV6sMPPrbuQ3SBFLT0pw+mHeS0AZlbVdrJr
yidPojSu3c78SUrdmhOME/pmiVwFVwlZ7IvltutD85ZHHC7yUG7aZeXdltt+lA8M
Zd0OuXtyrvId2ckbFiaYu0BycNRN/9n+ZsoNYpa+HkkPmGSzhSarelG9I5hRSwt+
nUvwVuXP8O/CoZTlbPrqli0C0yGqDWyU3DQuItt5+ml5HoVf08VCGxiOKaMY3KVa
7OMRtA0QjKHKGa7r2nUj2PMI3Fk7y9fg6sVs+WLiC4W89+DDLgB/35jkLphWrreT
gjCagphV5Tv7QBxqNsJb/kyJzAuP5IdnB4F/rVXWHEGKGfFp9FQbYBrkFp9kyEPq
V8YvqEgvYfWthmfYlldXLBFPW2BY/tgG0AkR1qYDR2qKknjv2wK2AdDypi8zMeSh
1LQ9qug8BkJztJ1uPMnRNv+1o/wZ0D45QPeQibMDIn4Kc4D7beNqcHA36CynK3Bv
PfAQRdyyJwWfQ2oDL2bPNIv7+jhZARHIBfBA/eihqcju9lULrd6tGLyLQlem1Tns
6SQdjYlD0Otiu2xgBzm9F4yr8j5OLQ4lBvDCkxPIYigsZX6F2jbjj1nfhwdrHBSP
fjSrjREsufTbl5fFWXEOdGA8+c/5VN6vJJOrQTfny/M+addvmR4Q8d55ew7yyBN8
EKGYBmsKA0NlPDHmzXjToE6VaV+DlTCLxSZlevTfTEdmQDQe7Y7vRcDEh0fa8C4X
rKTGTVgRKH5rtacZmtih3dNc/v4FPsJ+kiXRAjqzeMGny+BBDsUZZr0bYQh0YDwf
HIUpXD08pp4Z+MYAMmFItr1VlGvxEku1Mtw8FPBl3V3LP3SzeadTVIsZ9ovmZ1Gt
gCUdUYQoGKJ6SHtVUQTrorg1EQgE0ZYvkR+2po2a2VmBH+hENIuxzuQ386+CnG19
fUdWDev7tbZxcsjBpS9a5B5uZv3k/CTD0OJiXXaj/VcgoBkM1ctUAM7YtLGL5FWX
fmyiRmfVTu/OQFuqfBkIOksKGwRFMw9YAEDUrlq/U5Bqe0R6KPfVrC+qD5jBtdD7
1hKrJ39Ko9Fgq+KxKdN/h0wqI6IT0wRnzlONPXJ/svlmNW/0kB2SRmqxET9VuICs
5HSqfMVaw3vrZlbf7q/Knj3SCUPPvrlWRFcMjk9DklNP5h5XW11DrZ3RCA/t+bUT
toSBGy2lnX2YAEoEPNhLsEcc8MUMIdopXQ6zd2W9QlzmRbreozePfWCjy0GwOlTu
0OHEiiB/6wtsh35rlgFW/YAt/Nx18nnv+/kpuOep9vzJpb0HtgT/VEideoyLPtGi
FgvIu6nSqS8A5TqTgZDpmBjAg1lpuid1q9bSAJLkoRObVmpiTnSSJBXEgWIF55ty
bzWhxzgPEfWGIdcq0LpHXDN7hoTigkaqdrBXr89osYYYqwCkChiXdh5Irtm4jnQo
cEOvY2KpePs1lxaWamo4O0JcIDRz8t9VFeahWqhT/r7P6v3XdY0W4FJcOcSgz4nU
LcSLdbnOATAK0lcvbZ6AoAegk/2e5Hp+5Kwyo9aQP1mhjUYl+6b4gzgd/jSmq4Nl
YKrYhBa/bjPmHqq5vBwk4ow6udvVybkNNorjiHqBpeqU8euGFn1UJdyKSwXibhLs
UI9l+l9Ei2UJiD9AH+9uQOGpY4kyCXv4AqWqdhn+x38jvKgt7BWHn4YyWipqm53Q
fNaQ8RIomZPVnxLtlF/bvLCKLVMLynFgCdpXhWwtJLdEmjOqQHjhKr0PF/n3C+rc
z52PBbNKoCLUPMd47Z5Esdhyl96w6ZHBLhLW+f7UbYHaCyJHEJcAVncOsy4cSsWS
x+LfmP6ra1JFbt/ZCkMLOon0OHYm9muoejJdyyMFjuU4Q/KoduuYIIY4PU/EZLsb
Mysv/RbCugiC5yv4u8WpVsc6f2QV/pvfkQYhCVF+KAzGNEtFQ4MUDA4DyIv6QyEg
qtqZP7XcoTqUyb3EqX0sBc36M+HhxEt5SKulKuJmZ8DjNJzY9pnNFpQxNiOfFPn7
l5kqupOWsioLgD1GiEGCkGKDmXr2crNVIX+Reuv53wpc++E+TYCS+d04XTnBSVXC
qB/d+x+Y1Wv83T17vw1SOqOivv48A5N4HFXI7cmly5WQSiVFE4HmCK93EqpHCNpQ
KdNEDdRO5Aun+jchd3X5e44zoZ9MHnVdXFKiBIpyZyatjcwvbMLWgeVvUIXWRDmO
navcFFV9G6Y87rMp4ZRBFgusxbWSjWk6sHiZoJYxjOwdi3KZyeaVkmE161aR3GTh
zpqDfIAVdu3EtLMEeleVKzqf8jEY6MiYc+8GQgQUelJxcDeJiD+NZXrxbLqFA+1i
1ar/+m8gUijlBjXAuVQHpH0mQy2TMXiYdgXFvbLjuQ8Cd4EwvMv2wiKTof4jZNty
isv/BIv0JSo2OLXbsn/A+sh0rY8IOu2+hUda+MFathotO1QyWXNy95Vaff+exx5N
yylja0ZfHuCMAh/zFUsFtJeZCnJZR++lJUsEuT8LMp7omRdU+ff+5zXDZJErE+LS
IqVYjWfNuWOyrYi9bX3pmLh6ZNKgXY5pLU+QuzfufxpuzGGyJ31x06JJ+ng84hx3
sVLnSOBpc7rp7+SVjFI06zTUSPLL5ZKzhL0zw7ewYz+W0oXUTSaffJqFcpMj7q9q
hM8etXzVoVVPyuEUQgwaHRRkW3XuJdLZIxEn1lZUcnSz2Fk0KrP6K2JZQj/t9A3j
I0FsnLqac10DO/Lu4GvfxFxgVTbrMQROuNwFdQlyyXOmZR6drkJI+V1LiYJquSba
ZXGWcajXqRnDAfh72ue6dib7KGaHKg1OqEICdu6LxjxTfZ0OroeM86jJnJrzMYWs
kX24sz3KNdK9UR9msWOL3je3moM9b+LZh9O8oHf2JmaSAFFR4lJMbtM+hgIDt+bu
6Srr5sl3JuvsS3qPt9XhUtyMjKrKzMUs0fomzQysWL+x0WQyCe7mgfkwtYobY99K
Hg8NBK7orz4aEaq+ZIBi1ZQ5pl2cUJGodJynPoALOG869CW3PQ8UNfo9o2xjb/1A
xJkaHPZXeVUJz9W28uo3N3SAIbfqb+25J7ZxmgIAEWo1URIwgc7JyXIxgtmM83Qa
aH5vh4kOfSaZFNUe0ZVhuP0S6mHn4fi3M7LuszvkOiwwGZ3z3FwdKa83U9qq36G0
Qb8OZsR5H2cZIwWJSNp5OG1azBdeQ6Rzeh3onTwVM7ZG1MsUyiZdYlHB5Bp14wNB
4hv0jyghYXmjEDO99qKLYgxbcSGcAW12eLvdS4wDqRoB5HBz5FiEshSw/SpV0NlP
dUBPCgexYh9j429IcFgevirf+jzfhlBOeXrZSwTvT4OtXFLJKRoEriUdTC31PC8A
JloPwcylXjzXzAEw5Ez5elhjIyZ6020+PrwIVSF31h750lqnYNgBDHsA26Q/4z1Z
ftcvqXP0mTnGGJOfc1hXbiRX99LJLGqiPPkD17wncrlN62MMmJPWNKn/ZhaYxk6s
8tETqOoDPrMXXgFIRgV4r9hUhG2F+/PUDsv6KHRo+QXM+yRyQMLja5q48ZeIkoEW
i3Yn2SFY/HWC5K1UgCT2DUjqS0IXxrCFbCbfPoOku81dZoGjHg/jrtfeoEQIQjSq
yiNz0vYOa3PCvEgI0cS7GHFoqmChPC5CsZ7JuyN/WBz7ZWyZS/aMC4jLv+vvDD1o
j7jZ8gC2Vhqm/fgPjv9d3CFbNitdRcM4pGU20+TGfGXN5YNzmq6QeYf1tTmq4aJq
p5LpAx7H4gYl4eEC6uYM//cfNS/n0XeZTJu8y3UC+2qZQIQwfLNwJ6IHPSsDlFYt
FJZGdbv47ytuRKeeTAAM7fQ2xBwJcrzLh/yuPNdvt8KkgjGkE1Scv1p1QjmAGoQF
7LEbYOyXHZ+YJFDEuw2p55hAsdw4h/drWLhI9vE8B2nCsOwx/M2JdTOkI/R4VMc8
k1ueHubq9tpV9t7w8pKop6iw83HMXLFcvY5u4u2nyONOd7ymdwpK2j81dfn3K4rU
JqGuIZncF+N21BgvsQGAUA3ZxQTaZJ+McrpZkJdOVXJNcPZQI2vns9Ko/pURJUjs
8Jy7h1IELpxe2gGAS/IYHLwj2NkxMvI1NWIMsJEiRwvvy44dD3DH0JMxftdZybcw
CYp126Lmw6Bu5ZHgyKGWkXGdMDs60MV+c9BzJOc+xTGcJ/A0LX7smUqqHkBp2TXe
k8x6mKgppALAj5ZCgexyo/j3Mw3ctXqSFKK7WZ4v09/+FhoTldMa0oOH0WUrvK0V
eFcqKCnj+1j3kckYaLw08uvp8KUthBX4+uqbMd2DMRafC4YIyC8aOxXgeONUaKvK
ruMQlYAqBT+FZzWOhvTb9/Qosfy0Zv36HhtSTbeP2Be2npgGtpzb5ntdaNV5Tx+T
KgSL733iY1aEQgkcQETM79tq2MbGEiIKUcWchrFu1oqp3Foj82ZL0XbLoX0NEhAS
AhGcXEI8ke7qkdsjFTaNPuk6WP0G7sVV6xMFzqLteO2eu6/EYvgCuz0Twbo4SRa6
g6oM0JGKhxO86nnamf0VyZQdt7y+kO41GmDSqfSgNZNSN01XQ74hUbPEj5BUP37m
lxw5aT5+lan6PwyK7ZGWaMVMEB8kO1BrVW3ydeUyrOUOJY63o48RPEn7Z53HIbIU
4T2JkqLJMZxMv7cwCe4eY3HvmALBzr0mbh/TVPQAVaca9hERGSFmy3hjoGdkTT6U
UloqoItWRJXTG7yicZ91d3vkNLj7O8j9vRked+LLpNwJMsTm2ceg9cfFEFNh/bnJ
AuuorvW+ZhsH+uA9v2HZTafN6YwEGi762NYp9uTGa/adBJBAI3Et3XKSvpuDFL+F
63+9+D/hbf6Hjg0sVwM2uKGONeODBaj+EefbHPKR6KyyxAZh1l+rkmMfUR1IofgN
3kvvq4hVx9L8+0J58URTAx5ExNdLP6/mfkOghkebsMRcHFyJCSiAnvi67YrMurW6
QBgNmiaoH4yG8oWMvvBqMKleRs1+G/+Wd2+BklD32wg9GXI8PIxcqchDJPdTqaBj
e7ba1jaGFbEa/Eg1jUKfGbJDbKxO4SkGwmB2KhYGWBlRerFRUHQ8zFDzHLAmc8ua
O9Tb8PcE8s47vSf8f4N5U834fLWdiXKHbXRW0BgvTCcj1hrY5qg1MwAL+7rsBg61
uYyBG05ubE5iUJdT6Wu1lPpYi4C0jGfXHA9qLAZOKwaNTDNSGxk4z3aRK+Pb5SnO
r6TMAtt8FyNnRLRZCzyaYXhj0Hl0g6YAl+PRTOQmoHwB6IRKxBINmKAL50btKatM
Ivcp18xPKE0wemXOnKNRJ6JFdMIIEc0UuwGpdAa6rRexA9DkYseGNce0r9bHeymv
PvY0eRlUseupHK9WrvytOVWiaw8InfTU9I+Boypnw5cH+tTIW5HFFvmWM6OGdCR8
7vGyMm1weulZn4hpI1pfQCHODuduN5phSIuo2mc9pBF3RpfcOW0lHA8RZa8Mi+3S
xVBLgRkFyJk7Dlaa+kLt3g7gsuIyLbPNQigC1bwBZpMBw5rgbvt4NQzViscXudRn
9Tzph/93JyOkE6AOWSmCpSnL/i7rxBCQ72AeASWRihzRg0gU7NFFCoPqM2Q02LUf
zWMNWW/6OB/SXosshijex6iDr8+0+iDu0vDbJwGMaIKCZ+uiw6rk6CiC6cfvvNin
yZ9MNPcmEa4BclWjhkKICZ/BOXiEmW3Pig01SYKZ8Fb/3cbHFHXIspGYBqxdOvzW
yzP8iYffwPJx1HipWwFA593M1wZEsLsWnJFAXZzC6MC70knspmWZteeAIeIxDgky
5FayEDDD3GLsm17+EHyUwzBmEVM8DkkIIU9lHfIvDzNeIla2qOdxHzGU5/CF0ugD
pzDbRV2/Vo649RUvJCVmmUklTeS2jUO18xdwc/WdnDtlOJgCSUzTzv2Vt+4yMlQZ
YHIgUlJyj6Q4lFbMYzdsCRB3zjLE10rknV1f4i1EyFnzIBEbbv8hZ72U+tgIlZmj
6gjM9xblPRnR9NHLKlRq0mcK82ZPQqf43gZJ35RLu5nf8LH4U9FOp+2YIKS+vqev
HgpTaEokV2RnlQ35PW1noBX3mIBTj0qSOFXpi+mRVQzBIFbLL3NjjCILpuj+8NTH
jvZzBY28ILQCveqt0RAotqq8qvNUNXtPwHOX5/0OCB23jdQg5eozuX0CVV83F13r
C/TF5255WlopFIH+hkf9zAh6C8EE2F85cL/gztlHK7C2V9ChMnw5bqguUTZSyi2N
fsTayH7reqgJIz7EWOqO6+yjOf+lLajKz69Y76oA3XhGviZaz9JearYxn5QBnxAF
ubTpSBZ49zZF0n47SSV5+M4ZQp5lyOOl98y5bKg/t50eNlgZ/Vge1O5XB9lvVsgc
675eRzqdBPiwPpfXFRmuMjzI8sLf6rijiHZJbhyihYLuu8Q1qXKvj8Cfq1WmG7Bd
XFpzW9SLfQbx4AMV2zF8if3Ii83yUDin7msZy7edzaY+0qu+DDvxwD4uMPRnNw+1
AOUskoIVz+FK6I/JMBCQ1eoX232yjCGelhLmH7U++Gf6kJ/K2lq0V07Xurj+59cb
JzBF/7S8sjql2QGoW1ekeb2RFmmde24O/aYblFmtMKFiFFlTGXBOZeV2yp13wb2K
Gt6VyHE5k3LGbDu9eNkkW9BjhMkoj/9wcwkovwERKqBkAi+3Bma20coP6WZLbTsb
LxfsSADAfmHBeliE7jsWuo3fW7SXB5ZQjiqPwZM61tIwXUSx4bmtmbgRc9cM7Lzr
P27KzmBNDV98z2WzgePQXXZpvORaUzlpjrD67F0KGg/PNoc72WWqa5JMX4Y0iJ5X
ZcQs6MG0RfZhJG8i975A9c1uZ1OvmUz/aDt1z3Gv8PHqDljXRk1TLOTvkMv66o/+
B7CTruaVB/k6rR0Sy9zy0I89uOKDZ0zGXusUukdhc+OgtHKqHgnUKLsZbK1BRaM8
3hIPPFx80C0HQVbeF5p/tXVlkU19Emc85jOqrRaNp6PaIPxGoe12UPoKP6FUOeKU
DaHC1TIlEGDJHKIDUDuAGLs82J9qGPahQcHXzb6QSHyMf9wYa4D3XL3WKdibFsmJ
cXjcuDe1xIHOvc1j8fxkM7qeHykn7vrUVJV/B8J29L8mKYHriIOmKP0UFhGyOdu4
gaKFnOHblXz9Ni0/hB/1csjyAG0OgLUofYvyKz84vBi/Tqzm0ngehpgrIPKCHXY8
j1TOe85OJwbAjtsXeO8tBDznZjpUbSmt0YaXUNXE+ysY2ZJNnKNH1boYzo0iQBI6
WFp2+cwdkZeKpxXvirZcRaRkfOBCnbkljHv1cBbEg6oiUj1170IgAos3z2uXfIZy
8gPCln3avPJvAgIsTTXzXgNe5ubBgjm6bvqgRzGSa5HRJC91yfZEtePc3NekC0u+
LFWLCcFSIS9Md2pzGZ1f+c5MCqdEQ5sozvFWGH0bTujqvDbX2PF+y/V4T7OC5Ktg
3mUyI4TWCxjI/AlsbZFynxRPoY6Lnm8x5uv9eAcB9Wi8uqhFqYRM+HTxRihtJ1uy
EBG7f2m3+W0axoTkwfRtXoo8FtrVePJKkXYLKyC5BmvlvXPseFerzi9stJqT1BdE
RrnUmUSw+eBE7yVjv8fjyCNRYrHCWFNPMdO1vg8MHLw2t5z2tOV8GhIHgqSxb87Z
y/MwzQT1BHUn2lXpgC30UiFwpQB6f+UuCNVewDLYyy8dF+VKdOnlyaUUL7y6iNso
b7eVYm+jmsQTcQbpYxYGLB0XIq/PYenx3bd2Fnp5+KN5AVTKudAE5mycWZv31O8q
wOQ88KblG6Tm+gWDZVeIKwUbx3S9id66bKD7Ber2cQJWQz8pSLyQRnDi2iYn7x9H
VLMJCGBQJ/CQcBFOrgSOydcuMTPKXfF0I1kqNV+RUaZdAwIw+B4m4TLHm5UTMFZ4
93qLvvGZzLhooYPNFfxyOvtnhBkr2H7vKvCaE+kayXmkA7HER5/4mFOitMdeR29r
JYtP0s2AM/XIy4hbRyZFjLC3zWLvVy0Jcau4A/Jy3UciYQjGTGzzieYg+hhZnlaK
UHxjBAqU1adDflj9L+XKoY+kSgC3LQSvK7HfzEZCI8JARWxbPi1GYU5rkgybRNo6
NXC+yY1SqaVl5zAHfaeFT44YzYpURcifkAFHoxcymsG5H+Ze2JcFDOZNazutExDu
EWXwDH26W8dk8EI42Cp1UIjP1Q43iDeMhnOdPXCL5xRCGJsH/wYCwE7lMhxBPTlC
KEgPZQEK3scRq06hECVNEcUr4D5MQOZaJ+HxqJewPvbR5MzAKm4FCXRb9pRgnVvP
yKHJ3w1M/Jrp5O+apSuPkWfWZ5MzfRZHkwaaufaGGsgkUn0hJEQql6PE5UlC2POv
f0tE5aWd+XnlswGz2XA8dEdbuqN+rNCvVGdQEJ4vCKgm/7AQ/UYytsfcqsDsogi2
y4gCWkNTsKZMp+FVEXno7Q33Df3kKBeHUPLZBwzXv/gr0Ha5sc19rlHWR5TPahwz
2WyeTpHeLwnun2hOivwBvmNmZJoCg+tFNgH7P4Bz/75lYElT5Fc89+9/m7ZXd/Gs
2fOL3ujXDJ7YAU3MBYHfwbGOTIdBkDTQ+nPF8CJN3pc86LZALyWPU6PsWgAmxZIG
9DfqBIPo8vLN9K6nqJWdqFrhlID4X+LR/kG5cBRiqhkATPOsUN0ry1HO5jKhI7Ty
qKeVffbuv9porH3F+4l94V2oIIhO5p5W9O9HX4Butdj66a3v+E4sYY64QUR9DJi7
0p4eR5cXENGuw1M9Iulo3XOEE+f85ASCied1DtvYAGQeZYtiYYVFZBL2zqI/tGT2
k6FEtdaPMnq6KTTnCYw2XiSgdfn30A5csTziYC1ovyqM69uYK27vGy6muRlKhfAj
xu2T9lFwpXrloAP0zQh+COiodhx2ontl+O8Lm1mqubzwVBCUHg86Gf4sfxpukRqZ
OpxifJB+RA3PXTXkeUuUitZtGkZXgOeK/dDlJRsAsjhWJPo17lq8WD9WNIoD9HMg
DywNuT8WtDGGThS7DrlCzJQaoPCum8m1zgsilSQzQkkF5k4Dv9JnWErv17c9AY0s
gFizuasLpmhT+3V6Uxe7QfnQOFNcwB1fjlH4qxBMac3BIZ2MuwNHOs0VmcVUA6Jr
NYOeD5pHdLOvlzvtVemr0IFzLXLXB86i61xSpK7U3dI6l8Z56zYrLw3buLKN4MZq
xQ4iiHouy+XNtWw6ztoqfhDSNBjZwpdPA5SIl6doFWT9CS150RjwYojQH1ss0vxW
OBbeeipW7XMhH2HcU897ce6xqnlrtcR+04Q2pG9prTZb9zE6PXWBeuXAc0BcCPE0
0m4sCCwYYxKRtDnNJcuP+2QwoEx7vr6D1qcyKEwyHFL1P2YqmzohuaDYgpgCB0Qz
4X9lOVrg66GmRJD+YD/lZhIL2LPRiurrT/aO5/ldLZZZeaZ080zZJfvnXXO25gB2
T8dySBiupCnJazhbovNj/AeSveC9w8YP+lpJYQq4EMBk1USm4efNAXssgXjJOpHu
WUbzd6K/Ywmu9w5ARQDiLSEwveAyzBo1vJgkUhM3N+HaBwDM8q7UIbNlVdk++j8f
DB8THmmihKqlchAfgp+FIcK+g2d02NRz5Klrt5d/oT6yXkErz4zcHlDefXQuMnre
G3HjkJGDYqu29Q3Nm5MWcxnE0OBVWKECAjFBHFtA6latTjyXwymH1cWt1VrGcR1x
uaAzdAGiRI2zzeZcGeCKwO7cFJK1AVNvGtjolX4h68+6kbnZnY/9Bi1AnstShDrR
aWA/DD+7CJRxlo/JmwP7pOlhhc08j4nCum4D/4+qphhAr4gjiiFKVLRZ+d00OOG0
UkpLcKcNdki0XWG9+1MRupCznm/pQJbIZLYMC2q9fpQmtRciw7+1Sy11hTMyG9wp
MKOlQUTSYlE72EaaY31bu7LaRbQlZP/gUpYxVRi9/agPiXMjfc/GxrTkhQg3dhBh
6vIdCVnSPEgovnV0adyaKQeXIX7Qczv8S1esvrVApl6DjcSv7ZcYZQEndnmYQukS
mo2fARdaAlCDnk1wGNfcHMif0KS5dtqg/SfdkYaVF45jl5KzMNNBQqgvnFjQ33hC
vCAbIOPo2lDrtLbMHtT8qoGcxo7QCKzj4BKqTe8JGoq67GXrJvR8WbKujmFAFWNx
EeKjwXAkqJ2Cp8kL2l8ksxGycqE4nMw+CTRiSq0yLDmLe/EsPktCPtPEYo5QdYgA
LJEPIjTAlPFyFpSidVCURZLr92lUb0rSJQIIj7UGmeA3eR52fOcTDPzZMMyDuZJw
dBu1BL7nn2ZVxtuEgKsKqwO19AW9+cp9+eOghr1yYIXEp8ZkUm/rZ28RPCmQ8d0r
PszUs8WS8R0WIXn+E36zPCY0/PQpZiuijk/JomQ8t941YUHRbdUpufBy1p06H4dq
/1GJdBAGfMvhrx+orf+pETDwZqUAlj4kI4pbff1XwtbeBiTVyw2sv6e1Z88Ikw+I
i/yuHqapQXa4rN0G3bY/OiVE82T7UfxISijcPVgdGt0pNb5nq5qrZZFOY79HQ4Pp
7APf6/FxNBNAn50XBuGDtJiL92BnepdfBUPDSX38RVGPXup3HVlZNR6XjFplY/EO
Gd41nu78THh6yeLIWwwuzu/+KFFcDnfzPIrsIRGSRMORhwOw9+1OH0KC2J4L8OEX
dgl6LEBx1wt6uqJxk+q6uiE6+5/rf4UZnqSCCboxTbXcVXahTgRpTVskdjyOQqme
2H5BV0odRCF1MoetcnKSeV8vRPYn3p1ACUl6IuJ9Oc6Ps29np+6y+YPsjlh7EphU
Txk6mcMa71Wq+CMQogex5C6MzcqktZxa9ZQk27CPm+/AJq2M86kmyY8XP4Om1xGt
t9kkJvtcds1p+Z50oxj4nkr5on8/MAz2bpdgblq1xBlC89c4deIV6BmR9IqZ8NoH
mZDacfXrqipgv4HkzZKi9+Cuf/vx1KPS8gzTpSHxuRnDK1KRG6lOVYD4pW3TMHhU
zfinkKFPi0SnaNOebPJT1YNSgr7c2g8eDMXZ5oC9pF+GCrVhAZWI9c6/ZmIVw3tv
2AkOdFzslbFirdLuthayBf8Pmu552J/IwPnhLMuyf1jLT+iyy2qYRlIhhHJwoN1y
XxwdjEQtP+XLENaPjrX91C54oBVBKWjhE1YUwVOjgMCsRZDtSBxiMr0SSWs/JiKJ
8l5eIObHh7sVKDou5essTM49fz4fylf4e1ioguYhhYWalGKH0BRSVsh+k92B0v0H
zsTz3Snz+pvD5seyPhR8l+7B3Ax+9nI/R5xn8iKADgTojJXN5+5TZHUHruQjmmyq
bceWWfxhqNFZTeAjcPR0v+6xU8tOj1bkubQSxwYXe1BFmJ+rCAnb+ziDwhwdrk44
IsFwgrcBHQXs+9XCLppSspkGZKYUwPW4XbSMTdLt/tmY+UhxFnB8Qn0oYT7sp5Kv
QXLVCx/kXnX6SjdH3yCM1ZJ5AjcvC6JnmLU6d4CpUFKFlr7MImpxG8pBp+tzkjp7
ZJaBHaol+uqtIGYPo5UYZkbUeiqJgsasLoFza9zp6HFdr9uM6kzQq0p2yAHOqHGA
G2Hs92bjEkiyWDuPwZMdG+0Hx/W87YmWUjWbd6ai6kmRUe7MVHWbfB1ejUB1BPO5
3K2DGWFcnkvc6cLPrAbz6q8Le3HslrrLvoR6nsK9P7hanmbQF7ofszZFF0RIfUWZ
BK9Wn3DK6SHgbys6uqm62/SmTQf/w9+bIhg7FXvHzDwIG7yL/eTmsTutVglq0dSD
bep+YG34Th1qaQ8y8uAoBUkXcT4xeQDg0u3eoLr9ri+0XXXDVLZwBmweHyOZqjGF
maXG9a1f15vw2yAMiQoLdDpSxPRi+DQmcG+b/NDlzned8NynpGEq2+GFUBzLKlDR
je+nk6ZyhryUg8CHVc1QluEnz2Yhb/6nc97F800GW3AHVsFpRiHfY9lId5ms2tYv
JT8XHSRtrIpWiT92oC4wtbq8EP9L3t1sZjJixktOg90wnSTBnl7rK7yUwGJCFc+J
pepX2r1TZq1oE88qN+diYzoSb8kJqsqr8NEexDziY5JufOO0j+/QrsmmZ6NFf6ws
bUBzNOgMdIJMrcXkAF4jbDPP3PCfYa6lEmr1oD/ydPAh/JckyS1TDoa3mvaLISxo
SbT1AIqceGrjKEvkFiGUoH4GOslrQsEbxh1k7U3H6AWuvEHmB8DaLUb78PYAJ7EV
AnJ30oK2ZVjZMjTP5F455vGdCLMxuU6wjoqk3k1wJ8yKNHhEJkKfe6QzRKC99IX3
VpyaWdc5e6BG8BpZ8U32ZYSoVXwCbYs82hm1axOOXR3MhfCatuYxvo89WsKG2jfv
GBohoOk64Zt7u+8hbvJJV81dHc4bfSdWZXWIQ4faRwQ82d+wuRbAHucAu+Xxhb9U
ChjH7E6o7SNg3n/Aj7euZX77/bxn19+PSxROY1DKMBG2yxdAqqFVVmtFn/1eo5ze
UWZvMLzVgpKtOfz7Ddk0A5qERFP7am0gMBns/medGg7zil7adF+8PvhuJ3JTFOP4
C084+SejFIRgGtMqHdN+mv6poyqXnKk6PT4LLBTRYTLroPMJMqonY9iADP2IonJo
P5J+Ts2VLGK5wxitSy2+jyACn3imR5uB0TrwHeXspraHRUTyoAcWDaF9k9GZp81L
/m4jvWGzUqAfeWGghI9YIUtpZWn4pNwkvAK6z8vQt+GyS8JAGID9l9jOIt4ePD42
klk4axXIAMTAlUaSXC04LXUK7YhcmVcXQnDyWXRhfhLTALHm9nVM9slwa/Rp+XsU
X7Wy6XLEHCs9MIAVo63w6CAY5CWVpWHceGExhB7bA/I/cVdX1tgGuBOz7flbPjyR
/+mft2R+LtEJeqhRWkZivkiYdgPVQeu2hfsXPJEUItrFBMlKuStf3iflaf0Eulw8
J8QijVjpr9TZMbO6OAntLw9RjIrZwnqXR2UQzneT9n2P/E8AyW6WLp1IYUZg65ru
DutIdCcuDgdaRIdRI9p1o3NpWrqHK26uhw96R/Wz7K70TjDFqtesPTCtRle3vgn/
E3DYKFvLaQVHqHAoMY5cEmQUWElxBunHuQ8Lq6M6G26atRgI+m55n6D5T5PxIzdr
IBbKkcaUHwPhZ70UT3PcTTbzaUpA7SoptXa3KMyZJEW/VbS2fOfrS/w2OGCe0Mqd
NkkH/u4+9Mhlp3skLq+f6+XMzWbStMmTOSpIhbKZWnvd/77jH088aAfbgBABrCiK
PINTBkF9A2BEgj5YUajbwwwJb7sGOP4AmH2qXbQmu9fvyN2oNHWf7+1SjxpLEc9C
1UcLaBqKeXMOH04X8toxLFDeGQDs1GCBovoKAX6XqnhvwIm+b4C8v5yN/mUZqfa4
QfPA483rBtDr7fW1iCK1gActWZDJQij0t4qrfT3S79QN/5lQynd45/0H2SOOEpqn
FdB+pM+e6atzu9NArxBr3Nb92plJKQZvn2gsEnNkL9jYA1fMHJqSdr3mwR7Lgn1c
BZq+C/QfJQJ8pqc93VN/cffxEXq+hUFRWUx6nZRkbVm0kO1BbplXk6KHAHeTXmAS
81ZVJCVkVxDZgsI2TtWQeXYdPJ7FQYTbHIIB5Mj5Xl8XC+gW3yVr6BEtsWiQpAuk
LN8Dekh+oYifTK8X8VW6pORLo+HEdLHEh0P15HPrf1Q4Kp+zHPRPWtwvxbgRYf+x
twIqOzKuHLgj2SyDl0zAaTwuWRp77o+MsDkVuV51hDkWjAE9AgkYXIDe6deAhASs
jsm8DL6jmbiIfttRM8Ep+/1H5ySS0jzwtWQjDhsz2etvQ7U7xhV+tKDGoqQhI5nt
+v19ZZdnmdhxwiDpGWdK9UnOreM4i/5oNO0yMHuJGd1s28zyCJCmzXkZ36DptzXY
AFrSh7yrazx974GOTptVwyv1r/xLRuLxwjympkUunw/saNQW4T4HgqKpTKpgK1yR
lGijBCgcYFbIdhOtVytEQ/PxK3++FxQ0qwGvLebOKx7wSib+Dh6C+CNFR76tw0Yd
9+R54ZSHnGYQ4O5P6SRQxLD/6R9HBLs7Zur+mW4mF2mIfTLpKRwRqVDHw/G7LNIF
YVV2Z22aCKswjY3b5cR1Xepe2w6bYe5x9+0jgDwyZP2XWuRQtucAlVUhHu000scs
wXe5/K5cNJ/7CMbonp0JP0LksU1IqPHVFiMWaDpNsu3hAiIqAKKzvZ3idro+5Wjl
sSsRcp8zBywQVenDXvcmqhmWYGAiCO9WI8YrCCRkZiBhSwDodlbHCcrOaE8+9QfE
gypAFXvxLc9PM0iF15GbeKTcdyq+pEp2prO3qMH+1CUJSvyANwBeOCCs0YYxsiZA
dYopzft2B5Frx8I/MaXkeD3S7dkvqHRv/l6tWQaVcNOH1u+m8oE00H2pKsGrZCsX
SBqdPEd7VPnwESwkNZR/4AzbN1T/Fmfi2pbEeECRy/PRiDev1U7nk5JAvFv3V//K
lWROWDLs7Erk50I9szU4TfWs79VOiciy3GFxTY8dSyBgkLA4vdAgkMEO5iLbaCEk
uQEdPsLy9Jdt8ej5tTLk/gWKse8zPWCIQY7urHOO4H/HLh6XH9jpK5/5tkJhiFsE
G6BRn3h6YADOPkjqTwY7PtXVxf/DilwG9bDE73We2czTxBCA2KER/NtwiW6soLaK
cnsEspIvLq68nTeeHd5U3LxWR/vu7HcpNuyaceLkJwZOKBYmN4e9N5D03iIKhkFD
lyuk51pj/cq9bPYZdmzUmsdO7oqr3cT3BbdmMm2T7bFT4yj7uExG33NIotPbdqAY
crIYYtRjAPhF1CKurcpCm4Ojq2FTvNWiUFFMZrIsDiBNWdbboRVMJgcqy83G2u7N
cljMuFeqnOiqbep1//gjws12I2SvocYD6PSXzcdQ/4CO7f/XASicAEJ7F2PjZb7Q
d+sR4DqA20L17t7zllacB0O3j0O7bjqqaVhg1oyhHHnL+VjWaf+HS4yWQDwYa58N
VnFNmyeX7yLiXFF2lelj+0wKzUuZ6t0UCgZAalTiFwQluNZBsWcVVmvY+qEryuB/
acCtB2PGWfh0f+8gJFgLxaFd24J2nZS5rb1cMMCD7305VO40o1aaaffc8iWwmSbJ
4zR82VbMXMS4pb3v8MizEZMBkxiUFWeP+RMtCQgsHEHK1MzTjZuMceoC27WW5PAS
1fb/JKsd80uAehZDEEeNaREkWQ24NjWjOQlL3NJGuE2gJUiNtqZBi5xHcxxTHmKx
1Hf1vB2IfYA7sAKdwRZx6wsUbaNGaQLZADyhs8ptkB78/YvuwKGhYJJFs6d5fIMR
Sj95ht/PuU1Bei/4BZrQSAtr58Q+4Zskd6mr983diR+5r44PvheH2utCF3HUv9UF
BEZGDWwGJUUY833FjoXDAAhAOL7l90NXXTaf4wWSSIydMaPYkYzcScO3ntK91AKh
beQDKZZXiCzpZbTQHzY0xlQmTamNVZzLuOVJExfcDxoNqFyEC4/kB1hjAvmh1vfC
ILfCXAN1UYHaM7xwUti0Ug0S64JmwUYvJ1MEQItBNYS3/2WyjepV1d9DTSQ7lOqz
0x0S6l3mBQWbeeeMF8/h+/2t5nc5j886z1MPq2rQyrAxXbHiZiJ9RkHPduAs5T7S
me1xM7So6SdyHZeqO3dAJGfvYLKzKJ+uVXqwGSFQRCBAEZ2gbLjjZpQBl8rSg8rR
Urqml5exi0C3Du0A9ynuFGJdeySsuTe+Ab0FDFoCtKpt8cUht9oO1MFz08ZyIaKK
CumJ2XHqhUXkY6MaZlnUW+3w9uzcxnh3IFJgVEXxhEd8UdlTh1K6hL//cmZSGKrC
ulAwneE950r8/yx6mNHfhYo1aQNT7nc+Lqxl4EcWUmykRQ9St994U9v6P4ENR3sP
5kpWBio+2gWxiKWxiR6Mg0H2phZCiz+r9euVhWqG6SnNlhBeHw4i8HgmweZy9A1g
StEdzw/zTRyjAW0dt3wVSLEakzTV6nFpETk6UhUrFB1DqS45SEAfoARmQWknz1y5
5aOs1m0wu9s2C7CqlaAUwW9By2/GELw0uDgxbJsQb6wC4967ACq/fb80sSG3GbRy
q2NVqtDPuRZfuw4UrmpssSf4FMfqgWEZv4A4q/nrJjK5cXuQWNQs/LXQPySGtJG0
gOtbSM8v6zkzadnMN8ghUeUEn7K1MJVDTVQp8gRCD5WqCQ9JKGdV/mYxafAtBSvC
YAIgLUnKqqnffB5M+DoX07n2bD9jodmmXdo3rf8MJSzmZlyeaFXs7g1Qvilph51g
c/rtTLJ3gWlkBIRrp87OIJc2UEduzzb4ihrmfGw6KBuXBe0BF0Sl26R+i0CvxyY3
NsmAHH7tXNZbnZFsmD8e+QZERr1NCRbRGf4ugevOhZKoTDB/QOz5t2J0MTsXZmoc
YwiM63CngRwbsX0LXBlqMBjGB6eN/64SCGZtO6YGCfb5isbObrXt+dslBGrgXw5r
oDA6hfzcPhIZD+H9b04w0TKrtIlq5DSJhz3nFveCbc7okDK8hVd8Tt0F0LXM8jWc
EZVBTi/RvIt2lDGe52DGAtd3UeMRi2oXFnkuaNQ0TnoAukzkPgkl95WivfCKyH46
wykN38VxODJYAuWu1GJrphgW1ggBO85CwxHZMD8VyxQ0Yc+ylo0eyfl8l8gZVSPP
rDxrOhB3tJlIIkmgzplPpFR4xULYcT1aPPPqnKlzk56EjIfmspnGYBICJC0gXKaw
GAFps/TfjfLEs5KQ16CM+jqnLIYebO8DAdezqtBwOaxSmNvrlFHREE+YsbfSDBBH
42jkSiuW4qLRP6bSFVeTbOwMyuI5UnJ7BNAEvXVSQEjhizH0/2kQr8x+0BcnLblK
JXT9NLAUpkrN5K7GQtA712YnpLpUo+Rn1lrO7mPNtweqFBElOu0kpkU/7RjyyFxY
G+r/l97ADLORy3v84uEi6F55TmRN8NH0qfbIubV1K99JpXtDC3lcpx77YruqZ0OJ
p/8mnG4BJZd1qbyh+Cjuwg2R98xI+4nOIBUw1KP0pE7+SS2iQt9Y4q+yNYViMHNT
oIraU789cL2xSRR+y0uPQjfSrpvGLUq+7eQWB457JT6PQJMjRl5zC0t1HXBeLJzg
CSXL455yR4RH+k1niSJl4dSygT6YZr5KaVj3lcJJCvoiyZQS2Q1Zf4n8TiDiAU4I
bErlFZzZMO6zPmdCiI5fYT4zBr/1Pgw/qEFTmScMgWeyhgMfNBL9d0dFmRx58yLC
gE+lS449n17W6BMVY7j+iNM87l0UHh+PW5LVhzDQkcxgVksL60e56N6IT/i0r7Ra
OL5/oMqi1SChbbVpY+qLV6bYmrNY5NYP4xbntxQUejTL/7yI6i4Dg+HPfgpTMhD2
j0oA0wESOKYoJNhK9kpyjO/wEhsNa8SJVasFH+lTvCCKth5dZbYsXqkVvr7ol5gk
jBwCzKnegzDLAiopknHRgLvZWxckRnmfGCmBh3J6FJOya4DFT2rDt6b3IcYtpWBB
Mf0ewlXzjLF0DVnoCEf8KZAQ7zY1FcqS6fSrAMzwCkJXXKWrfn6qoY7yH7HbIE4t
xk7+Ae3m8eu3y0+i7RXJQOz6R0j28uYwwswWolTpKLCU8TouX9rhED34024QS4pu
X864NWb6ihWKFH5OAV3OS3DeYmCyid0nvhD0d8OF0DWHqjSCFo9z1WFvau70LKGb
Yab/zrDeRuSfAP0P27c//SoFlGisJUZTrFQGk4DLKZWRtiQILXkV+jb2hLk9s7PB
dZQi1yZFZBTvrmc9qsG9J6SxKaDhszjpCajaFL/7QlCxuOqCl7e2PxAOmYIgK9Dn
KBCNbNH3QR6CjIltMygkLs1Nd3ExNoS6A9b1B8CWYHvZ07kyY8rQShgnYcS+FaWS
4EDHSGHyrep98PkYw8E14Gwihzm1wSsxeA9c0kqepfPmQfolcJcY/WHey3vF+nKc
t9yOy/AOT4K+XGAFJvUrNCuxAJXOiCDvNPWhEpYUXErkMFEvzuVHG2iWvvoPYoA1
OsB+YVFZ+5TJG65GD+C7OIatYzD81Bs7+PTpcScUbNnQLwG/zqh/35elXZa0HMZY
nvtOYJIwvHjJ23VTKBtBU3AIyKB12aWtdaM/5bPLWnCJeVhTwE3g+AgtLoWLwJn+
h+t/TVspWNOFXewpShEtYynKFy9VVQWnqkfmAppnH5itZ0QhHIEGpeSVKhwtMxNV
G+cUGWOzen9Nr/rkqvU0pCB+werH4zCYpRgBUSfZd+JzN5CLyPKpwUpS16U9NG4f
B9S156d8b/Ml6GLkeycV0dVWZrAdNSPDsiBZICCC3cvPg7Oq5pfYhuP4VieXt/yL
31ryXZ25YtmBhy2fbqaFtKJIb3/swXrYuCnNOReUmdre14jC7X25Yrl+J6wtFApU
iZAjCxbMq93i9tCJjLd7LHhPzfW290pr/ympUriuuoJKap39rJQP5BaOYl2fkz5t
6UAJIbH+5vkmriQWk6QSBuCQHnWq6HOhXpCwQ9V+UKxtyz7cSq4tRRQoRyGyp72U
3//O3qAyaS6nMI7YpVVwViAe453crtEE7A2x3LRFg3PDiEOqlj7vZHavVvaVHJ8Y
9ovtognSL5tOBt/4Qs72aoMjITVbONfsRzm+mbDVHks6l8b//AckbUPWfVp+RZjK
Z4ifVg1lYWH/EMru107rnMbX5AaGY61qk/xyd68okAAEKvYAm5nHGQVB9CnR/hKm
34hs5pwmv6VRmUEh+OAPRV9ulpb5OGEa1kUNfWPUPHTxOOCr6+GC14sIMVFiFw5B
R0yYwdVL+1AoNAMNBx+yUxSVefki4+PSdmO3MlYPyo8M3V8wkpQkUHkkuruXG2Kb
GMdkXMqpucCuQBmtoQHMIwS0aXuQ3hl/udjhZR7WpsPv/FBwr03gfbI7/sOqy6Pd
A73zW1lLhhQtte/LtQxSPqKfm1kjVK5/rhVD/O9onjjD6Js3z9aO5JasMfXqKir2
ckan6tjnYa0s/znrit5ZutQFSvIR7GkWbM1yQcWYtzaXR5ELCHAhBZehmTdzoH76
/YNTuomkX4HoMBfLvM1dRuYUHuUE0SqTn94V5qxvsykdE73bAAjbNaNrCnHFlu39
YtcMAVTuRZY7MCFSdcnV850b33zGMqkxsrCxpL1ubwRBSC7kh40S/qn5h04QnBck
F5NefwOHwIdAohAs9W+/J50B42jRm5BgKN3ElieZ318G8Qjikt8QLr3KjfWRYPij
IoUPMVC6S8/7KPUZsVGZPndetv5HtIZ3WtRFGL+TFGCNtxHOec5lNXzA6Wm2VVx3
p1W/R6V+xAvkmW4T2/Ywr1m/0wkS/Mr8RQXlcnG6mSeyXIOEg3el6mvVkKcDdogP
S7sF4VyCpNm6BOQVGl7NH+wuDX5SluDzl/3O1da1EA5hjTPvJh00k6LYGntibXr4
M4gqBfFsDsnOw0FcfBDVaMng3OFpqMpggqolEayOG29LPJEmdOBKz3bOvaHvgEQ3
BsvZjmKhstkUA5BrmU5TQwByYtvcyDl0Z+bHYixFZKuXejV409NtaC+DLDlipOqo
TGXQAl5vxJcK06VoRdh0gnso/PkQfAvqJ5ZqCQ4v5518aOsvVFim7rmRNYzU/0ee
247A5JjcCt/Hz6pG6jwhDujcHDHDqdKL0z+Ju/8TE7vIglY3BOilf6+mWOZs2Jjv
dXLTWcl60WGZ/EON5uQA2HQRg+AHnGCKnguUAcX73Ct6pMIDuH8d7BoU0ZVPAZRh
fZDV1Jyj7rvl2TDjYIiUQsCx6pD7JBuN/paGiulfIWjkA7o7vmh+efdtIjzNafqp
tgXsdyRXM13M/NbYSNCOFWsLAlmdl0zZxxh0Nm2BsOTaD4hymi30cy7VI1exH/er
ggpbFF3Bm3hdpquBkObCVb0sf9igvQmDv9Ev+5Ii4cmjjWoybkBp4K96/02Sk4JA
vPPkl8NqHjAbEhukQLLGfGjSAtVGXQZxij7hPbOOGei0vSWbNIeSZphpYUw9Fj3V
row7NYvlPvrpB3qSSfRQshO/aablcel35hxuR+k1Qlu2eWlXLPysv3Sq6mCDew25
rZ4jht2KMgpmLVj0/rfuEehC7r2P3mC8UVtnrrrz+qk2+7X3/soVhAmebdVfD/y0
RmId+LnlR2lhR3ZJIDq50R7uejoTI30xw1n7P25u4gvOtAHJpvA4/dxM4fkyyKLt
jrCzfP2o4LAS/KFHx1YvretJMYTwWvTm8FbcwqAI6uB+E2+RZMeK0yuNzEOydREI
UcQhm6uL67E2iqCZNlwOVdAhVxmlYjaagVVAabQ/J/J/nEl80TMwA7qrqWK+gF8D
NU5+vSiMPZWcphcr16YnFYh9ONDMuUFBSfHlWgr4FKc5eiPXXtVj65a1RqCNAIIM
1t1kkYQLBngQVWPUyI1KHr1jescUB1g3iMd+HiZwHZ/FRUwKjiohnSq7AE3aat7/
VqcrK3XllHtP7JE8Mi3QJZxLVURnDTvoCWs9spc3Gx3DkwyRevZbfnTIbs2dhucy
UvdDoJ6HaZd5PCtyYeaw/CMyF9WeUa4rCu5LGYwBoYBfRo8lJn91htPPZRnp+pIL
8Lsr93wkTqN6JW18FEFeHgtXymT9H+bvPq2TzG7BXYwi4nx7Oi2B5AYQ/a2sVeog
IbuP7gcm2d9vKdw06zMVGY8uPTkMplxfWhGT3Y0Bj9caux0D3kzYfLlwoBnI26Yl
+biYksGFrincaTJqDvjJunlolYVvQyyyBM++p6cgJcw9zmjllbPtdCkFw34Ase9n
R4v++klRPuW/cCSoCgDJysFwfbiSdECfbc/wQqqYNPK+H7JjFy+QsxoSlXO3Jjps
xZZ6L+Iz6bgqJn4yWsTsOph+6rfFxV5zfOFhY/gWzhmqiDM6m3MO4k4K5z+8cQO1
IY2GsKLCnk62vAsiYfK1qn7LMlzYTt1JKU+QktqzaoVVdTKmUgomnCPuO9dFYgn7
xzM+Bkn3+YGEPA0HIyV6P40HQilMwh2ZM7bYAlicTUsLc1glCd8cH0ZnR4x7Fy8e
tgNNQq3eTcU2aBpXcdus2wg9Sc668ArKV/Dx30rjd4GNeA658guYb4S8w6KVgnGN
z0QUT9QbOCRm3MXGKK/xK3ShWtb6B2qzvU3uwlr1OcQAwqb1unQchXFbbVhlVzVO
FGczrYQHS1tzz6r2zw0bHcsBK/MasIh7i4hYDr6c1Ky+opBP6CDH4f/cyUf+qS4K
HjMDnlRLPNajTvy+iIXkuouS5tzgwXdo2/M3kXCJn9g2d+MR4PGQHQPffOE/gWca
OF9wSeCWl+4kPBmdoEQM0cJvlCUUywWbW2yI+dcfYx2YdXVzooW5w69b4XRxDSMg
WFrgb5xeMWp7u1IQEM9hQ3lbNHRQktvns57mjGVY16RU4BkZLRY1jwx1plVmFwRG
pV0FRR8Hq4J2N1qJqgCUJexCAGKRPNjQii6nrp/uqQ+S7fWBo/Wm/BoVctGRZ717
eH1+H1z4ovfaWaWnobMYlwu5bPd6DU2+4cP5PX1J0woDJc8w26VzLmKOLEcyPY6Y
RToiJvrFXk9zkTC0Ab33RdfS2kvTvqGG4H2DliWP9ZQ33e51KdC8gsobmjcll4Bv
SK/JTL41vb6/sD40C5FeL6yQf23RXUWpwSMcMZWjPMkEzzoQ+Wto0r+bcKj/lCdA
37nROoqyV7mtRxgEsaMo122M+Zs+djtDoyFrTZ7tjkupMqSE0Awd+tXtBd/l5hVn
H1iyweY0ejavqHZFg22unAdBYtas3dRYqE+PlHiZ+4f5jLC0NXdenOSOl5jzHuXt
mFZqagnGjLcf6wGmdXzMadHUHHwrdbUUmpU8UnKSRYGD/vuM8Wadtq1BugLNSYMf
Y28b9igNgWCo3rhE77HhwLefh2bjviIqaV8WcUYngDfcnehjcGq6JknveRxrgeea
bNAFDfdAaiJGEFCFCR5FJLT0MK9IuHGcpGA3+xD3KSh/GIQ7UgHeTYw/+U4dq/Es
oUtcimavlraduUHIVxdV6fF5QkpCsyEdaebWrYzwKoT5dAUIt/jGkS14Xe3dakes
uio3ziakunpfEr5A3VcdKUD3XIklS1gJk5UXorE1WwOKA3IaBfEJPUO3htNbHRy0
pG4zl9OzYX9HVrWnWKBxq1SVn1nctVEoVuYSZ0UaR9xvPWQxT6ouLEgGa6LJjQen
VR7ByNQ3Ej1/x3qaXAjWqz7LFYyPAx08Lyt1dJzBJ8hpBlX9H/8kfArGSEWnjFFR
D7OvtfrqmK/CbnINR3QxwXivG7eNMOah92kTlVmvzb4NWwFPAojC0r9g0BnmrSJv
QCWOwBypPzVpXV0ri1elsaRb1xjr5Y0xDb4shD60fg+JMI9p5E1PpXPM7DwY/ZTP
vDD3Fa0d0c8kIY+wu7r2ynEjy1fshXTswB15yH82Bk62KTSvefW5WqV5xvh09i1I
EcKIJWE23TjarmKS1jR60kP6/lgZz1cRgrR/v+5dNy7GmrL1J6rYJeOGfqcCzZ5c
5+yhMk5bFmQKrQjM0DqXdAloRj7fnwJ6pQwP3InxKQNzXw3Pjeq6UE2o2WePK1q5
5Ut4pEG3fZiQcRbVT7kjVCZQN7s6U6o+Vqa9cWIREw6XVgihI3Al5OLOt6wwJfbo
AV+fQ1WZxFMVm8R7i60CrrmVycNVjeDxE6KNz2A63m9DUhHVs00x3TyfZs9JLO4j
Eo7eUblwW4VXI4z8LQ8wHX9E8qeLsNXoSJ2wC4JzkmxlXKVoY9XB6AAtjM30b3DX
bC4pL6yzMH/wdh4eAxQuRj/hlloJk33AZfxyQ6KW4EyD20YsbJ0X+I2J9O0h878K
ijv9wUpg3iiAA8dVCGpZ8Sdg8B62wOf0pIIo2tK8lwZZIsCMPg/aBt7TafzZmC8S
Vpsha7yymX+rppmKuCTGhbMR5FfktLtBBjMKtNMEk9vScBaWw8/SM3b/tipHwBjq
jzrE+TQO0f6Ld+Yl2Mh3qrLZdh3ntDdcOliUXQzse6iBrC7L0iFhNCWvk+c6OC4T
dAnL5jroCFtqSkY2YDgM4nt+ZfGkwd4y0/NKTGjCT4ZXcyHFQBZAkJ7ck18aVu74
MlxBvpW57xz12+GJw9iE85BXYdNMxIZJh42uGXmwKp7ZKMiqvrCCdmoH/jSriD0S
bxGdX9M0cL4w3IKUv9v61xpV/rQWOTrlAovDw7RAWNzoA8KzqEym1s8h696JJM96
poklJRnnbtFf0h/gKIG+CrwaGzaeOcxANECtW4/+ZsGsf5b8NgfEBOPG3Z2f9vZa
1FgwL4v25SCyLRxC/kpErmJye+wBGNkBs1axMogRn/OzFcvq4g1kgCr2oIPQW4W3
rsNEEnISZ2pvJ6prKoFHXluKr33eWl3U27D74sJ6bYxzcuyO0K8/KYBNhvBxI71W
v1y/PpATjY7bJIpnIv1iFT91dKR9KHGb1n7sMPIrOsb71TGTn/KR9HqXAsKAax3K
9xhqAzmWXyiNpwQ77Y/Gpo7D2/GyxjGZKMwvDlVqtsD8d2jelmV7XjafR+Y4hJ7Y
l3vmWy5PTON1qwNQSR6Q7CgWKu8YhjYXZ8yDeAsJwL6tHoI+xwu05uvJetMxSAXm
Njt1NwFTPovlBqa6gFO5pExgO/+SbMxsCtVLQGjVnH33BDomDgxFKq0R9CgTl+0L
uhhcyotPvZvAW3qTY2LftpJCvhJCQ1CnD6dBL/n4dpF4a/AOUU2q4lGIBnL2y93H
3Zf5RlVGkmrxXDL/DLNclEoy1gLPpQYwEehlLAwOU227/+zZH354AQCijv/Oc37g
ckWWlsYKTsAc66qNZlmoGu8wRso7fjvbiThh7H7qhfkm6l8Cs84Wd7n0Phi49bka
7iFOhSOdFFVPHwxBk86B3j7DLzJ2vY8+EH7vQ+Pn1eWW1hm+KeIRRfNU65mF1imH
3Z31NXLsK8inzak9JiZyhh+j9n2rO/sjRZLF7v1jI3h2DwSObbKUv/NSqKRAtInQ
xf7xKG2gku5Clkm26k0+lZZdB9CJR1C3N3DdsSSwT6YQIQnPXG/dOnuzcbUZRtZJ
ww9xIE5/WbYWZXKSG9Xr9d4RucUrQdz7dMoflP93BgI47ON6pryLcCpUnLy1YnCW
ZR2TwxXHYB3PJGbNPsRtRL10aDL9VommSfz3bDa4036rbzSbivPSqjDHTqyxeaj4
jffrrsUbzO565EG0oQ2+4ghz/XGyp4OEJPsHp8+S6uQQvAV2DEM1X2Y04NSHlXAe
ni1SJOLugjDOxN1pLTKt3PLBLgC+rjk30+r2NaOkYHpfb1n/Aa4Axbww4ZxGulBd
Nm27mPgHxvJvPykue4iOuY9mUOH3jS0PRsWx4QLaInFAKc0yo+5kSfluZpLZzHKa
P5kpCXNXDH+3Svwub72+SFYuX9B4JFnE8N1KtFtb4AXhQPatRHhLWccK5+fyLV+p
9Ihj4C3RQknePjELnuE3BzEW+z2+6kvlyR2Sw0uH1EQ7LjQUjm8wr1oJG/yPccbJ
Ry9thpXRwAAHjR47eJuJG+tNiur7tjTg/QckCLA4ltPC6dMvKayXNluxTqG+912I
pEK3q5DMrag/gjexLUNR3F+AIwlJxhJMxWoMTkRYLv6qmtd30PvxLL/D6A7X1luM
li7hSQj9KLNv3+jwBIv9yzcSPX5v7gU6ywOsizf4Evds9M/rBi+jVRlCz0FfENgp
06TqfoIw6tWyZsNXMR9NuBLIgxiwuTLJzqH3EnVKUkrpDDa71rc6FpZJgYkFsO5X
YKcdnt04OgQX92uX1UmBqd2oADoiPnS3dvB5tM/BSG1fs7diiC88L1ovLsLVSqOi
CSIY3z0I6tgsF10jyzmjE+Fvlc3hnWUSpYJaRj7AwNeh9jhO+wsmc160HePGGr1S
lBtxKpdg0eKKYSYTjJZkhd/sAavQEzL3WuIiGxxWTG6jcQ9//JjhoIgMx0di1S3Z
TzN7U8zQ968uWn9H2zg4cnkPVfuYijRpMXwPaSToMRMYqKZLXewiEStJAWklNEl1
nwnd8YCxjMcZe8Mnm4ihLTBjOH56xbVdH3Qs8dqvL4owZ3BngS7OT4rPcAdpWp9g
5ekXEUVZ9gL2ZJQa/TCmPtFrI9po9LoAC6qBMNoYywDAO4p1Z1GKoqNMPW7HJrA7
cv2Y+VKZ4fv/os0H2To1yLv50XMY6FybL5Uwza8W6i/s9qyl2bpGvrWtUH+b3oJg
/NyX3kp72ZSHiujMd0bVgH7U4+o27XeK2n/0cVmEkbGfNMsYUd48rh1hDbp19daQ
dIg+pP+fx+ntF+JDQrfXkxVOn5OXzRsiTLdQG27vqcPhYLJ1PCUBILnhN/OMgDXM
GaRLCWP1feiw5lPugWjtihrlxAw4pf8xP7h3xF8oAqhWxAz/XjywqyLJs85FZfZ4
0JXwitQ618RUCOwcEXVdGZUUsRNCCulOBw44bS7ZCAdcix/ZcZ606a89PSu4XNAk
aMWOyhML7xakAFgYneOmPQHUEEsVM79fZj1t/DmV1ed3LjRU2yUg0u73C+rwRApD
8O6sIEjn6KoVet5fbsbwJtJXkO+JqZk1gCMFwVJaFjxgOSp52+aeWgonRWxxFjCy
XkhWWqOVnKpJtw9GtZM33ks1E/JWjEUg59oEdoI+JWQCScLV45sS6Khg0LvESWHA
VkO3BxGsmAHtInH7iW3VzTJZV9O+UvE36/hSFugtSj9ja3Oqqdq3P3RVCnY1rX8j
72DjW/Z94MkHlBW/VrIpH8Ao5estqa9rzrz8PwsPRWpNdmOd5026l4rbq46cShA5
25cirXH+1Kn2Z7OfgcunIJcOd1txZhtrwEUkGxUrolNcwhjMhyplwCAoSvTu6wla
GC5JSca3n8yAcptBcYQjyKZTa2ho/f9l65sjp/wfbFxzXd7s8zRpd2fe3v4jcRfx
RMfYMxMXZLCDQf6qeEv25NckTpiCEIEKaMkktvFEPfVCaFvxYp8IO/xnwpyXUmj5
uNWG6azBMbX+vssDsB4mWAFHvcdypZB3+m2mMSVyjT4aRXC6/VQQqR1gHx5FnPtX
t8YEjQhsVDiA73g01M9554I8xurmFb9RnHo3GA73Uc126218JGSy1rVilHEMpil9
r9Yn0pBYG0+UgBtwxfLoh13j8iGP+ANr4agGyh28rGEmmCNSJ8NlRrur8Pdiq8YB
a6uk47lyo7SsJ12Ciquj6frXraP6oEh/iS0kfWzLXb99HkkaPxNuNt0WatmJrGEc
vO73JHZpLU4tnTjMZSb9CFOhdI+et0ZoVZcq49y4C5hljPq+YJ4V95UgZBjuknyU
+i1GiCNyPyem3Db6uFJgjX6bshZMjOjK4cBTwlsbh+2TBtKQU2vd/6Dkh+rhGYDi
xNRorMSZXmY6+CzlY8pNhMGds3W3qUscziW8MH91rhprrWjg6O0X7tCMyuc5Bf8+
0AZM0DZjDv3THRVu3+waVw9vmPNu/KwJy074GjSM6+OylFkbB5pEHgWwl/Dotaj5
91fC/0VYh/jzotWuUDIsW1340YG+A2lpf49lwjISsGKtDUGRrZMjj5uHIpiGxxmx
dSd6xxGDO5ZXby+gczpvobYVhv8fXqpa4CUhez7JcCIZ06ip7Uefk8gEdPd+Ne9h
DWXK4LaoX+Mvvh11uIHsJ4wa3Sla60a+eR9JIuoP2H1JilacEQgdGty3F138RU0u
QQg/wDrgcHaLZ1bjh5cSYvjopOD4h6Tj/t+yK5UQoEXrBgMzIbr+9vjehVvssel/
0ykqgWub2ZgFmnbg9YXg6c0XxEFbz9aXVRma9Vkta2qOQtPHiem4/MGrgTdSINhO
6YhuxOHsaflPD5nS1/Z7VXxlI6yb8XsgiDP3tW5rI2ZhIv0YUoEhP69tD3+hkbST
aKHpqUq6kaLJpdvLu6mcLHyaGxFC0XqGVlk//DkwktaoJoAQjUV+mN9LCZzc/rRl
sHwpABqsIrG9z7P+uvjMpk9C574vsSipqi9gEFq804fJSYK//C9ani5Nbdp7MXh6
nwJiEykd+wgZz4dazRur673UrOTEyaSEZASspLlxAWzDaTWZ1FYrPGAJiGkKxSaC
2yAncDC0qbN+gFepfBFFpWDco97P/k2yUmt/dZO2o3vSFmLaiUcGdi5voKeejNX9
j6f0Qm+4EC6pw7VM0wO25TBfHr3/L4Uys3j2MdUQc/JrrkNv6s2KEbpXn9hQ0XAo
o/BtlPx6kw4v7l1l41ITBkNWC1ocad/kCZiOHgQGbOHTveFDgWZvkIgyzbHaf9M5
KrnFndapKkxkSF/NjW3hlRB8cY9jh2+aBQwcXqd9J6/6hkzzUv6WDaMsaEuJStLs
/7mPg0jWWkCqPk6rhCfs6Nl0ZC/4JIsv4PKno40CbJ7Ug7xPZIJTca/IvmJZH/XG
CterS6Uq80lJelk7pFu4IDd6nBCaGZ37N6MOyEJB5PLgoBxcTfnNwp8RNCll62B7
fZ4kbMxhOq110kdk1xne/uRrckTIIxth1NccVPKfTJfmcj0sH6udGgUmEhy05Hd0
FV0OsjmEjOVHnNNGRgKSnbx+Di5qkQkrKbvNW83TkJ8C4BGM0iLHIED9ZmPfTWBK
jSJlhXZCvt6Ij4PNVQksHyN/+j/PthnaSAA9dBrK0X+5y1ornLzWkoSDV0Yw4avs
vIo2AR4Hw0/4cyILoUZiP9cplDWCOXyFmdYXuPgIoyp73gzAP/uM2RMUiMb2Qs1g
Dq0GFNAPQze/TaD6fQUjwhBgOCnTIBLvHWvfot5jScnFOYFOaLcHsLa672Nvip3i
6NDoMZazDuoL8SKMY3s3vTADZRXzGXDqB/j2TRahqlHMwJkWV1FT4CELvzz8GIj1
dbRDgiqCZQRufD59uvFX7PZzG6V8CjH3C9GArhY0SshIsr1llGGG32Rrk+cuT0Oe
RqsadHa30AzJCv2HwSQakU6iA+4hd/Ty7YL6qirkZc8RzaC0YhtN7GpRKMcDpvDt
lJeMIZMxgzPNsYI8DRoMXKfpb5R46zBvujFNq/mBaW69nyZ5rM0yojSOj/gGyRT8
Fh5zdYbvQGJ4IzErNDjvBCyi1cRG2cOZxUFH01sdrPYW17FykRsN75iWsEBKW8KL
5Uj1Rn0DdutLzncPdG2RSJj44ynmsAUsa3oCsXEerztKvxe/U5BHgFsZvrRPkDps
9tc4xNa1SALy2h/X1iYDCvia0Zs1UsWT7ZqSNfhoCAcOee+/2HFN36La/zlKlivQ
TlZwQUvgR9NDGPlvr4h6mEuyXB0IrvC6et7kBSdSHwQIuIkyOrexxoqYrCjZy4I0
nyWubv09jjuUDuypibeZrJj3jxYasUn5IwGE49D1rW2k5fYBfbKOqbmAze4o/Sj3
WD8ouOvtrPpImgd/l+Mwq5W9/aL2gVl6WQHTphV1/F+Zjv2o+EE0qd+qrM2D+vqw
hFeiKC82DvSViVx855ediLVAPD5vmfdqKDpGfHK0DWz5P3nTIZ4RAJJRq4zWm/tB
AtyjcT5MPduaJdaY3U8IBPeb4L5LcnkqMKryOban0aIZZDmsGF6jr9sLcjqISske
aq3mmxRiz3FLnCr6rn5/RVy41CShr/0pjmteIRMCEMU/JQGEMJFJWQ6x5v6dkqJe
GCzxCoq3g8X58ObkKQ2ebUR4KmiRsAtctPkorYjXVPEq3o+qiIyUpdON/CCvPnrT
BAI0f80qZqL5SS2XxJQYGnUZpcLBCYpQPSBgeEnZTiA6Oi2t2UxyljO//Kg+ARJu
LmnwOC9s6HEtgG1zBBUvePdPLRh9PU8qLaYFFeJNzVmk/7tpj+RtZVjcVHjz35py
Z485fJOt1x1DOn7ZYazJ1jNhFrrzIRyJpn47mZ4pE0Y4KmsDe1DqnBMLHgXT5jTX
vD/I4hVNqGaX//p8He2yZP2dnh/NhXmdJQjlE6UdJILixUEtBJO4D6BZslu5DAJ2
FcKDjU83W4cW7UK2InfzAQJBzKN43lOcoOwXtHLZByneHi19UPUYdgu17W+Yq2f0
y+Wpaz9lLT7qlxudoMTbATZkxAYmhDX3/JsBeYDHsl5bXeHL5I2KX2VEeFXOS0GH
Cy3Zt29zW8ZLRB7mOC1TuieGLPTiRPw5TG9YWmOVWpWskZ3kOUCXQ9Ar9PpBHWZ8
UInblOUznAIf7bo3zuQ2ov+QvxWGRS3j1+8fSof669Milv2Wfkt+LnjOVzcP1y11
VKx4/rdi+5gB7BHH8gD8MKBbmtZA/XekwF35F6u+ItGB8PWDtyogZ9i1aqV3nJv0
VUK8807x5Ps/UZICiUIP0quwhXcRPi5ikigZqwdrM2ESWFwFVIikslOFs8qMLEm0
RCV6TJrVcU/px1OQFNeogttLzQxF/IIlk8IuW5l2ZpJpYwcFacKgbPtC9NI0CLQ0
h3vC6CxkDu4obSyQs3cuhrdY66Wk0/ergwURAL+mEleuZvBADwGRfyGt7pH3qZlo
iayv9RnW7wSOJFAYpncDoVfJz7UcyPnv97FtCLQ5OG8SP8Oe56b4+90galgyD1nP
BH9gwXz1pJiWvjdY75ow7day+5NG8mhYN8DIutMGvowdVh+6hMw2YtKETp84BUt+
sts0LcEPjBZxGz2EwjzXqdmoqz3NOXRLSm3DG65LNcOHNpXOCt0TYe8eWEti5hMT
dAZx5IgiEMA+uq0a7cWlHO1Rp/NhK5kEIHrvg/RpS4ooTp76gX0sanV1TardE9JH
jd/NB5ln1VyL4MLwmPGOPOx9HQWu5odY2VoungeNtjHKlVE0VQSoBfAro+gqNrkT
1nTcc9SsSltN0OpXe05nqFOT1doYZ8O/j4L4kpFk/oVGBVgsaKZFKnRTvawbfuZN
a2+OQYCCI9ck/Z+zy9MfDJawJgXnoPu9XeooPSFNF9PaBiuveu3CJhBRkE9i3ypb
Jap5/KnS7EgdO0IqWGYnSm87KQNIQwC1IG/xIsJNlCfVQxdQ9gRSc/l/Klq3JYlN
5t1jhYEM3F0Os5W99X1sw4SnSc6NApdd2NOtBsLqmMGcVi35Ihnup9ZNoGWF7/p8
yh7JsFmpdHRGRNdGsXa3b98bXxBBb7noZyS8GgD35mycbblYMz9360a60ZchLELj
8/mdxS4sDWi+w5K3q/QpS+7ryCJslZrddHinQDrFOVttV6noRMCykPd19Xz2TlNJ
3lWfk/+X7xyogPBJ/Q1Dt5jLptssFFKvSBHTaqC8gi6cjOZaGCbFnSoTZrvJZox4
t+aPD1WHs4+pBOgGKWR9eg9fzKwRBtKfRZXENZrxqex+/7Atec0nt+q7egow2tV2
3gHJCrPDZgMhmD4i5vSrlhlNW95g4cwOknDXZKL1VzzeUnP3h6hgz11sbqKEC7Mh
g+n3eCBg24m2aeLidDRTmDghR9ZZPWMeTUANKoJXcoWgeo7YYReET4vFWwS4fs1O
H4BpUliogyaHNC9n9JwwZCDpRh58noF/C+EVH9woz9kCr/ZpGx581eStMq1cKwlT
QmKoEHqV6wusGEYnbn8SXIxCIeHuLcuupSlMz0PlDYuI0AhS1z8OwjRv6XyyXmUX
fqvOZQ09/syY001X3ZOiuPz5HZ2co0CmeNLrP1cjY68etJLW9xnBLjhMIUQ3pTK0
AdQtSXEl0Q0oVTtSbjekFcwcvtPJDH/dBMQnGnhjzH0Z2FlHC4vLga/SwnSTTTlK
SrsI2imnX3wEaaSJHVT8ZvSis+pO+wrHSF56QmHYrHMceYfKcAwGuQt+okEDLB4w
k/NtMV07G1CBmJMsKkZJJjpzRLyUEmRsxZYMaJsXtPd+neGBMTTm3m5MByy43yVF
zZxAwXstqnp3IvMa3+mZjt8WPg0RkKRTrDysNPatO3YFgtBRawQl+ROdGZifuipS
gn2aLbn2ssivJ2nC1lFcYqenAqVYRvMHXtl7jtyWsfsQix+PvKK9PYz6EPPFk3fp
vthFTKTAX5p1a6SJjejF/rlgrZ78isEQTCIOgXwPpKkYFYPIHGhX/WWBT6uIaV0B
9R/JAoXDkNgiGzCE6nMYZxIe4r259qcy/UnKm/uRTz6/foS3XLOJwVtU8xscptOF
Fn4WEPN1MaQPwnFoRqteFMRkJoTZ+gzlSkRnQb9bsHPT1GjH4ssJlCEZuqJJ56bL
0/UZlBaZ3ZsSUMVyogxLtWiPLEWbemo1oTs8WBYnTuYDKvZcGmGWu/Muk20lZl8k
MWfIeKtBg0iyhVKrf24EsqNPwaAgYY4CeY0OAba3hM2eA6spIFEhXW72R3JMMarE
V4XllnCKAb7cytujYfKW92/33RK5OBNgupiah9it4yik63omsRVhYRfyjmaSs+Dl
fnst9Yec1Vb+rOan/1aOSGSJcO+YhHkxqd3dDgLfJZK7IO6bBaXjee6HmoY1In4d
zAXmYZTXaOrBRM06tK5EdnYgalciGVOXW5Pp+AxxcadAmch3FSFNoaW/HPEjqzsQ
nTZDbRP2d2fWzpZXA38EoukTeVWbgLA94hYESmv1knlUYT6geLBd/2cNt2YgaBH+
ji4zJ+3cDbGDfA2Ga89PCCyEtHTrXWDVNPrH86yQVKQ7/U7xMkW/LosNRHjw7nEh
Gyxr97Ik1zGObXYnT2apELRxMno2ZUPMJh5liEo2xGl5F4/dIFtK60dBCAsrPDSA
zVxzycokhej9TbhPz7GjJ/NTEnCg+n2KXBwuCkHNQ2VQ6I5Bmfmx+1oCIX+gICa7
QIyyC91SvMt5EL1xz20bf0xeB+HwfbcCtMNtg8aGXMk62Wkis7k/FyQIU9bHozde
Zo1yq7nEv7gKRBZiefGDrMz3DVPXb3eZit9PXA8bWd7cBP6A6rgDopdxseWr4RFe
GCSkktElvKUKnwwBL8DkjSpkbRI4JtXStHZP0fdelKBzkyBggWnqz9WUEVFotvTq
jJfyeqCWaGaUKhw9saGKst0lme6x4RXFam7MGUaCWxiT2SOTT7Y/9Z1FnOSQhNS3
ITsWivgCV4AaTdrTN4b+/8wpdWDTc6pzjA53AhanxRp2mNeLVXnzju4JQaVjC+14
uv3FduMvIRITXfRh2ssu6hBV3XYBjbBFA4EUrjzdttiuMX2cEkTrSsbwqf4aw04P
Z0RiIdchR4aPirDRZsLnjXW3vbth4MRlZqcBNPoehVPvwGuR71JZmhbMWtZ2ymeH
ZwOQReBHOR6wDwgbBYIkegwoDa/r2AmhgQ1PME6YeFyiFDcMlm8QxxRrJw7ZyVcn
/fAESlXH1c2D72A383J0UnydFKOJ18wW8DOKUAqQ46nyrGmhHTlJqxtK2RNr7OsE
tvlCZQRSsiOFHJyw7mkKPNymuY2h25OjkxGSMSK5iMHbobRM1e71E/KTiIdCPJnc
EwQz7Xo7r3QxygNQwnHRmRnfQAreSz9eDQUc8BKUj2nie9Nd5kfg/c9EiRHG6/ZU
iug69jVo4C6tHLJMeFHmlh1i0SmA/d52AzFdOWFNh0to+ux2EMGIEY8iZ0+1zdHq
QOIRMFiHZCmNE6mPxHFI436D1MRgIfoD8LwQWpJxqJ+YEHvrNv5/FExS3wj2lrpd
cYVIkQeIDwcxT/sTRzfuK4180u3WtB2731Y6SniJgCxTng31OyxdIWt+cc0XS4O5
T0T4a1GKwfXc1xPL91ffdyXDKBi+dwFOEnWmU2aHPSQycQAHY+SWGkMwpydw904s
ao3qAsYv7NrkF7aVIo+OJUyK8AVmzP0nEX2QARienV9OJvdkgxkXrrbzTm5i6+Wo
54lR2Ao2WZ3eG7v0ipIzADwwOQTks6orZUNLALYIayFhyG/bI7LSBMEmLWVnqOxI
ezkWBS8GaMLs08sfWNAGqMQvNtp+tviPFOq5LzS8/IX6jXI+pYEGqnz5Nf2Sf4mK
EAuxDtKfPvpQk9LC2CEb44Z8lsmf5ycaf6NDo5pqSoQih6hECWhvpEJDY7zHPatk
GjqdztOOylh4DFMxf3tDXGXc2+cJsPiHQg3zh076kcCrYCuY1eeOmaqbsJXHmWr1
dZFvKSnUzTbIFAgMDen8VtO44RogrJNxQ13WgZt0xzcDZ/eSLJZAFcIng711/aUH
klwV15dXNTPEjI+W+TvuRHOD/Y+n2Ld6ofKYqGAyOZlTCX7YKB3/sqvgrhWcypDb
v/R7fZrCWXyODhdhZ1vpY6Q7RnzoFKV49yMOvPLvI46xNNenzUud8ssDAp5ckmYG
SkC31kwK8LqzdcciJOOEs8n2oNNHM3YHyh76XHgv8fRByxfDrlikXSQ+kSLTH2FF
p6UsYebT4Rs5Hmc3hZuokvssDXi6CTJZGiPKw3POMGbhRXtMfC4KLWQ+ykZqfx/L
9B1GVZsecjkHyYIkuR0zrgdd5ZUA3YhMwOyIfyV5RsVJciPWiQD2HM5/Nts6l5dh
11eNLSwLxgNj6KF8stb0RB7+C3yxGg7Lg2LLtW3f4/Cg0872js/uf/a1UtXSIzaQ
qnlNdIeFNMqhxGlNVLiRX4DcgX4gtcV31K/cNMg5EKQcGRHujJqwBXf3+docK9jR
C/oMrTgc4eWI0OiKmIKlyOMKNnNqBOFRoAMwROlEs1jfC+sANZOCag0eqX7KEJ8X
M0ERmNWsI7pQ2f5HPTGxdV8FcF+oEzC4BX///QY67qs24kEb/ebpiMETt05pGrZU
uCvCKV0NnTNPokHXjJLwkvYhktfLn/T+klPNoIfxC4T6SLIlEypllpBQRPyzvXIW
evHQztBNQlSS/oIYdnUliweAQSmBkmTpR8sShfRF3+PiibkUC9K0wWUce6EA1d5X
CznbLmWd9P+bvFHxNVJBvKh9aP5gNuCoLVxNvtU5KV0fnBLUFqrqLP65xHu1ptR5
12TUbptiMnW3jNMF6i4SiTD20IlLXqwB51blrVBf+IVDHFN4fT+FJFHua7n9NQgc
h+0UcRILRw451fzQkGizXH5JNrOZD1+kRsXSCAmK9YxObnSaoO+xCzg9qPjHQuct
8G+4gwxXtTdX69KAZAfaqIeiL+MYZj1w63VyJYQ7Xi6xeileOzoJ8/86XCnusjEq
Mfp7KQ8CHMWs1yHTHjIrkzZ6Wv8r9wZT5ESEsrslDQRPHM5sAxGIU/gmTF7lSrC9
mwLdLLRqwlhkzzGRBTASjtjhwtOyaTW05YxpirureN8xLQfNj+UXhFGFP+0xdMCD
5EJbd5acK34nL+qbJjAVHVocKTazJNthXHox9PvB4E+bDTptsqy0sXpC1OkxspcD
y/T0IA9YpCiyXpLUU0u/Gkjsm8Z1pppZKf7azw452U7OpRV3ZUdRjvY0MyUVwYaQ
50JTuVsmCc6Z5oyChcwEMFKLqzUoXVbJ3E2UOj9+Y4rjNXQLhcyFI643+GkP77ty
krE0V0SZFfkkpU0oZMgELyRXLNORha6vRezdEzSUVIPG56nDJZ2dK3hG+dZPoxZx
2FEZKIMMLwuNpHAZTjbyghBKYkvKMN7dMxnUdpnk2pj4qOyxPs+x5dGTS38uff2H
C6kWPN4//oyn0JsRqitmr2dfzrCYX/9I9zvkq8KKcZYiTK+kPnooK9mpE7b0vjCT
qH8rebhA7s6purfenUYwbd7GwFKg/dJBqK8/PqRt+LW37sRNNYwn/iGAMjJ94C2b
5BRlfTRbgkqCRvyhdp61MPL/P0Ac3tSTddAzw2r9tbYkt0j4PlF1s4ElT6yL0NxB
NBmVJgE5FvB7uk0/a4GtL414mwIuAnQXe9gl9yqLr6bxptndwKN0i92GF3iDSrHz
z0wnBnuRhJuUTo+k8ptCDzj23dKDISfIIMVVtXh2K3WYnsv3McfYVRaj7GV8BIGe
cm+qOxUsxLcmA/Jr+iY6U2O7IeooSizc/VZmbKlQ0x1uK1o49IRrS4CuEGb075/b
g3evMDQuODUd0xcLSUnPehB4eU1nhpqUZHkzJ/3UV1yYnQeHBDRelEpzRvCLyrfu
PE9hZyNxPDkI7VNeCSWMHq+1eBTzuMczrQ1Ik3YyI1Dtk3qSkj+JR5lZwgEyyCwg
5o6rG0X0xtAJuvV+k5E1jd+4P2988f4o6eC2lJ15KLinoveCbFFvHp7ELzTbdNI9
mFFAcbsBA09/QOrs9Fk+UH2uvwBr9paNYby80eGJ90KofFLXz5l8cZ1kFkF/mmZC
4FIqZCzoDSKw1RsbNFJqhlhYZtt5Ax/RsFeBt0fTGEKNS24f37uoquLfrdAFLZIY
HlzBAIHwK9//Z4f5hKDoz6pD7IdD8Ip1ctA3S3rkkDwyqG413KF17gH8oKsCjwF/
CUU7x4wyEXR0qBVrCSPfJ1HSa5pxwWZsFVbNMMMAcw+f/9mXe8jvd1X4HiifTJ6G
/G5PcuQi56fGuciLgrfFfuySw5GRgJHd21Jxjphk42cKtvFyDbaevHq2ZZPFEM/y
rbZFNmwB2wL8x+ACIoWwdCx18H1GqmnyNQh2xDvYyT0nHzEFDR3SG+mUxskvq9HI
WEecOXXIPJcLt51UO9BM07t3vpCZUHR6k3kh3qm4x5Rw26GuogOMaVCgGEngkbjD
PpafqFd1+CtAHv4ea+iCp7QCJV42/dHrkeyogIIeymgRG7mYS8jwCYFiaSS+sFnS
ZeBq2vo/bNh6Z2dDKu006va6CWb8AvpD5JPPDN6C3Bn/C9GD9TM9vqjiDRy9wPfJ
QxHn25tToYpJjfgmFo54b9OwWZ3hnkV2QT6r8h04o4edOhhvH92tgbVVQenIgU/A
H53qaIh94nkAWl0v4UkwME+w8XFdYUA/q27QY0YxlKVg6GvPeSwEXuJzlV581DxX
nj3Z5FhgBK0OlRg2vtJZz5ATN30tF9yP1p+pcw9TeeCziywgkXCQHKja+kW41dvr
DQBOUCruCoILqjkMCWwHeLIzqo6A3z7HFdhIIsDlt5wDrjiPiTjCGCctVkt9lwgw
xDLpMQWBNSCF/Di1OKfmXReNlsnfskpADROZOCt70fdhBQiA2a3phGNbm6b0i5tf
4+xbAohFuRrD3UFC1TUSxHcScXSMZOZDhgwgkcaPE/oMVJjbsymZ9WbfRwta+yhw
0pkBfqlOUGGuZhFpbmK6gKmbGYkH0bbe9TOFHcIBr///9dFhQzapLUpHSvBjOg+j
qG78IqsHEkUKN5jyiRQPuIPBsmKA39UFi2mhQK2BJxPR7lf8Q0RRjdDFliLIWxOu
Yy2Cs8uHOvslBwj0kTIBtjKwkFGhWB3EHopmNfk/T52YSvcbVP2zpXFjeO7ZqmRE
teWlV7YXtqJrFwxVmnPkFA1728ekg/Dx6UX89MWXIWJNuy1YZP6RYHq9BTf2auXu
7MjVYBimnaTIa5ghxYUTnPSK48Bj2nW0iooqbuxEO2SMUUULQoqoHmuk+kmgNCRm
p/UDXJkS6Y9ShNB3QKbsGdDuVtnd6HQ4OKDYkVVNQF2Q6gFpjXGElu1+PP0SICwB
HaPYPbPDKJrSEO0GQDJdsCVtQsgEwsVRG6toPHo9LV5pbrCvaZRhXgo+uj8yOhE3
iYegZblkiAlffkbkcUN8wPOxaOWtUCERqZgsGteK5uxbgu4r31pgiCGNLzstiBXh
LpZo7CGPnh55v/Oyky0he1MWDNxZ/vKUx/KvWcVt9tLYCJMJOd3j0v5Ga+M+0Di2
O/PqxZ3CUkLNkiOWgHbiMRCGDiapaWrzvBPaIfeu56YvzN6ZzzXXidzRr5gVCRJ0
2pnt5yygdJfbPB9GjOYBefIBkeXf1fHBcTDlyeG9fxAIDokSWz1gIapLLCgLrv2a
DfOQr+56KuyZiBy6unMo+0iel2WtdWIAvINamX0r6zywza3973wPeCEpTNyJ7FCm
CVAwzCyiP1r+OmKZJtNrFbBypdZjCTMU4l61dfRq3enisBfT5c6uIZ0kPw7zrxyo
sUsLXLHozxDdo638adyUAVv692qtvwQEZQhdW52Gh3Bf+odcnAg4a+o9oCogqio2
cKyfZvEOLyIHhI+IDQRALYNFQfs9MtOv9CJmw/ALUiugKmGOlsfOt8+u0hH1zfv6
MQBMvLF0/FCeKSSNmERazvcbFHrxqTzGt7EhnknS4ikMu+V+1d0B6JjuGpeCmCBs
1XWEzyruw9219AnXfoHYlwEuMWLwwuPkxKkzAxHp9VIP70PDSk9rFKtMJHxOfnxi
jRAbmyv0dAzYdmh8ggJnsd83kDQuEjHC03jENFuW0dHKgq6lqbVhVFFDs6gzq58l
1A95RhiNzveiCovcNNhqe3VvJ7fzIXEOzsTkdW+nbJfqHVKYizHUNrGerVGPPxHY
h7Fj7kl/T6cC94ELGG6ugdsz3wI2Dgh/wfj8K3wmHQvCDUQOQwD7EwL+SauYEqWB
7Om1m1YKZKaVe8ANIJOPGY2qd3j7xsBJ/ZRlP0VjNiorwY57PckNExivXYhmwqOI
Vy7qMP85pGs+w0q4DeUsdLSiW30HayQksdrk2BUz8K7ScMiU8JtxE9YMe/xKmNJ+
q2w+8hoXAHNSXFTWmzXuJG10o1AgYr60TQwdlQGCA6lIQjU22N84eqiwN3q/b7r2
TlALvGX34ChfdQd1CrY/Sc+ZD2uO/p9O9p2ncSmeGxn4wfClEa5r78IBRdgEKjoa
15oBUG+s2GGOVBSe1P1pws+vKadrPfuIopMPOrmawoTt2zMXaznnyFwxJzuG1umc
P17W0gruQYXu4+oojSemFgtdnLUQ3L2w/2pGb3Sdu3dNreg2ktyJ6lqI8HzbXxf2
mqrbQTXYBkU0ge9vYQGDBl6NKTalkHt/ttNSp0tNjNJCb/jIb7atc1OKtynnv9TY
jy/XFJkUUXvg7+BuqsrPuXDSmbiL3mdTNFoo4/wje0/k4zQSoX0N9KTOmKDuP5EF
hDAk66MPtagMj6dtryaV4df8rB9cygZlDyu+3DsAkQWDjRAFpDDgUyclGvtDjKxv
X0yt6Q1L5Xy2WOOcbdk4xU0anODT6FQJOzK05gefaOz0LnVDNYoKTtfDZTM8y0U7
0sCBHl4HacjL7N1f5f5yak1mHLtawGNJuARJtpDXd0Jg4Ri3spPbj2yJNJbkuj4t
kZ6t73FHkeHpFPLtREWnTZd2aCMtKgbDvFwt1IHtFQf3DCOWaeXWTNPSOqgvmGWp
TSejVedPccESZTIaXGm0bquRIk2FwMMzPYXF6EgO/6zJcaU+9gFLTwIkz1PYt911
rDLHKZKOVufwh9gSTd6lilNBOTD+9uXLYkO4Yw7LOBaEYMIfgD839pcxQiI42BfD
+AQQGSeS8IgmAP188MCI6I+raMXL5xj6Yqm4tnmIYvuGbk3lHTe64hmoK5fepLc8
qoK7D0QzEfcktgpPwJ+vEFaVRgt2EjOLS1WunMLb+OC/TbZb+b5og7f/ezfM2iDd
pvdQ95GKVlXAgGzLxv024cUZewNp75QXQX3evsfghlHaJzjEOWlF09dY0uN8kHwC
pki7kkzEYeqK25kCtlM3ObYytxV90D8q9qLVcEKCvDxU4FoCl13dApT98mDJGGEZ
pCgApqc/SjY/lwIED/qT+ttbKznrnhGEf6CmX0HIcAKLDxbcuBoMkrisJ1dgMXLE
u2jarUthLTEljIMQiifXfCJds+kPuj6s5VWDQQWG9gZwl6B70G7o9Ng+mSAgAS70
2+MHjdFUAM8E1qt6O/BrunP1flhSbg6Uyhf0UZ6fCWPawFZ70niSMKH5EceYfzp6
d7XcUPIVg6CuzM2XIW4KdYRxn+cDNPJ6gIoY6cwJJtSPXhU5dUrZfsPDhYEpHuFa
QhGwwEN4KJhkkLrRODDLX6TSxmGDCJ8jVjkgaFzT/XBCfLkNXhZE65FwNkjjqlVM
nSNye8GDaTATad1c41FjLK3kEXlWVzMbZ5O0rLIEbnRsrtm8b8vWk7OZ2ehwlW5p
T9nEqZIUMm3/V6xuEzPWAA/eZjGi++aFKZjrYYbP8UU2EquoEPDTvMDY16I2I0Dd
Qr5HF1q9BkzyBvK6I9UxGkendk5ugSfQHMFx27K9hpBXQi4c5oeuN2nijKmJ07jY
LsU9YaJDtyv0RM6OxTg0Vz5p7bzn/LBE0Hsy7VmAlVe3WSr1xDup9W2QpFs0WM/0
Fd6pqEFeHd4bjEJne3muHKmoO8u7z9AgHURf8p0JurqmJ/zVTmslVJSfGczeQdZW
uIEyTJi8IuKfQIVPOIoUgOfNmx1i9zsMMNe+Aqf3cH4gwKqwcYCAGQfNTnG/+tS0
FlapsERIQCmx4alod0kyVcRfJg/B91Y7B7fudgl8ilbOam6e5o/W//n6//johRHD
O7fTxh/KFlCyf1EVArzYXk1wizLGo4b+bNPbaVwP1rq+0qM4Tr7Re7AvEXxtapKe
AQuvfnLv8EhOaX6aL2O/qIktwX5UoYy4+Khco4oNpxfF+UVDo/OL6o+Y9b+IKFIs
L1TXH4dGqeuNSUT/XfWunjenk64SlFZ27ZkRtt3Hi3QzPoqP+kqqlp/yg6YzB4I1
u151aXqYKSTWVffiE1vvHzm7t5Gn19kiG7G04Or1K429luLoPr12jBqchlsRt4EA
/MB1COkh3TDv/thY8Yb8VuoslSKFT2JurYyUF1aDNgFEEf8bLVKmpEyusYbXTbN0
H5jkD7RbC3WjpBRm4Ai7Hqpo73O7tfXoysMtLDCnMQmFYweQvGl79mDqwISm8Cgu
1/u0y3l3hosxe2Ztzv5AJgvWP20GQaQi4fdqaMY50rD4Pxt4fTTpSQ7kAGh6Jqmf
Zj1ha6qtPDxCSLc2Aimm8g9t1tIaDuiYNn++3iHWhXtV6/eh2SnJMt9/dcN6H52G
/iA7b0ZiMHq/GGZOBaesqvJSe9akrsT4mr4xj9clEM2wea7S10TmQ8pB2sSGhxGe
8b7Ke0YKufpcl+5zC7A8I1A0ZuupEgjirZDFpvL9sFUR2vBsJY4HdZl+Rt3z7Scm
lStuxnfU7phyWNVwQeR0XsNLQKxRiFgvvxnhcwHeUKgQP4U1oZYIe1r3gnvlrV7Y
uKZfvUg7RRKzNb+bNfO9VIHOQ+T1GxPYghAHEbZXMkUSN3C2CagJqxOqUc2lLq6M
diNvoKkqe8lvzYOIGylNhza1lb7PTAczyMelGUtJIwzn04/ubj0TDZNOF1ajKbtZ
lZdfsoH5gysftL/Bo7alvTmXhp2a0yFChzCc2XUwG0Pfbb/GRqyOAN7TbHTMH+kE
oUfZsbnkmKC2NNbsLPoCNMbpDcb+60BUpBkKacpt9t8yyg9nU999nxyQ5vkoCWrl
eY9JAjG0ZrKoejfBA23BVJlTUxYuCJU+3Cojj3rtyQo8N5T6WOrbYRF6GfZQtOV2
fURxx8AUK+hG9rAB2zdTc23AH84+MyTfqCPC7pKWRDQSl37u2sFUv9yYwPCj51JH
A/MW8YjsvXUWzF9k0SjM2rC7faUZiGxnVysNJWuHEVLtCapReCEHW3qIVElcfPGW
RmPtFh61msbHfuPFcDKjSoel3O/csh6stOwX1KU9luWJdUqY9c+M5NlrWtX5ZXyI
KPj9SRasg0sNHLgHBqtNo3rjQD2F+FOZarpQ2zQv7Mky+HzOjfq/TDzfdKOS2kyO
kllMbvI9XFfBiJZhcuTSQaQiZeK4Z7Rj57DstidkusdL2hQvS4n05sVi/XVLJbxm
lBVF5tTcvN3bg+NZsg7LFbnAC6XPk1qFqL0CFElrwArH4o4IUfWHWK31Ozml17Rt
+Qvr9U6XRgNhtV3hRbHj/w4zIGFMpIR/0j9IJ9N0cL60yCEbDizUG0T05sh0troH
f4WNnRtvBp1nTjGVhGS43iTBVo3mS+eBdMYJFdQ1awQPPwdpTKR13e7OIHPyhDHl
DSLBVXQMeFtS3JtPmwpvS03QvUyL+7Lv4htCp/hjap4+nuulLCnP/U4lQ80O9lyq
9mNqDOsJRq1PY/NXaNqtNqx8Pz0pcbRa+jXi1I+0/tFqiXJ9gHBjfhmvz96pveBO
TzsrDVlrlK5sim/KXAc2rdAINFtRO18Bemtu4t73TU+MWcF7yBjda9TC4wSRgKNt
bfgMM4jlm1vcU5qJmZBswV1mJG1gft4Uo0g6jYiZNg6D4um+LpiFi9nP1f2bEqrZ
OKE9K/+3EYXSA6NCwtAWjwBuoEi1UvQnsMUlBFaIy6Gl4+FIlSVRydcz2ZROYU+5
70inYDmz6iS9CTPzkgAs0ghs6ZY+W8+IfAs7A/2CI9VzwpuGuLCmtQToDhC6LmR/
dCuF7FiSRygRJCqfXomdJI5nXX4TrW0SsdQnG0YHE3aB/xPm8lXpyYe4T3cwUIJ+
HD2geRFWMbAj2jbBVBp+arZbvcdPszUKYXLn9KdJfXT3QciAwGfn5dB+uhFh+3ex
FoC+uqKj5l6C7eYmxR89boDx7YhG0XBhUoV2liR0e4kQ3SpBQbSxZDvhKzKHHDVS
X+KVZtO+BsJzXXadrXe3zDNovh91mJWDvL9YJ+dhcqN+WUxkzJRBroC5gecdTHfu
+HizC7LE0fjaPjf5WHXxXV7hBf7SHO4Tz7HnIPgvaUUEyhAVcjDiv4FkQDyR0ncx
smJRAJ+ZzfOeyHBPGtEg/aW9I6KF81+3R+VJVlkrnyopbDMecJ2D5wMCe11VmXCB
FRiq0NJiZJG811e2ilkPDVDIQ2oZ7VEZOrw5e9z2uCet1T5aLCj5dLs/VWN1wjsl
s4ucjbL7N1i7tmbRmnMN1YhtVbTJ3/mceLJb7nz7KvGozfiLy1tT1NJtE0dzVr/d
PjzasKob9vrzGHn0JReS6Ime/oxIFCOAAg3cF7D3lwDpFr4/Cr2N5aCp2wHUT9/0
cFV8tHd9g1R3XFYIip2TY2O8vQdlKnKeYivGavrTSDve58BMRkXYi1iT3n5sN6Ew
LSa8O+3m/eKdlU21Ld4U8G27nYjaYi1XaJMKEu2WAWkx+QGBrXSpVn2A3zLB9XCG
X7GcuOTcAwrxzF18fhQDhJMeYWudEUTShJ5vSvh7+HWnvODYbmaVdFcQEJ567waa
UbN9QjMfkvsoHGFqfcPOOpW76e3DYao0hSKtDF/iTyv2/WKqaamFCg6UEJX4FxJe
MzWVjECn9r4oxlIDb7xrIkn/Mi8YlNhO0RN4YqJbfNAI0TV3QysIHvbquvoPHjNr
LJQDplszgQLuppxMxEe7N/GIfjtI11LpiZQKAe1a+gY9oBof+YM0khI7WGvae0gH
DqMc6O2DofEPq+dZJXJvOQbUFOnqTPia5smyjxbWK90116UtI8BzdGLf+hr1FF7E
bQc6Wszi6zrHv8yX8gNbTypvbnXqDqaguweSrBgZ8PsrtrvON1FFahAtmEdqkZ8j
8S8AD0SIYOk/O4u0wWVDSiLwxRgLsSIX8ygrAFvuBDsJ3VkotLtPZ5AbrlrT+wmX
voG1UFOYFyw3d+HbTID7h/tstQekS4SYm4MambEYNwLFeMXsXoOR2W5zeDKThRnu
3MI7OB8kFo8Jf4YXZdu+uteBy8Ih+8raWbO4tCsxmVkRnARuYDTi+sQB9beAmqCO
OJCGsvRAGVIkdGGU7Bxsa/0tQZQfO3o6K1Ahziz9UIg8NF4QEPgFApGvmlpQsTBY
BGr+W6ygh8/Zbq0bEN1EkGEMie3ZNvg/EIrQYQqqhY/jRa4J2TBGvI+cz39ywsbN
DLJZtfdcxuxlyj7Fu4bb7YsogoP0VzggRI61AIipe2J5f10uqX58fZ+SgrP+Blbg
TCYhuNKzlBjhmes0NcqeuQqZJPFyauV/Re1FlJzAlZFj9KmdfJvmJo1ywN6IkfRg
isVO4CLCioHTGsIFW7QpTbPOktpQQJbzs0j15IrIyecYv6Un7VN3lRTJn1fqhCnI
BJGxMedwNFt6BEWmw6YK9Ips0cyRsw9+nGFrFIsPfsGXsd2ispeGy0dv23aXDamM
A7BsvBVKEqmh9vnANWwRlQxWkD8U87RDEyoGqqc4CqBklbAXHbcyJ4Qfg8Eb4TEX
zjf0qvu7T/mjDrWAKk0yzveN1B2R0S7hMYtOrlXhU4zCcykojlwtQfi5G7deEuCF
8/g3fRWvyLLN6AXDJTLJf6i86x3hRpwzl82QNaZs7/hPXDz5BeCMBUfKD75Wvapy
o1KiAn8uewVv/1PFkoxI4Q0RS4jhXF/xCJiG45fJAp4fMN8hUmxDWDO47OMYXwyC
4tFTiVrs+n/zZwk1m0MQ3WcVGlo/X/iHdfGPMYQEAghQILTq1cL7OYwsZCus5qD5
9zq3ndiioA+lAhEnrQZc23TFRO2bxgZ4uFl8pLemyIxFGrIFlPwrAg2QawlxWP2h
H+1MDaXieDWLBpQsKQMAOJGrwmLrqhl2DaHIBRyK38+DrMaVJrXIp8oBwE2kIq30
9ce33xc09UdaXioeMhs3h05WjQmjwsVci9ogyLor/69v89mG1emsvYq6VziPQpB7
3u/4MhnbtdQzvnUk368+u0MCNvAAIy9g8Ea8686ejzxo+Wx9TyR+pCihm5xEGQq+
skodSCLEdXFS6+AAoDn3X1+r7G1aXi5maTYEL0HpT7GPon4TSZ4ACACeAkl8lvY7
J3rNX39tmAZdPCecbFj6N6KdG07PX9lWNGTqyaAqM53XAswDXvkbsbns27x8iL6S
SyaqxZ+9aW338wpJehpIJGA+Kph9A+3i0I0FMwkxSoqlpMzRTDK679BhrGZ0+tap
O0bl+Wa3oOhB0F40/3g3Cko4O8tnYE7Mify+qoEJGj1hOLTbHMLwudkFSvh6uLCn
yIbkXF9lMS0QDlYySYWD9iza1idbW+WLpoI/zOkCufaw9+spDVH+OJ3PRmkp/A/B
L+pBl/X5S4HGwrehpihBiCMS9Cg8KIGUBURye+Yy69H1Q1c40XVbiSXiFg5Vi5P0
5sBA/2IKzsLHX4zLZ+50XkIGRo/IuVbzcDYoS9eEXDP15x8tsM7hGmPk0TWJEPqa
2PRgg009Sy6IVOsjPg/BMOLcyYzE9538pbdZajsRcjw+8goGWJBNAnSJJL3ibt6U
ru4efvDbYqYbjHm73g7seE/G8kWtoNk7DaXagMK0gnt4NQxaEnE7CSSZLRoNKJbw
PpOmd+ZS21XxcOgTHsFwg+2NN/BoZm9KLKPH7051Cq9SpDTtM4QL0wrevoXRRRuC
EiJb4IY7GyJ/qbi3NL4U046058I2F9xZWjXRXHdX7m2PZMWRiXy0riNr6me0n2SL
zrSHWoQZ6nHpjR54d7dHdGtM298tKicsVwgrAgRTmjZWutWyJdZqPuTG+QQH2QSN
+2AvAuJVv13Ss4n6gTQUM6RWuUtogTBmKlkqcFLYuswAA/FKF1NUUTGk9FgjPVYD
DA1G30ErNsPkoLdrohmjhbMwhu2ogeOD/9t+OpwJllhRmj+i8EFcYJ0ccALJ4Cto
nSmlrlPwF/x0Ln+djtjY+8dkFBHVj0tJunPexBuE0jEHkUadlputWudPX5ZqT9BB
XcrcA+52uwMjUKyt9Wc60mzWIaQUQjN+nPgMtqaaZgg4+RyAk9d7httbG7gvxPJC
aaDWYxQlu30YsubvHcdGtON4Vu5p/ZM1YM3Mh6Vr3ita64w/9gw9oH3jQpaG7luc
v5hlJm0mwySWoPOM2+hVybTfxgN/OLTBsIjm/oyP5BEaMiMzeYmdoyHrckdjqU/c
Lsy47zgHpqQWEJTn9eghBAj1WOQlueTCEIM9qLQj34Gt8JzmmpGC22xenpR0Z60a
uvCYznScc79hxkMDXd6NzmHynYIH6s1UfRj1buZIETX6LxE/njd7rij97L0X9y1G
jtTSnjFM3GBstWS6YaDHsGJ56JKuib7iYA6b02nblsmPdCKOzRJdm2almNvMz3VP
pex9j2kJ0Bz7Fiwtpxy/CmopaVbbOnyyJqtY7LA33dqmZ5wC98ONujX+ucXrkhZn
kGoJnDGRl7WMvn5ohgrxd86qk3uZ8volFqpC33EWJlap8OQX8jzgBvezHTFTKuBh
ycBRkPBM6uu6EAIRf28ooxdIjmODipyQ4YqcZV5/CE+PfoY5AFlND6NDyJrDw69q
fv2HhgNLtIlGinTBdv+NT814e9SzpSRNrHeCZHRJVi/qX+uiWH75S9mlhj5XIhsa
L0eZBdSOT8xHzbi2YqnpFvIRBRxMvBrZq7yzITs/wQ1xrJltMnrBc6L4AlqGK0C5
Ws2PsNf6bdLYj0jr9HC0n2cVMnoFg7Q6HwgNMYCDeky7kCRedxgyQrkmZ3riX4Ma
c7lV6OwIG7hF6AabFpsWZINrYN8IBkeeFKeJvs7q88sYWy/03KiexSf5i4Q8bFHh
JlUCK0+llHPWNHlhCRS1Bj71cff1G8FBeOdlA4H7X/VuY7l0g6kFEbYd9LggsB9Z
pCPuIxQzKaswWzfDvKPW7Acpn+fhOCS7r9MW1urFwBC6lUw8nn9U3I4ZoEDa0feK
MrQjLLmRIZz0lB5VdCS+65FxF6cW8IUA3G+Gyac21r9IWiKjvtp+8zx7ySjBoZoR
5PmvBMvPCHVNm4x5KnAd2WJ2yDRj7PMcyKT/i4mprGrA+n5Uk/ZTRSXzQqqCs9NT
0YMdBDQf7clyl7pdiJJxo/l7rmb8ZGMn4fPuzYm/ylFRt45pahwVMyNhxnnlTcbV
zVh5iS8epIYKvt3M/q8UkAB9/eOoQPhiLxukI6eZ705TzQN7XBNPtU//QQtCwFt+
Jcvt2MhK8Y/oSoLYyphQZ2JbiRQvjuDPxW2rYz0uAvKyL7fjnjoyxVTY1sBAGoaN
tcF+c86B7f6F3p8sStoPqJSiMcBT1GWWZ2jhBVqjelUbX+4Te48wJ2dK9KIXa0qR
ZB7vkXeiumS3EHEKWU+EYYjI5rSu0CpaFFHVzfoVWXektVjWzS4wQF1gqtxqOOq+
H4clIFX26SMRf+NWS/xjI4xLznEGljlqdImIoJ2hkgUJbctaN8Qx1tCyAFuCqqpf
SftX4vYIxDwFSEgdBXFmPbYWdMm3w+lf2IwlIm5GpqgeILw/NUJcG0KEAnj7IxJH
aBZH4SNoZHAlTCZzlsam3a0PKQKZBPbG5tLnPLpCgIOQXx1lIhgan+r8//SUm/eL
lB7LU/B/h2RyO3QZoT2EYWUcVVZado4pUAsYStyM8CKxYlTwPuWcGxAvIC3NQ1wI
CcwivG0tL84MN4KG/IRrKaZby6KXrY0fphU67ysjTIa5VeaSm7WGAkn6dFEFCg3S
jV7ARxHKYRTkbo8FhDW86PPlH9AMhZvOMfwyrJXLrn993U60e42af1/6/RB8V8K0
UqLsx/bSnwFd4jxO9bFG894M0Eo5w0dFz1yIIuAYeKY6HiMYm539H9H7whoBw5Iu
3sCjoH/akLk3ypZiL9hYVbU1ZrFfGDAGYNepkGGceuiJwrqYDm4s1FsP0TX8Wkqh
SgYGFmiJ4lhmRf6UgRei1PSpE87XM2uX13mqL5pP0BeDB+2kIBc3TFRhJo8bGOn+
gX3PfDcOb6AFGlQL0yfqlibwIHa7YvuIynSNK1Nt5XCU0qrHL4YgwtVAvUGX+iGM
If3WABkC8HaD3L/KlVRFz+SMdOMvncr2TKhfbFjIqN2x6q6oQsiT0oZI+XWUOTso
AtxB5GxhJaJ8DdvZKBH2Mxwe04r9gncbg0WmcC3IHGlcC8g+cX04KAhFxcvq78EB
/utfgyO04bfcwwMfTeSAszBn/U+4QGFd/vYvfG9c9VYloBShWl3vf6koILbnv4Lp
CsokEYc53GUil9yQso8yQKHNv/HnN3EYvfeLEUi3YymbQb5fs4fbbP+lVRUZ+Lhv
UAop85G9yR8DeAm/4SdDvwfjJH/pw1mRlP39KR0acIJSVZEYpd/HCVfvPzGLxKs9
uIvRLCiGUZDWSM/oCgzd5RxBirjqCqUMMM4Xcd1v0cZsZM06X7LOsJspP2iyJMPb
OjbPQrk5MJAkQZKtFOYPyCkVmPVDoLEMqHkdDPWxQPFwPU3lfv52d24RXnAkoDc5
DslQL1XmVlX5kE/iqHURIzY93LAxAHR6qaL3d3MRNf1LvkQ1J5DoskV1E6AF/N3F
3FDnolb5Az85GA9OXXxb2nk5+hniKC++iQujQ6VRmPl6gPgofAZePu7I8GSIwOyn
t5QkeAsJnJdaJ6aLI+1ky0HqXzMo0GEhRz15lf5yXe7zbJanNM7321JND8qhOPrr
qxMsV3MOdLptjVeg5JZ/crbUPZ1RUWbE4cD+kP5GzFiiC+Eqphfus7VpTivRaEi7
M12QN1HPUu6XJ7PlwTmfxDXPjtoHheJETl9TXQ14Tnq5PR8ApPtZp/hGGschwwxo
w3al7xtK+kH9xPtMZZ1yaBAy4Rf/gu9W5MZVcs9/sNQlav6p9XH0c+2mpK3D595u
sIffe6zk2EoY7utPK2ufRuQMUb0Hq7Wy+5eZodCAQBuJwPPMQhnTC/zXw1Cpavn5
8vftARygVqXM4NnKMBzDqxugfZ5F0JrG4zeuxSB1ePdHO8s9QQ7xoIyBYfvST3O0
1XrvDqVuIpOPC/He3MKuM6qREIM+WBF0odUDIpskis1WzevswRTJFHsIgcrhygkN
9ldMY+raprHi1RD0LIVpgB5S9HNNRL8s0i9RgZwrjpZAFSaWN0mYYotL4zyCTanq
M2CANs9Us1XPJjnDR8Qz78ZtVkutMbg02eG9nTxQyIWezyjLqr9f+PjMpMmoi+FO
aBBYKveL1AtAl4cZeVa+ydwmTHUpSIu0VASYTraJFL1E9lhZme7EuubYaQ4elOWV
w2++EbZyVb/Bm0a2sr10sfutFN6IdpV685iIAbf+qBJkKBnpmlFATKmA8lepovbG
izJEnvCNFVd8PY1TDtV03vR3EpWkqRSRpPHM5rtfENXtOREa+r+PbtM/coa23GW4
00b0i/8SB++IU/Gu5Cew8Vi/KQ/ltWguNyQD/ucbUKQONAOc2nKoKBzM4Z5vAx2J
59//nod16vFnuRfkPsYXawyByqiL7kNLtg2w2pL5R+XTV3kI2eLBOO7FkLwe6O8D
pRf7cVPtN9+YL3awKP1n4YkdsDWq0GcpbHKlHLQwpS27jZvfry9qg5o1UBhP1SQk
iq55jiUsIWi349NZZ7+m5pT95IPK+xdrfQuZzA8bKovzEDNa3hNHZu6LbfhZdbcw
kqxwcKodwk0z9nv4deZANgCfSl5LlpZgY14lQ2Ps6qn/RQjO74CszjlzmsG8YNO8
g71DlZ/whFl7vAG0jAzN9mvBmz6T7SEltn03z72HSZIzUzYM2CsuvZbM4IvOgqY3
LrZ3g53aHBGgrsYXv/XiVnG4YuGUXn1mmKczwurAym+vIF3p1hBm0l4bBTZ+dhBe
Cy1DH7OHR4r8DobujziGKZ3s7udZkxauKfY7B9SccYOiXjqHSH6T7EFGiM6fTlvQ
BBMXCxbt2Vs7aRAOX7zDBFHeauimJu0dUqSKiDLtQTa4ii5spH9MJ+sLxJVb+eLo
x0T6eiCIEk7ds60lECNRg7XO32EpgzzxGarn8J/oQfWCcLFqXqrXoAfTyvB7ZKHh
eLu+lQo1QfCrRdTjuoHeaTZ6NbgAGA567f0FIzLoZw/SFCogBCfHxP+WBYzz2bEC
WSsQ+7HbIwDjUDveKEqthQ8weIshfrUdSiDh3+HN8k3L+A0/quIZqTNVyJ0OqtLu
+4UcrIbFg0scWiFIuhZNka+AQW7esoZHY5lE/25r0wHexLTrH3miEWHnLflzaPfO
Es2fI82IoyHoBbgCjso85oNS4noDcss1/a+jy8bJ+iTymK5IiMe8kAlywyQPtCWr
pO3R3hmzDGgmVjFVNTGL0PCV8LZ9Bhd+B1Q3isAJkO3iEbnZmyRQWYtt63zl1zW3
f8HthIJPq0v7/hhvi+XYrBanh1n5Y0komnYulJhqWRXjt0hB1vXyEqIreZzFYyT1
TEF9rDxhN59dTbzFWXPVpVTh9CoSs+smNncX7MFlyDalN8v+6pindpJKEkv3G8Q7
LEeYliKJWrXaMP1SJZV+fS3sAa45cTcW9iwiN0Jd/+lISMAWv5HSTvQD0a9G+ifC
dFsj+W6CCYln9Htw95HTCyXjy0WHaSCWuvtuurO+Y7RD9a8PKjzr5gkkKJYRUDFm
7SlUvPyhyU0NgoMJ98+oXdGcKqPAY/dYxRtvqetQqWEHV9TYmOvFzEIMYqyUuDmF
KBYx+dK6ZfAuqLNHIt7t1WMX0Hd1Q6EYW0kEGNAVUb2dIF6IVhMgkj1HDhzif66a
k7tCjl3YyEjkdq0xVPr63co6gxpvOo3HFccKFTO1P7/1mMRmku848nHQdJD7+R0G
lmxaSNsvpmGAFkrs7OYFzO4zJauAk+zte+KwgZ7+QeF9KRa7PKsca1/VpIvv1xIK
rc/ql1qQ2Y2IQyAEkgwQh0GQVqVfOCy9ailja/EV3thVOVJXgPddlPJ62VKCwW31
nUhT91qIe3opBUWRBS3K+ZqIF69uGhqmVui0oLpVHL5k8p7zrLVb8vMrGh606Dra
oNNSAQY97xnq3F9MPuButmquD03YatHyt2s+wfvK4jMPHBvw5epcca7kps4rQjzk
PBJCYLzBs029Ia01+X4jn0XT9J/dnPjbAS6gi02J3uWO/nP5f1PPZYUIQzc5sO8W
AtzMt7uY73LDoGaLJrWUrHTUb7WZXVjWmxscT/3Jn3XTx8FKqbPfDvicG3aMJKF4
2axVqT0iaZnDG/3aveJQ4YnBgxG28ADrOEQENuU4VPI9bfbrZK8s6vYTKLFheNV7
QV4lX/U4di4JK1DOqdDemqFg1iTpQ/NMl4KQuSSDi4wK/H522kqFy1j1lLTDmkFf
Shx4hUKl/krql+MHbPwGV9gvQVs0dCqWJhlpb3hbhuUeS5YC2gWZLTrBGmw/ock0
JcRrQutWFzVGaQvzzgUoMOpx10/MbusF0zDsX3KFO+0ChjST8pWWmQQ1m06ImkwB
O5dbQ4KIMIEIJl2CZdTp0cQdfdtQmObp0rV3vkwVqQCQyFbgGHBKF8PLEAE1s3Fq
bMmKHikoZRnWxpX49GoLfYYE31Qjg6NVS+N90hARp4YJTq24FLU6Kq0XJUY/IFAp
o4gEQ7omTeZdy/QeHdx1v7YDE7nAYSmRAQ2CC4+x+46552uJP9Iz1F4WOo6QMB0k
efyUhJQfyRvQxlG0ZCpkn1ygzhxQw0/1O7qSBtFIOVTjUV82ewUn8M0LcDERCJcg
Q2ZwvBCKmimg2beX/3SGbpYcyD8h89tDuqFFQDNWPkWovC/RXheV9TrKjLijzI9c
mt5AliB56POM4P6UBAdmrquxlNTEonxeaEQvQlgrnxeALlkOZZYrq9AsSAX2/J4z
aetlgH1Gm6P+B/Tq3YEikobt4D8lxHkKOHpaWmJBy6ZG+D/IrrO13jZhnOy0HAMZ
DLt2j8DNh5Hxa/rPxDI8cKNW77fQv1TxZdYkUuFEwwgrscyer3cSo35r3WnJu8gn
3huU89khU5UCfqkjjylAGQgaUytSXRfqKmhq+dWKIWxDb8D16djoU8akC6mgYB/j
d/MMXh1SojWBQ/E61V8sbXgDMSdmAn545MMyN+Q7AjYDrX7jUx7vw28nq8THl2VV
qVBs7SO2B8B0khB2+1n8eVvIpifAAD7APN3/cHbxP3K2ZHUQay+V1pktyNxskJQ3
rSnQRcr/woVawTvUCwrHX681G1wgrVQWQMwSu2fiBem3x0zwJpAXRtY8zq5omVYj
K3KxKfyrBRfXTtO5NH9JXbo7j3kzzdSwzI2HNjLDBZXz4D9HKD7bpg8SIF+Z8JWg
MU6Mwni3WkOhOblS0sPSde6nF4T+HPEhHIUJ3kMWv3cKfu/J6E+++xblJBlNuq4D
pxz7ISyGW1t6tj7CTAGgPNrKqYMlbyX95I0ZqNYdk7Cj8ZOsOA9ueCjqVZCD2RLM
rm21ZAglZfUd6UAqJO6PbXkHrqQx4XXxA7YOWtHD/3qb5gAmuYC1UNPtlb+NhaAp
pC0KwJsvY+a7/2CCGrdMxnEaFErV0GfcT2sxx1jVj2VIB1WNmsbs+k177GTSyG42
CeEljZZAN0kli63a6cJVt9XQ+itP+iHbFdWSXhHg0Fq5QisKIo5BVCFTWfX1zEh7
uDkJDwRvhDEeKnLkGk+w0NebbhHaXHWah2NQXoaF3XQKv51VjkaUtxVSHCmkl1Fp
j6OkDPpCMu/P5hNXWD17pI2jIpUsUbn5nIrW+SLC6peLyycF+e/IZtG15LS/WC4O
uS47VQuNAyVTL1wYfIrFsouszgAD8kFfAKfUWucylqQ82jdyLozZRHW/7CaW+S9j
/+egUzeDT3HAjWN9ewN83KU2vnukmnnRZR4uAY2uSpmJFSoFiBs8p3j6mpddlLJN
kCodPyq/NPPdrnKrgrdHivs1P8LbllX5d3aMV+3dAd7JVGsZoIPTCT7Cdqqal7bd
UqqPgUP0d0RMmSqQAtTDVmADFKRQIO2DHWxQzPfK0yvPZ44uuMjpDtesA04czXw9
vI/qHdY8ZSrwpgaonK3FBXvgwA/9E8bcLaR2gZXHhnVJe6iWZw16nCrJbBdktO/s
YarJ/jvelXmw8FzMIAbAN4+3KE4cqcmr6yLIcltHzmxBtT6GgZ2CyNy49YnKgQWe
pgzbcGO0Me5JrVnl9JY09EnDUAM72m7MYkDNmliaLTp4ffQrZrKWOIOvrDca2cIM
5GnwxKY0uD11dZlwfYGFfFiQ4hKrW4ow/mn7GDTFW+IBYClBr2FQiHb2hbiMAUtZ
JYsxhKz5+i9wArEoj9iN2Alm6/mrZ8yfoVvzJhkPg3vGS8MdnQi6ezrJ+FObQPTX
+iO72sKD5ZfURabs61UkEuPBzRe9Z1rVnFpxcmyJlbEAzYrQDXNUjc6+S1b8K3LY
McAxCRn467UobzBHrfKD+bLvgv9QtbYW3b+EH7DAZ56aCwpUu3Coh/uKDnZEgIBT
pOFn6ANBKKKv3afwqqcYbt/knisFBmxGZE6QQ4HIss1OK4rjUU7xb3A1SuwBTX47
BkW+VIK0BV5oQdm+YLUf+kXre5HR7YZCMBHu6DNHGeCeIr/m028v8H+bCR+qQ1cf
mswdLI7GziFcvOOMQE7XX/4lZpOYNmSSrrCUQBAtZskTAmO1BRlATMX862CRH3dp
V5CgD0Ir3vKScJgd7B7nFledlhIOSJULspR6QJ4FSxTyqza7vulQY75NjfAmDzjM
RHyaVNvAjUQLj4Qbw510YGQQUC/7Ddz+BhCq+tn/6xKKEhXZox9L7SwBcz0DXsz/
ml233umMbKxLwVkh18wEKoauCWoEhnZOqMi4iWKSz/8IFEk+RKp7N/k1rqxnQwAh
V7KqInCfmslQ8AGA5h1jSlR8f59IlxEEtOFWostiFcz3iItmLBhnHOP+a5l5soLH
4nqoRMpzL3pG+NBdWry7rBP/aH/beTAnT4jmuS01wwQdcB0tk8BXAhXRif3DVeXJ
rSwnRKBgvPXLkt/AyjO9Vvald5zr7cQoqAhMrNhPZnzBewGIw7DrlFp3l8+U8H2V
SSmBXUaBnF8RXZjFBGLW90aCa/jX+bAK7JsHkxCRq0H8zx1SO3NDg9RdJtWp9O9D
CNs7AWCkK7nKlFG2YBkblejTqLQeHvdpf81CVxAbiaTdDHMkYqzXgn4CCQogAvDp
+jrKltX5Go4wodZ3bmucwtEdOPkGI5ifiEaCK8jipDOs6vOHax1I9O/tAkCHHwEL
kARZPTVGxL7w3Se3fdZP5IUQ3WGNYcXo5o36dM5CvK3hbUkbDWnq2spe03rrOX5o
hZ9/KsEGSs8DWHT16QYI0vBzSGPterWS3PjXW3NB22ld82iHK913SQJei4q2wvrW
LNm2YMcX+3g9J0yqllPcpJBsCeGOr+oqOBnlj1aXoeoKa+WyQbT0WtYr3wrkKAwa
7m2/Ox2908b/wt7uuimBoAqB25BcYcvA1nVRp1Y493S907XNtPtRWHwl0b1r770J
5ryJwsa0SF4xD0S5xiN+4fNvsUPubnIpAJAfcZV7BHXjy+UPGZ+R+kmhDBe8o4J2
btVTxzloJKZgBWrDXsHYAYJBxNrtE5bHediHlFhm6XnmofEgj46lT9H6BK/YpngL
UtcuAFkpn2mVr73iALLvjqvPUUsmMRD6ptjz2bAiicG1pDAshjCESo5nAiH2Tepk
poyCyzbFSnvlRLiINDpBg6opNG8Mr2NUFsJK2kVKuPizcsErt70Fbn90iMQQQjg1
nP9n0k2Tcs3eicpXuxsnXoRnvTk9klYv+R0X+waviuNl5JnokRVqi4WO28fUfDFR
PYwcPHxluWlKv/O3ZSTRdu3er+uQolB4MggWjnSbhSA9V3frRcEioq7Yw+a3SZSD
SErzWFBiG3HoEQUercA/TqyXGL+Ng9VmaKL4UzoOW0p+Gij5d81agkAZThGkNlN+
wKDzWKZM+IhxHUaxCJN4QgDGtxguGPKJcgl17ePJ3jlI7ziqwkww8jKV3jGu3ELd
Z4joY4PcjSmZfvGcAI0mrsfSkvgNXey1jY5uGu5i7vPTMoT9mxJBelTPG3YWXLoB
ZAqEHqko1GgSJHKffiYtYQAy3pF0+N0U6Gtood5uDbEcmNd2wDJlh80xZkfwW0PT
VkdDPJZSCLcrHyxwZ/Zi8qTClABIwLjB6OJAbBX6Y1BAIlzClnfE6oTKApCirSvG
B3RIIxw0g1FPPgDKfvPLq8fbNGPuthNxgIYROzt+uZ05djQBNsMbsSNtD06a9yaV
5Itj7ntw5/yUKazblCwnwInHJ+Rsk0pwsRexajdafRZDOAYpOVqR+Z6WXPz8Wm6b
eLxsQEQQyYgV9I0WvHNi2u36eaJy3wB4/nX+Vyk9l8SoewJxyD0a3g5KjiGINEDW
VnpI2MEQmu0wTzKS/lA6rkTMsxYSy+S6z8ozicFoCrUnyvSqEugGLDRSsM49St7k
TptQJEeYDdex81jd9SoC4tdPzWZCLX8XAkCA8UOWPmb3b/A+tDk2THXyC4luhHz8
vsoPfck5P/teDM9gTXiPddexMOYS27egdyjHAKS3a0Gf8CapGIYT6R9lm8PMZ3Tz
A+uJJ70m8hlQxeRcnuwe9e+7eTa7M4PLxC+2Ey5YjtoPe/odAHFRDaMepLqI5XZf
gSph6ZkQjOsJCeNGq3ZmwhoogU1r6RuQHXctyUbFm0OMkwAKm/SmNvNbSlVbmTnI
YBG+YgZq00qnz8bUHhrErJ3AMOq/RBkxknLViO9Cr6daJMw4wJc3NXJVF3Vkf93C
X7b61ZoJkEHa7yEmm4rsOZ4X3HONiH/0gcXxgXlcRDLl3OMuMG4KgW7HLRD3nlC7
52pk/yT9nUNehc+O3ft/NDEpAhfqT8Ungf8YosRqh/wB1pP77j8hr8+kOmVhRqgj
ssYMuJF9tBh6PB7SpqBDsvmza5DeR3+2QI/j7RVjURjerTJwsUwnHHAxwwOLcf9c
+8C2c7nZtb/xv3Rj0aN/p7mv3lMmd5lCNJIZNkzvKfZGEt8OVeV0ksrJQdloVRag
fgy8wKc3xnj5BI/tWreYYEU/MGCA1NcwU4+4W7rHMdWpyxYSqDquBTcVjYLpfgsw
ETsG44CvrYIFxKIh9khHzVXijtcX8Lbdp0YGCaBIIXvnz0mbxYCS17Da5kj/baME
aXaxnScp6TyqP6SyFS9ZhvDldsFZfKz1mLWwBzSyrnT6gt69s3Nrcgo3coayFaqb
xqsmeUMyPamOa5m7Ddn6WZLDO0sXtGYFcKIr1pFJM9NUrKiWCGNu3Odtezlclr1x
TStjMNCGxsBDT/AJ2WGk7YQFI+ur475NgtTwuTgFm+5UwzBveDY5zaMrm1YFxy3/
RTy7PHq39sJF0zpAAmcXMmSJYN7VGrAux/r1JlysHQx4Aagwu62JmSeCl3OWm/yu
3UPZfj/6cMyZIvqxC1zCPX4aHvmRH5bYhIg4BgIjebYOHMT3wlTtIbjyrzALicYk
9ZjkRmNu5yNIN8JgEQwbg4mh1IKXMiJuzfTIJeyOvR7liU8pYmMMxiJfcptO3mKb
o08zt00l1X8cKHzoF9yoTZQHOcDDr+vkTJK3vL3TfvM/wxbtwRh0XwulhMVtzEik
gaf4bxJaBh92rdTr0qKuM07yQYgWlXNRtuxs6ApprZSGLf/1k9id5RxnlnrkfdjY
y1jxcH3q8MKeiILwWdQhcusurEuOK7KrD4zpTqbtCbfCPsGep9jqtaPs3qCmXeMX
0MLggf7eFcAB/ycnKnRhLGoE40fsptJypUoNJmAiVThQvBLbaxSWhZl1/onlBY3T
/aCI0E/dU5vqeLdZ9efXOfwA5Yk1bfpqmuYjuh2O8HrBJ2cgePqeF231NpYMjI2u
MTR8se8mnZEPR0v1xSuDpPRVKj+sPDQfgp299rVTCf0+mnnigWVya9WOTvT3jyxd
u5pPfZwLefAdtgOISIqZJDnWOJi5iSlr7DIHh5py/1TvHhQmVGs+gxVASpWLSdHV
yMtpab7DccSe2w/igM6VRXyNYODFGS5H4MWTARzsEAp/l8SvdINvylE302/NC9ky
gLWOzh+w2fM5jlHXrdjnV/+HThazKqQzNHswR/8NLwJfXvlsYzdMXe/hrhlgLr+B
n0dhbBxs+9mGKYAXsxjAhUzCJCf47NiC6KTSkhn+ZFM7ZYxrvTniWGpxCqiORsW8
rlBFNnTO5AAbbdh1Par6ODkJNkkvZMZXdmZio8pa4LRoObUt2zdETXddD4ver/ht
EbsY3zmE59PoNQf0ouCgAdmygnqz15ssS2V/ovtEw/cxTTI47HdcPtzWas2t0a0F
W9dMLdQanqXZtUw0w08ERbkbIVWHmtfi4L0sEjRvxix+1ivAnb185Ug4vR8gdckx
4qSPQDhSwPZXuwoEa1Z3xD29YTsiO2PgqUruLcg3hi4/ZOuZe0AiTbUkkJnuwbJC
yMe2sTd5NGMS9TQcm66/QUKXdpczJIMbLTi5VTjVlFse3EN+64iP7e794iOUsspO
MD0qKXoSARlRv9ImxLhNdOCZZmKo3CL/gn6Ty7zvWs58eYLCO3rInGoYoXg8CfSY
5pBp6sNNxEri7J8CJ6JgDLwdR/9uCP9DsR6ojfpwY9oiy0paILkLU8ahML4LJSK6
FUFdMqe+/z5hJhNwHccuRmWv7iHVQu0aRXOCY+47U9PbDTpGmut3JaL1bn5dT6WI
srUjZZnjDPHa+Qsh3ud3HW6ynNo1PcyWw8t8r67JbUE6xbM4JPy+o/EzKK1EnkqS
GcBWV8msg0KMjstWOBMWt8RGYjjqSIBuGw2I6/bqIdB/2uVWGK/LnDKPi1V2677q
lLxZ99ei3G0uyQi7IZtTdCQumeUkQgMXWGutSf0NixUxWHa532S6Tc7l9GTdePtc
j/2KDSv4s3bYnIvv7m/qnSFMdBFtPtybykCNY6SJbighHTD8rRM4AZZA8+Modpuh
yRAsu3p+gADUhEEJPzx0/9ZF7AEFL1zsUvjp0G1WLGLJpVbpfQvTVWAOcD2waHCL
+u2qPNJqDWnpmGYyVSBevqkBjSwCXNxwt33x+PnYTqIpUxl1gAVYycqLxETzkm7B
SD7n1LA/K9HfsVqraVwAqXwQwZhKORIabYZgX+Fu+r+lADQ/jz94eiAvugkaiOSc
UJ/lCP3cyros8TvNVvTWUCFetlfxq6vJhM1VaJZyDMPfJO6GLzlxx6HkQlzdNESH
l8LI8VW323xVIiyHVv6xmcXxN1J4Mmq2SFo6JHkxw76HALwDGGTnnjZbsnIeUtmY
hdatfLOgtXfTr9mvKVo71Qsj7URfxKUAr67GiHP1Qw6GDF4B+G9rOs4aL1JUQB71
0o4ey8RsIeZbXDidxPCy6u+tve39LvKW0MmG+MEAk5UrOwE3lD0YOXdQH+D782TD
lP502mVwTrHmwlnqVHTt9u/KFNuRe44U35/i5sWAnqBYd8q8Qwt6oJU22mhWpczl
FMlBk6aYNKKWwGzWxZm4ejeWv+44Q071oC4s9QCrhUwWpfGnGl2rnAEqW0rFGbCJ
WLE5wQNYLaXDxOU+YYdQF8SsjTxr4qxhYv0VVjYNCvt33qxlDjxRj1/6IS1znCll
243P3NyMEBjiC/JLf1BTQbLF0BDlj2jSghbq/Zifei+wwi7LvO73GyznUhUgEu5Y
OhyrJUE7WQh5I3Z/0AcnPQ1jBAuMPWNOeInTgU2DfngelnMfPFAPd8ZjiTKXnDR1
ss65iewkywuOocZb8Ey0q9RavtFvYxsM9FubK3ej97lB4m96RIQ1v/Unqw1d3PjY
PFdPi8KynGsf8/21jpk9tO9YwRtJUn65Iwvn1wkGuy6SPhtpJ/f0z4YSEj7REDzP
JbYv2lbOeH32wukkPeqD90SYrfvwbHOUKYQ6dkOzSWNf3WtpSzEyo1gAMosq79tB
gCtHtB8UaI7UL5i5mPgAY7lP05c6riNO5My3V8mVMjU+GU6Um1wQg2L0h1alWpkW
NVXLqvFp6JaeWxPNd6wjTdpDwrWjXhveOAbgKPDOFqAcgFdO3BujWvYYopOLJDge
9P48+ifvNvDPxC4aBSfuZ1qcYXzZLVfLLAqAE+EOY5+x9Z6yjcOXTn2gvp9gNoUD
35t4eS5w7VdinacqUOvBsbj7jupeoCtfzjJp7X8UeVIC97muAHx27+Rtqp8QoeXB
kDf/UDe+oQOLbJL3sAZ1X2Z3E3JdKyCVgd19+DbA+ZjbnpQRb+KK8nDErIB4hEr5
Ne6SPsRYTsY0+pj53rZMEtvPQ3PGiCkRriRPD7DmgOxkFl1Mm/DfmFNKCsHFs6wo
VPdkPt8SEnpyy4wUk531RQJqIZUAY8vLA3FDCeNaUnW0thA6PRHjTjaakRmdTzlj
V+EYdeuI96BKJgr1SWkTuSfp6VRKeoGFhoPujEM/n9SxX0y2/Kt/X2FXATsQu5vh
cyEJpcP5uFuZKupZ+bgsZ4IJMvqwkkbYsOBxoGCX2h/vLBTM8ZcaOFb9Wjs6Ae3k
Jpo+kpLtGuDJSdSTrYJzF8KWgbB2ysSZP0e6G8rX4ELp1Ia29u2isn8qgbZm9NMv
lHzuS+P3ZJLku3JnpLFZbILI8x50qQGl74pv/SOxirP001CaY2Sk1AWzn8T6dOO7
t/Wqfl0r3sVQMaGUdHQdHVVJydomUk7ZWFDpu3UIjv4304lyFZsXBERUz9k8xgbV
4zgm6bTuCs9jNfRWcIKbAaDyYHDfHxnl11kAR+WV09eB1/k1K5hVNCInoMx7YKyc
W/Ogot0PBiR5AaiSLpPCJpUrrwElMp9qmcCdFfzQx95tBk0pTb6dkRVUqy9gJ5tY
MCgGPsdCrc+zDDUiCxDnPZ35uWGabp9dnbE82y0dMoNcoRCoXdHO8PrBvhTkD/4t
vxHdnyWt5pYq0k3s0ad50IZhIUodQ76F8sMFpiSvbZkaVbpoPRPAnKDPp4wHlO6z
f5WxvIGwFWi3wTpNtnAECrDu8ah0M3HcTWifb1i9J0PwERWLWykC2IqVDyjEEfKL
SAgvzDerhflPuv4drqRcKt2zUCgvDsIOnn4lx1D8syrJ17PJE2OBDH83Km9lqw6/
pU/k5gDkzoDtkLGSqOZgLUYF2XxRDRg/uh1DI0VOcupKufrxwvz1SBySWy4AVutC
WUpcRynBfYCsYI3oJF6kUQkoGcn20/oTc7U2qz5p5U8PHXxMUjFTM3RPyI1/2YdK
FyCKz6EurZDbXHQagQN0u//WCCPEJJrjEiaqv3Qe2Sq7uplde/TKIHeiM/K8nhYa
t2Y5FGD3qHWW1BgqqzOBIxk3BenqRUm6xxn0bUiWYsjIWi1KH4VHEPlHz16AwGkk
WZ1CR1SirSm8wRtVcl6MEdrh9OeoTzhczM3kPgJu+v7xs/5Y/QDHyH1grOtbN1uE
8LZL0t2Ce3xwYmaDqRStbf2dEbN+RTh/cfWvybneNqA2AtEii3R9kqQtX2+suaLu
atCfrVboK3Qp3QsNILMNPpXTaKL5wOjYGN+cg+VlZ5KAoSnCLdPl/c/Jznzq3FvH
EG736+wsArITVqmBBSB4J6MrRV/pMxCU41WLBSSGPrKrXzYZn5Ixxi+vAvcrO1cn
pjveRJdAyRd74Tzv/JNyXV6gKWrxiXmtTMCYeyVyx3CxdLqejK085B33gO1okuqJ
CP3JpbTBiCwPvkedkYrXhY4mNBDjHPlxvYcTMMkH/wZxZfO8KwZOa/6ZD66yAFvK
cbKvyQyedY1mxbbMnIlXbzek+4ouMunpf18hg9YpxXTlmoBrRRapIJqDXBychrIO
Dn5ni3VJpf4GnW3IRfU0iaD57qG2lR34AuW7wtSnxXVYrXY/MPczoMyQIwZ/3FK3
vODwi+a9aBEQSWUooA8/xA4xOkTzCaarP6WVqpB8lClsP71MaZIEcPBHfu7IhoE5
JeX5h2OHJt7fmn6/1qxFNOHkhGxD9oJmilYm09xXzeyCF5iqwxxaCUI9dwu1Xj5H
LvyheI1i4wdnwqjzD8xGQmTgC2GDC5HPxpySS5LbbZxHVnSEtyP0REC9+19mENzS
1lMzFMk1KlsHrIak7KimxjyvyPJMYsF+dzX28yHIdbFHlKhcbd6kzhZpucn5hX1b
3T6rAPxrvDQHxcFoLGzEfE+opQGZtj9u7WNGlWF4rH0TMi/IQBUUGd4sWLnHSXMw
y0Gko8C6jAVLyD5K20TCoIl6pwKeY2c0Kud1d8tIukoHe5yUr8v2z6W2MJnI0+JV
Uj9JqZgkg/ShZBHhbpkqm3lXEjJlL/A44WHVaqQBoDYm9vL5J/TuQC08+0lp2ivX
AnQRN9LtrPez3RPD7rvX5voyeSTaHW7c/OuCcf3FTsxEzxcnP4VDuiFqkCagwvm4
CHYDP8jVqLXFy6nuzKlVGY9X+Kc6rLOEuz5D7jKwTi3vmPGMxNk4DtZqo0NISy0S
jsW4tYTwYqvdZIDpYXxrjrfL0PFOFPGoTnlkrI9lwlxNH+++IaC8iBgOfSs3s+6e
UQPa6f+q1z29XauiAkMxG4uu10Feg9vB0ACU5w3ErbJMfYjDMQ7pwhZ7VReyW/6K
IHi3rSoO7xBs6umq2jSEayr934trlLmhvR80R2sSh1HxGXl+u9eTAGIxl1ecyRI6
LL4AXdj/TagwCuM5suxo5wl34UW2tgKch7O4f3xSsVYUEZBtlCZ4KCtL1+0tz1nk
uAyVO5pTx1JD2qwqoK8ah7uiY5aGCVBoFsMuObFAF8adqxDk0OnJ5/6NC+zFhzrF
BWk0F/hJBDilo70dlDwQQVZ+A6eJHz+72+BKnqRBy+VZOH3RJscWyEl6weOOW8UA
Y15C051O24OywYIYBxU2lfIsvg4cMBmffqDwZXSUko0m2x0+H9FXyTZYDFRYef5Q
tbvnOuMCe/c5YkJOiWeUKNIZBAVS/qBXpoCo7ycCSqw8uwvxQ7oaSj6OaVvE9W5d
wtuhDXF3bJKnxjh2w6r+SLWJDr8hFAjs7wVKS3Q6aBMBGexz46nFIv+LefvFYfg4
7O/rhGk46KkOQze0RtnLi6BEa3FRQ6fGZrZ1kHbXhOp9hSskv5BQz+nC3/Kes4e/
ugJGXS5r7+uVA5UCe5ZYiiyZztVcXmqN5ylzQTEyveball6aUotsxad0INh5C+rs
O5u1DecXseaXEvk4Azuxf+xRd8vT1wcoYDCCfo1SAIn+4HzHZaXFKrAdszeHLrS8
tQFwPKDySPmiRcsal4GdAlFJtn7ObhTbRuU88PHwYRXCHyKX0D4cOxnD+dPp/sp7
VLbCO1iy1/HiGH7j4Ga1Zv9acILXS7vw2Rs4OLof9dGZzbf+zXfhIyZ5Va/8XPYs
w6yAiVU8oy+TcRXdVEVAKUJIem+OJfxyE1nW1Y+GJp6cFov6dlMoyRUlb/K+KIhz
aEpz9UhWZDlM6nkUXhOC0AbkMrCn05xvvaMNrJ2VRGpOvIDo6FyVKYUFd2VOQMrY
Xo2EreyX298g2VUodV6kfOwzoZqwuxQz/kKFoWSVcFs8PCAE58I38hiN3gUHNPjK
9+SpmA7ComfWJozPSvl87eqBjElKnWvTdTnx8yYytdm7hIypCWCNQu3JK15D+cN6
l6FDT9pD6LD7bzgv1KsxpiShGzFkg4TOEO0+lSFw+JceJ2RCzfOs3QJt5UnFKoMa
1pQ/bauwmpHkR1vdK8HdPamTu0M7fypgE9gblLU8iV98kuXa2MwJoVzSyv1Rvkc8
NH842AJmi+Rcn4K9b/vgdNWqtLe3JGM6Fy+is+jnehbcdb66JYbdX7jGmhqnwKqH
2FYSjKCX3/CZmRK+Zh96nmeUr/qhn8UTtKK/K7ch9W91FL6m+ZMrvNB4B7arj9Q9
EELvKnFW8+gaILQq5CNvHBQhTLaJITlmkMMrLk1Pa258diRtqPomTT5ht9T7yYN4
d4tdqCgI0GQetaQRQSjsn27U+4xO07423vNhg2J5Uk9THvqTL5bbogUEhdus6H5D
22hm3fLLCkUvYH4cvaadT/AAjqleD2P4DQvoIUhIxlVDI/oARMDVh+MEF+CJJ8Tb
ds/Tq4XSx01d5yIKNcS9u4IgizxED6NoSvO09eI6pL1Vw+qrbNYUbbov3uALevPU
5WdEnrLK575epkzvtCMLiRFyDKiAFTwa4FNJ62N9atN3Sci729lVNaVAua6lnWW/
BMvm4t1DvVOEXuXIx5NmYu4OWWA1qnoL9ugFDoLL1haKauJHwvf9zIrMRLX6CxG9
Nw7MTjWzM81f5LXpF6XUiIe/BhRJ6HHgyNiBlVY2fa+bGCCKCdQEWcbGXxk5qGHg
YyBtyhkjfkN5QsrVWmQaDinukS4DGaP/dblpOOxZD1ykfIeXpGFUqydqVKDU1p4M
NEpNJN4XjfhyCr73sqRutwlUIdKZ6pxgl/chGxxff9L5xZMMo12wuLnC8qiGf7xN
PPxWVBH134a5SKwryzb1Eou/xRTNfEJvGIiOFT9ZVjTNMF9lXScUAwuGRRnogjC3
qBiQdHB8bvC6c9l3jGW19xM+HUxsfv33jwS0cC4ceSMW8Led9vh7WW2AsUpJqP6u
0XYxJTsf1w4h3Z4paaXXJ4dd6Nn7/9Zd++iwFlCwQXfVtc5YkpMwYGy6E3lKj4Zz
3KGpJ2YHNR8nh4+lLlCtGjgjvBqY8Q5uog09JJTaa5NBKwysUwEmOu0rrlOuYyIO
ijOin9AKrWxcQIJ2N2Fh10stuAqT6W4a/33Sn1qqTtIzZNC6k2db6Z/Ka4FosFVW
eqoOy1nUjGDL9mAt5mOiE7ErMN/DARKG9m4mRT2yMJb/P+ngSCWwn8fBsjn/xUV7
zMDiyfvt8RNN4opGeVZ/W8BEsGSKBiuvrA25h8HIrfeYkRHtra9ZB9TZEk/+CC+q
m4LT6NEHOCIf7QKYU4GuANmPi2op3HMw7SaNRTF8ZfTq+JzEI8KDgJ/FHwMNEF69
rEER4b3Wq6rpJaCLbI7FRASK0gwLpnaZt6AI5i7QcpMrrJDk8n5D+ZPKZFUTt/Ym
pue/auBf4qrwE2wW4b2V08PYlLqNkspW7GlAZzALEIJg5s44qnB28iPQsy6eVjY1
MrTyAoeuHuvQTrF+i1ErvYofbEgqSMtv1vDil/vDYaIKQ+IUKp5MDTDrkSPPXYuF
demOT0aI5wdrKhYhrIfYchlAHMAnuw2TukEHgQ3JeC3+TpG9KSlQ4ampH87p3N4o
QSs0ad0VgWvdNgW7XHL6RSICml7EM0YI+Ye/GYH4j61Ms2vkYxoo+A75/Y9fV9ZP
RINUXR4WAIdjFFpIIQitDPsnucZTKQQ8QiyLt6g+8HjpjU5RXPy98Ov3pYnnVFHO
yLGt5B+WgQtNsuIALHHykhslDovyqX7E1GVY1YMbhhIgOioZk9LgEA1waR/w0iZ3
Qt2iaZffSgC/G8nCIlPUcYjqKWLDf2jozUZmOHCz2VdLjTagwoHd2wSC4EJDCt0f
i/kBRN3N6iHLR2KAYWkdx1+whObXK53HAUXhYkTgZ8alpXZ2WrIcETByrnPSGdK/
YYFta3kMLaLroLrngakloz+I3ufdIGURlkYcms2NrfYy6jv6CUR81ksRwvNbfqoX
eULRuzX7YVBXdkI/B8Jj8J0TdB8L8Bj561J1VyaRWbpgouFKXvGXR+CAPDQqsrHW
H0P/AvUPHnep3qzjZiIpVTGMWE/3Fl72Nd2HY/I4c66ZFB19TNGU4nVPNk43UP8n
gwJFQNW94JbQ8gaOiOvvV4IFgYCzliiu/vk9TdkY0oAMagNIN+poLwxTkZbWsni+
f29YIBaNRAb24eXjsZ4lH/S/Q2qpzl1JHvdODv91pG0rikdUJdrMUo8nv+0tFq4s
jpep/NOzsoOeO3ogoNwvDUN/3R0CYnbbu20ivyYp5DxffKF3hS0aPoQSHVMkqF5K
T0twBa45YlJAY0YCIjfPolOCf+cC6Noy4A/OKnuvrbeJWFsGLvsDiwBrydixTcRW
sIqAGRh8eYf7MixC/reuguYSIBRmhnRQJ8lXkm7pS/pBuYA1nsXPN0Y3zW8tLiX2
6qFsDwwkzKUX+FBMDd8UapBxziAen+DqxypMDizGEhTpPsp3TyA51x+5dPBuUOrP
0sCCdIuKBbAWCOgVyVX8urqCxB1S3BWh0Z5sCCC3A2Wj8EjtUyTGN+fiOI4awINO
076+JGwJPiQT+sba2XRUg/WlCpLatayvA+uRQq2df6JRmoc1qdhx9rEchjdyQ/UD
fa9Aoko1XtOlNm+XtciPMwKvxi8YgTa5/ae8MUinNV3vwDOJDQfrskzkVTVjrZbf
qAlsDGix6LHxNFHTdCLeIQsBF4CKvOM30PUrPEiO+OJhB93wwou1Y64twZzuHsCu
avH8mtMJJlyML5pkEtXIhGWKUlZAbZusTX5ersQl6Pm4Y7IPdfR1IHT/pwKUHtLY
+SWpEL6ecc4g8UZm82rFZotZUUQ5Z1fA1iQr1IjuoBOyN5Du2ld7PikopXth5Juv
d32C0hVKQSV+/gLmYLx5nb7m87PKTqHzbHUEEZOtewZMHtR1a71QNXQq1p+oXhfh
ZrU+iEZfnwWGv+Xe/C3CrRO0+LWzs+70CGhUnmHtxAg7ZqJdV4OUToOXDNjfrWsW
zSnmIPCYRwEKPOaR5SoL/H1d6E9qCOTC7jSLcqqOiCsOfREpqOpS1TFiSCMGrkf/
DtRzif70Eo2TWgX7CXNxM+fuC8OEfgTL2pH/iqm+LiV8zbnwB0eLu/T86bFR0pTm
88g2C9p1mXpgBwdaYAyj5OVIWLODry942HB8f2y56LYHeNZoENfihOjAeuiBOeG/
TfF0JJJCkxRba1ncro3kuWSJBSXgkVrp/PeiSALBvKw3xoM+VoNK95oN7svydXvT
QiQe1F1pJYcnWZGTyegAhbi5OK5BTSnzSPOPD7hAxKQMHDmaX2s3Drh2wWVmxTbG
qPn41Gx/PXyVRLwTZPJITtcRNmGahwG40JbIWPJZ/DO85H8up9YoVUB1Q+RyYMQ4
lf8LErkvkeHOINyX1/V6wKDlgGdbKWV+H5J50184RhyPw0Dk/DP6sG2XgnKXSI/8
Z9Ta0AeNi/ftEiPPDlrHXkU4FusU9ifgsJSeIrFgA8TiE1xBBxDqB2/KRTyMblub
iIF0+yQ10I25DvJf0qfYTHMnaI74OCcwYd9cVAL0djhE0rfr18+Ni0cWneRNG6AI
+NprkUWWfcHEWN2wry2/FWMGmxocMxiOK//KWpC0vaWIIyTGfQEjB1hMEI+jQSN6
mItZXVRSSe0WOQnN/wCzdOpiRc6i6GBWBLF3RM88iDufWOqxpoyqwe6yEf2Z9wnR
HQp4UpcMu124x5hfdABX3UNJNPopT6hOHngI8jGqrM7mHQyIa1HKe2wSqe0DYVGR
LYXntsjbWPmPTmDJ1gqBeOPbGq3GPOMAe3CqrL4IwJPkwqvu1Bs3XujWxkjzERns
Dxon5mFna2VH9iGxUJmqqcfr0CvDE/jaXcmptEy3Dr/lS0KiulRt0D0N+sS/faAM
rVlQSaBPKZIf7be7Rv2h1sezLSOW+5eEwm1w187aoAi9CNyL1MKd8IU1gM9bXoI2
l5MjjKxYl9QTW/d07rtbXS4THx3rrIEXMvKu4cdsXDmJkcnM8RYWw0XKVD+Trkhf
pL6ll2Omx3OiGyO5dhtEc+1U5tfuND/ZlennYXzW/m+YlCcGDPlS3jndl1tw5aC9
/9hYcWKPenrPVH2WwkODVlxSwNlLP4zkQf3zPhtdzxTgwvGO6mf/ty5xpMvhA+ee
TA8qje+8sp1dMNsv3nwzcIPDjn+n+7MdGiAr6BEIpbTle7X7aWiGfF9e4us/9Ytv
ruJufnksZ8kjkZV7SWbIDLATmg7HNbuaG6VfDGeIyJFf+UyX4vvyaeJiREbI8apN
D/XRECe1PsZvf7OF/HI05rg7+rlobzvDP06C7QS0zBHqeksc/8h2W7FaOu+SzEo2
ai6+ppInBDjKIq0h/smnzQhrtM8z84bJu/k7b1WpLAaYRsiNaPGdpcqqc2sLCAoD
49IPh9Exy8tokpqtl5DuMBG157vLS1a7N3ohX6khkuKQ7k7HXYxY8nTNDBegmJs+
1ZMIkiFLXB9Whz6068WKwlP0P2kE4wi4dvqWkeViw7QssCKNlZwYJpXqd7OnT7On
eBjl4admwi/FOTwUNy8SYTUa+TtYTrXkl0b1VbBoBYRYv4eknw3XFZ6zEz2LxG7h
v4a59l+qopzCpKpmmj/yHHY1OXeO1a2uQXmkxkXeC2K3ASncGg4ZX/y3KEbvXNCw
MSiz4fdPqCK3JaP9LSgYVqeIqhdf0ZDV/P1xs2k3WnIzdXGgH0JhZ+76HG5ivthB
HCbObFY/eYMkFsGP3pe721Juo9tlrerqPhzXVrwh37z4xLisj5xkWFtxUexZ+AmD
/39YbohDZ9r9SCuFt9ts6LHsfVxpUazCMBHT+F8LAH8ypxQv+TXdASVKrs0r898u
IIPUbEfDMrcfOGwI3Ft1wVemJLPjjr0rIDye46diTeBdQ3cBL8BplGrHJQraCn8K
4hzDxdKboxNggn6ecZhH6Np+MC2vY4UYisw18iudewdKlBRTYtFUO2wlu+LFmptu
KFSbPq0dE3h/J6bk94tKPAGTagg0TWVakU9JUq+TtHpawQ82LRup5IrF2erVLfkr
L7gQu45JNCbi5LzMGBTn/rU807Tqg37fQYZ0VyHjvyKjDjG6GRhbxLlWTKPWDTLa
sY53qrI56os+n6/ewccFTK6702Hfi8tG4hmydHBn/ADwsTOjO0dyAd/63B2pGu+Y
4o+PC+3cIAMd++LF9c82L8B6XiTY0XoWLaUABn3+jRoe3lDbOvBzhL/YLnmzlq0u
Xj6NocpgRSXIWvuKyDffC5D+M7+YkVnLdSS+wM8YHg+9cQDjYXORofeH7O0JMdtu
9/E3IiYe/AW5c1ZVMHbDktOb7InQ8d09gWRxXBOFE+mSpf40JKapReyNN52+SWxU
V4GKm382CGAojbOVLLuEGLgexo6ZY+K0yQvPxDjTTFsGjdXw4OnMP9fZtOsuEbYS
KhOtQkdvs8MK9dbnWRamM68NZJ4PE4oieIYNuIf3Uj0bmQrs05RedzDKNioDpsf9
JpK0vy/Ji5lAQuJUb2Uy5ZtEDjeOq12qkgmuyBBSxkLKLjmSRH9JgomAgUHaqqcJ
Fy4o4b4W56UdWsr2DInst+KmaLhVR7JxfgXJEBLt8Dk0uEkZo18Af+DdTmkQp3S1
xpsTKQsqS3IT7ai02lIXAYrK0No65YW/l6tSr2aj1ywguED4ENzxz9ILQS7NQ5UE
sZ4zSYhMt6S7ozpNszzV+sNwt6tXLd41xXiQiomwxwTqbxw/2wV2IVgcE61DRl/Y
D/4TEuTQmGxylUc+qvow8j4T+Rcplzju6rF8EWsOplsKHXCt2U3W+H9g/RNKAaFp
xgpAO3xHzTtQzfu02qKTOk/3RssKGkSUmiaEkPnN8NZA2qBIjKALewaq2fif5rMr
MKLyW7oxNzPSdG64xchVMgNwQ4FtGskX8syddgY188mAYN+Jd8fDyMsSvDI38e1Z
2MuhLlS3h89Oh9R0BgcDjNdpf+yua+VasC8w9MlshCRqEgHk56dLJo67NyNP8AXI
f4w4v5zF7ve0XRGLMBC3YKcNy67pVv6q5Q97Q7LD5Dl9vnqwKAUsJV/6frp/z950
utK88CJmhEtOIR3hhh7jkRJ8ZRdzGiFwcWduW04c3oim5mX0Anju2W7F0Mb7keMo
tcXutlDKXIXtbAjvE7cwdtFl0x2yJJnTRr/MMsHXpIES/L5l/PHwnDu1Jp3ro538
zMhd3F4P/R61EJK4RAT88D5E8WfNamCSstUXfLKZd/+jgJeYoPESeUB7pdy1zhzt
zX24UtGqg06dqaySo7qW2i3fHGxxG6Lfd+CK4L/+l0Qmj6WlDvOmti3wbvdGKioH
Dy4862EG2VBkZEvnRQQVDuMmQkXZiaXzUbWWpebcpuxv0YAm4J961d8rn1Q4Pgj2
EmTHQb0PNvV4PNprFWCjxMaGy2tkYjNwjmoxbTRtPS2RocXGVirUCqSkifFCaxDF
ukP/7uareb8nqA7ijgoaAY8Ve3dp8NlOTa6DRerz+rCjy+fcVkjHxbxo9cftMbxp
wkPku9zK3keRpr2rCPCfITpb5BK7XiblEmZkl4nM0aXfpuTRhFzSPfUT2TrIcSop
kruIpzlxTvQ7EjPHCyrAWjlj1CNme0Klna+GNdGKKQ28+JCg01BhX6+SZoJaPe3Q
3RTdtZPPXylinRbuagg505PYWz6hmJNpl55ai7crD+K8a+Ol1cswOyuEmLys/gH5
84fIfuwDLq9fD0pSLqwqdk5PJnqOkzyr2bR7TfQgAeMydAWoeD+5DGy2ujd2M67P
eXJ0+ow9KfOj9iqKCYh4R+E7IWxklq4o1MhEq8EuFC7nplXupcTT4l9XGdBv8p7c
MiO2iDC89Q2MGVxXZG+xXPVXDYrSfSHMm+Yu9HdjjGOng8QPoZ8bEaA5C8Eik0Lc
Smy/NQ7cf4kIHsG/03dEF4wzwgNEKPqw+wmWCLnqDTLveSdAr1ZBiIJnpUPMnsxW
GGC/AIfoPYoj9K333OVFZC6GqfbC3klQqV/AtUsY3G5j4aaEz0eWeyWJ0hl+WCVr
H5YA/tO6qQybcIq1/wDcqrkaamwggjQPZZauMCo1HJs1aGsvPlQAhbQnMQskHrHT
4dabgQCoUzCEFEYvy2xBVwuEG8luXCx76d91KsGpanzRX04BzkShvdNQbmPtxoMf
aM+JMiWmWa/g+1dZBc7QiU7DKmme7GkoOcIOO3dMjpUMVb3Dv064eR5fXEyFvZbN
BPcWBY+0GRzYwKWLhqin5EjNmKZVuFDPjXcELrtyrjnLZ45rN1JgosxLnimxpSTR
4k8fo86deh9FS6QRwigoajABx3Kk3ChTjcrPIRi9yg+tJ8Mhnv9LesQFaRaN3jAs
B8XUNrwyAtx/F0EuXbJdoJr4ZBwbl+Psc63AQKp7X/og3600xy+zBM1PQ1/xlSoF
58unegpDG9G+0kwF7xztdr2d1IYlaW3x/WYH5nMslusjfCoqx1z6GhplXm33YsQ3
CYGlDRz6a3lYyBWxB73SRcqr6SIB+K+aSzi2j9/aw4hIHkqc6rr2I+VCxlPdPcFl
oLWQMCxIu3yrbk+lsgDVx3U/ZfKbXwXUe+n7AsdZwEap/pfTWPCwUta6jTgHJmNE
Zo7rGzv1dsMu30dIUknykNTfUxY2RYC/+qXur7fBUwzTVcbEbVFoonpWPRYrbqtC
f03yaZdhPQmKqMIgZJ2BISQGnXgxMicnuSZ7qBaERj7SdMd3KlHlbqVKMZ8+mOJz
Gz0au+YTMSPADvTheSL4tTZBoc3krhZzbO5+Vi5N2A+tGzW5CqrWq1YzEE4JmuJi
nAdHuSAMPDmGVZvzIj2Vzn/DtmgkvUVRAFKpVX9xbn/S62X8ovahL6kxi3TxPK3f
Ub8So1NMyEV1vQhUgvt+iLdKGyVZ86X/mItDSmtCUt3Er+Ot+NvLR8MXhHKvNpzu
rAeqoG4JPz0oxdUQImxDZSbsRp0G1jNik+KEDQGp36JedM44+ptK3NufqOvZ4DQE
8BzctnQmCF4GaOwmdnN1GMpIqRW7VgHrSo17lhXl9VtaHI62L7Ls/y9yiVvEBE6O
IBEhP2/caHdUkl6VbNmcw7scjVtVAPZ6XGCK+HyO74/81WpFkRMEu1w7Na5TIUxY
vbu57+ZbZHzMty312STmGsRxKaAnda14vOv3zN0b8dByIjxz9lvXX2RvNjog1DgF
pkjB+Igdoyzq9PxflLvfw51tE5ug0InarDCqMqf8TUdoIdCbLKCfLKucEGYbHzsi
nV8fSEyp92k7h1aieOoi1P7tEWD16w0dukOn5oCjDqOWsRPA2QkNeCmR1z33v8P0
EpLqm6g4bBzQu4hcOYU/Kcx+otQnn6a4m2iEdGYAYAjtIprukgFn2cdAseR6OfXg
MdVKpSGkr/K7QsH14k6e/K8Djvf3cLc1bEe+GTwH5dYIlQaEr1v0gSOwKkuxKpTe
KaYQR+bmBxxWHqSEM78/Mkhn80ACbez1LW82AJUZfyaVpAoygfphqvzr4NdkmuVJ
6LiX/Fl95HfQIFUp1QULaoVDlrbdnm30R5kd/fPHplUJ2bkS5saDzO7OKKSgH6TN
t3wMFb+Xn9X/3m0L1bx5NNq0C2004iy8qoCBoZPwHylBiJSCPhjxaoZr92cU5RhE
iXg11nfyThODgeEdRyiYfxjG+cCw7F0phkNVBsV4SR/Do/z9R3gfHcPokeYJlnCh
GpRlAzpnzfQnDD/Q/6/3kjHrLZNoIYDNcSN0V8Fsw2uBMx3oGJocQqnHUEYi0U/O
sOlUzmHMzZBwn73Z73ZjTZ9zALSj6m3zd++tvLdy4wDeh3htTqUlzAtTAh8F5d8x
Vv7b/vkjzCKvJ2TQxnzzUvsiQdLwYB4t6Hb4MR84W6IP682S5v739e9Ex4r8SzKw
rTsx22zhonU9s91gdWRMruXPZ03qJzRuZ/d9vV07vxAoDq4ZVRxglHkPO4yVCtyP
6xBrrXKuYid0VpItkslhJcg7TJzZv93GvG3z7ssUC5VU7rl1VlsxIWQ35y/tzZur
pfzpL/rjrGDAXY9C//ohUq0sJFI9OT3irfXaxZCPkOlGmUPyKPCP6Y+AIrvrjpVA
VbFlRBuWa2ytqjRsfMycUIS49r+GICw8vw8iq3ySi8x+rrXxivN2B71C3Iipg3mp
ZwPt9cnLNx/6CSF+U0qn9BxX40VABnCiqr4vqLpKLe9ilcyGdhk612SjCA29FS5f
C1g/9hRCeng/s6dO+98pIO9dtwLKkMPRq1CahidwG5DeTSafI516ToRqEwQVMl5r
FL3utCBmZFU29SLA34Goo0VDASSfLdwDhnclF0iiktgMcUv6cPw2sp4ZLaqrJSdf
Y50O+2pheq03IXuDKI2Qum2Vvq9TzPNmmoSMGf7HBAzK4IYzGB5QGl0vz+/l8eY5
dEBGnD8T7if1Pb1xi4ugVIEO7RE81d+vfLWiLW7pYbEp70juZcV/EBrDH/W1C+hA
qtULooaxVPMixfgLsejRqB+5cOzFY9lQAlLtVyMPsZOJ5TWuojm/1KEXYUGwUpi5
QJBx9wUyHhym2pAgz/YdrZ5ffUK3x61eBjqUWcB6si2gqdjDg14WPSxYgVv2zQol
vLx1ZV5Ne3FKryX6uv9ih8IfYor1a+Vq+M7873UTCDNuX3eHA2/X9YdOTEHsiPqs
CjoIPQIbT+s/eNtoj6QOiNegQsIlMDDCmjdHPEnUX8jKQKwB65Bcd349Jb7pZKoW
crSsbFRMVlblKs65hZHrYE1F1AFCf0Pmderl2CwAzzzcLO0KpEVAKn1Ab7t+TO2e
Zf5LpucPuU45mm1cgJ6SYB2eEs9oDe1vyoUSUNDtIJ6tXvv47w6UQkXNWJ0RfKmE
W0FWWypAFWZBjVKqL9g0eKa5uVNxOm8qU3qCvghihnfMuypABXcp/UK7Q93glKkG
hffdXcehqdFQGfYgdeey1bnbLg7XKgR6TQ1ZKyyEg/YgIcSUVAHGMGIbYVJdqW76
dEmYVEGLk/g2NKHXBiWqQ6ca1eU1hpHCSH1hFC3MlJ71tjA36Dnkwb3OTbvPrG/g
7PisvdsYwYvH+gB6ZCX37TKqbPFZWKpOr2HUGg1PowkqinVTkfazrODU+7xiX3Sm
rafyOa6iSz13bbVBULhuTMGtPE8AOXN5qNiaO1f+mxdDkpByGbo+laOdMWqKMOEQ
kmw2F3xRWNEIVl6cNpMnx24QgsW96busLWZfYheDIRVlylXIT2jrmbAYkrFY5fde
761AfalFp9REHkF1shsG15qhP5153xRjXhvHL/HhxxIJBogZQ9WjWHFRPcAwVRmA
Gdkv9wTQXB+4mD5uertetsShwq6700+h6j40KWKwH/r0EpNEnixp3XYXu7XDVTft
UtJK3LPe37vEAhHT2Vv+can1yltdkoiSbwyirHHpjeCSRBWFELm9o8kEsZHykEP7
QWVqCLZ5DWIuEqF0o7V5AGiS02CwaQqFgw5+tO8HBB3EKblahiCzF0PvLu4YKsXu
XxyXteyowwj6lXhKWOlhEP6/pQpX0DVongdlE0CNtmANfHf1x+E5pi5jD1Z1kAgl
VesBCpaPe3zP4gXjsHee67suDtEj5nS7Ezpvb71/rxJ4puOeE2ZfzK3MsC3odAqR
+RfdKtx3o9AjBBIadCF5c59497w5443QawElzDSaaj1gcHrysf43flgdwkVN0hXW
TaF/WDspe3iHT4S8FsZHYRCpa+o+EbUPPQoS4g1h+MCqkGelamWHjlhQFhf/lwIA
pv9Peag4XOX7T8cbLr6QtjtWmrg3PlaavARMUsNtjRmkX3/fe6oa1ilI+AY9mOeO
lkuWZ4uyOjkF4Keb4sNzOJhgoj6+OU2v6d8Hv74YiQM5cEmJASXuNo6Wm20Zyo/x
dYCX+cpHQdM2P5ImXlS5qzUCPcJU7IcIsEk0kc7VWea/Lry/XmxMqidzM6Zus++e
XjpqOS4Gged+6THs+UbzN9Ey4KLefCl04FZbDikbZnuPdf9+OA+roC4v8xioCule
/hnmUKwD6Yl7S+gudioi5FUQwnHkUSmDqveLqcE7SrUIW7nLce/RfEFwTgnQT90C
d33srmySpiKAm2UOBC9S8p+4mWYrydHCNkp1UDrgN75f6c+aaPfc8bMIlRQ4ZKT6
Lab2JC2zvFal6jUesutSBsolwuTQeGXoxtZH5MPvfuBgU6WSXmhfYxK0vE3vKo5s
A/5Uv5eX1T8iiTkq41EDMbEBMJFneQtES7mVrZcBE9d9jCbNOee9oJi05Q3cB+Qu
bJw6Kl77gheKNVZ+lx5dTlVwGZrtkeWcZlV8frkQNscCnINE89Us2z1ikZO3kjLf
2ue7HhBtE7epUQs303+HTTP189ZEfucMKb2DfpHU1xsqEyv3WNye2YgPP4AGtgro
W6hmbCSj6NIBYFdHeJn0RzmJctep+LkJrdUmkZRFPgG7zpXH0Hzmhg0jk8NH9I6T
QEz1rXJDFLJfiXXd7oTFzBJ/HLMnV85KtiC67t9apV3jn4m5rztO3ZPCPspDJu1J
e1zOj+U+vGhpGYWNt1fsu4WsPhzph6h9q3tDXtOzIRi+8we8OHBPeeNT805I6Wz2
m02/vEBqQsZDUMG2B9mY0onVRbP8gENpzLpktyXcefiCExreti6uQmpi8fPjxExa
3B9+o/R/o6KZXPa4AUdhnRSG66lc1VxidHzyhlS0t5EM1WU6Rwyk87mIwwcyhUl1
KsQFFoitVKp5VOH8NE2ALTqfFECN0xkeDcsGBFLoRYsdqvQEvDbnulbi0tgyVNbn
ShjcA0sRNRbDb3s+CsViJEaMRHM5/yT/hW4gnjGdaugvwc5mzT9VapA+aQBX3pNL
9JKgtK6BoMxb2opzgB0zjH/WbAixswJefK9hDC4zLrUEn76gjoxRtuSdMe9cuHj7
yffgjkR9dXLZXQZFVuTPPpGPHQBuHdLfE+7gta4EHhwgvMhir0rakznZTuZSktby
hozvCcAbw2SACqDob3vpApBnzrzpez18lLqzf1G+OqETtAjjkfdyv/A9kgzcHILG
2fISWyxVdJTQqAe88QtXDyx1w7BpqSwkwh8RvdPV4M63tEDBpRpft2G9KpEkiJGD
JptHvdKoSbbMyE6NvKI4dj6PmJ573WkMV7hq/gxz8Dctv0eJTymyR7CPkDNqd0GR
RyhAaxo4S8OI7Sie0QgQhpBnGjBKTvBLvhHWpShD+hF5AQgfNJfV3jFpKQNUft0P
mD+Ir5Yi7PI8JMsQZiHvgVLARDEy32QnLz48pEWnPUckbdyDLhVjre0P/zHtICO+
/1AsxvGUbnr/Ed2gg60AxO6g6dAfzbiT1A/W96jVzFPAp6fk/5isGzvzkVM14i6a
TX3oG1DRevqeceOjwyK0yjspMo/PL8RclL2WLZazjHTLxubt/HmltKmw1zkwrXSx
z07E2QDXDbMAIcbsFesXYV+NohrG8KhPLi9cwU2Ro4GkYZkLRVJPbpC2q8p2OZ2m
cWt6LVbbrd6KPT9mbgIfwDaQw2zwQtbzz5eDmtwhZelMKIg9lV9m931cJUvu1faO
M3g41L42ts/rVKeDl/GLtqNXr+FEIwm0ROeNI3G+bydz/nHIuGBkc/l2FMruTMGD
/ZaPhbVYzxtJLbsAY5jExeWmjDUc4HQU1BUVLZ9WRE+IZL0EZqZDsPUyrnf3jIhz
l87vYkiBrMwkXqBxfjjmfU11gpRrG7uSNJ08YMnhbsL58h8bJY2mJffO7OIblA4J
ge+t5B5EMX0YbiESy3Iy3Moe1/z7KwXczFPBVYew8CYifkG7nZ1fe3u+yAKUFVk0
2QOlR/Mnb/+sAfIS7Su5IFeo36ba2hKVYg8MYfwe6EjZkFMoB7yqzga+ZFcf3XCG
2FnHufYhym7FxUmwL5J5YXJY9eE+tj1hYLkPCzUfmB+NWfzbTaonWmBUsj9PZRfe
jKsgYDUA9t2EXcH4/f+YmCcnqvfjvFOUOhdJ+DKc1pfCMJaOrqqSRvnFfua8VPVh
HG/nYiTf2NBIrG1WB25atH7uqSWZvWfckgwxQd7J+DiUdPyb2pD5mmxYHwFKHm+/
1g5FvqwqsJrsQFVjNRhwpufhvNgPnRsgzUmGVtP0fbaLzXWNsbVQpUu9CSwIK96C
OV8W7GK5/tvFGM32MufUKCcPjxAw8Ds/a6cbZyrYU6bnZlp/erIShr9Q3NNq+Hck
nViQQAkDXQDBcmb6MVG7XPUzWASEv4NItd9e8OYkgthvf3TRVPnEIJEgaUsY0DIC
ZA2HDPNesYPw1sxIz9/Pg7LTGDZHMU12M7FOX0tS5xh1yT2qKu/8wi3zj8v5DXEK
zK99+aP2Dy34ckMo2G1qqRmaVkNX1CYKlJ9ENtTySag+EtVzx9FOHRrQlsTQZtU/
AQAL7fYNjAf/aJsVd/ynD3g01homwEqublmGyhq4nfVPw+3ox7v2dt7nMDTuZ6M9
KT4vXPmMnZWWuOzsKixLGt2WdzkKtt1K34gwCgAMAoW5ACf1wlJxihmRf/8e0Xx/
xrGqOLiVgjdF3X86G1GhGzb/EpM7xpdy9KDlrdOYibjeo0AoAaXe5t6tj9mzxxCm
2Vnjo4qPn1zDBcAtnqQQB+3HBfQw41ZjOVNxUa49ClmEZtSKLlpg6UOi1yPX4gOX
k8CM7VOs654a7qQozQ5391uowd7YeGhg4gJTau0NoifW2ZP96Q5f+1LDeQuQA3rQ
FWxJb6bz7haHdH445jnARRlDjlNVnD4F610Nh9kPAulWYQrc2NF2ie2zAUypi4DB
DQ8HYsrL7Pr3GWZRjvRTqygL/n03g9AqXpoGwW2mhZiTbJM7PvaSlZPs+isFXnR4
P2SKacT6JdGMkTDXxIEcODms26yN8XxEnrgcDGN8JlM6EdIvsaRt6Uql2p4XYtJl
VpxBBS4qUJl6MGtIOUZT6j7TclddcnaDzM87SRO2G8lToGjvvFuJ5wBQyoJsi5Z4
Z8wN0nA9T+6MOpKag9//sj/vJcfGZCvJZVkOcqSWlEfXEyHc4OSiMBQrrCh7f2rr
vrlTiUPu2M26PLpqz/7oay2wSwxf91oNoP6tP3NGkEHSkvAp6XkXgLdSrwcji91m
dRkfuPcdVSvWx2HjZ3tcR0obRdQEGVNgILqooouW7o6Rp075PoOeuDQZl3Z/iv6S
HuWz4XUNeR+VGajidgK2o6b5SWKSK36sezduXBji2UCFGR9ZytfTdzWSNW4RhHQC
MgiQ9lhur+TaWxyOG172MTgWq1sVWijUYmU7ZTceoWTKXLsbeRukFoJjOT7eTHnY
DSD5sQdh5HSAYDtla+u10p/2qBcknpKROUpzwAI7S64zOa6xSCT2mYgjGP0zSBJW
d5HFCIf9gTArP6oig+R+2BH1gOH6fSFigjjlQ34d4LmkEp9JaBAs92esmCMEMF7Q
xxokPx7glMhehOqC5/p4qkmjBIriLa8Fpuho0Fx8g8gjjGdVXCq26t5On9kQ6434
+s1vnqT1yIRqGe8XbGUv3nlRsxA45C75TVAfW0vU5QXydeKG4W8gIU+yQIIh/ZvN
HEFfZPBhSZpskHKeGI8Oe1ymun2BIlYEknMx1h3yQyeyDWarhIk9S3sD2pwEhOQV
o+F2M3o2G2iJXD3+dM1xUOzULib6CDeCeBiA5cLsPMumUiEPdUXEH+uKORpK04I7
1g48UEBNGSSqbvJxL3DUkhmjLlj7qk3D9zJqiXIDaJnAjpugySPD6OaqWUticV+6
dCBlhQgGTMW8f2egYhGG7OS7qTa/vzTURgcON0cYyhJGB+M5SHp+3VFU6lPtebLv
AEjnWpgWx7BksxUUgGEXIXqIkj1+R+uZXj0ihhB2eKQPydpzL20gWOoAZ7sfgiuF
iM3D0GpfB1Wt74hm/YSdWb+4WootthnbGA891rNfiZN8I0Oe2mt8CBZVCo7QZnkz
N3xHZ8w8YAqxJS9whrnjteadcF+lFelS4xqwwDW2HWcsRQcK5H+tKyjnTyx8bPaA
mgyz92AnX7870olyR6YM1Fzvq41sez9q2TilDfB0ChjdF9pAHHNXzuviT0u5QRsz
YBKAQocCQAaOkxhimaqgztd8V5L1ZENYu0qqHL9GlR9EHWZyNt6XG6x/vxgSGDMO
ccIMpNCN7UTFy9A5hKJCpUHWhdNqQeOppETeUFlXaCYcQwAysXA9YJfjI/85X3FW
PpX1AG9dRQX6o+Wi13VhVqA5JpPPBkVcGpiRjtdmfucX+h4Q6+ojyO/z7xrS6ts4
GnZ+hND09/YreWDCR6RoAiW6wTynEYOm906zCPvq3C0S3MGUsjsytfyzOtZHi7l9
KGikLpy1wGhTFw/DyqeFVuq5/u+WLMFhSEYVCDZUQVW5gJ0/hpiYQIQJfjEOhUp+
1l1Wtbl/ohjQkV4dq/Yp/SwYDWD9/EgryraICuv3b/sxMWC6wB7erTggwmgG/RhI
OFzZVqOlEd+vHoYFEF0O3Q6fGvzjSRDrdLmBW5twrX5dykoEvus1DBgbJC/fEwRx
0yed2kqKWNKQlyTQjJSaVeB/+kROztDm3p9qQjx3hWa/s9Wl1c7vMZdnReNVYDi+
ISjeQcr6EWku60o6LKvWMJ0FOmA6w5foCuyQqV9IgZVuSOy48QjzCj1KN2OlFqM2
qgudtEoR5qlpuXUEDc3tVvRW2Dc8DRAERn0ROVZhn+bQOFOWxZIpCmrtw1OKPRSC
Bgl+m1oi3XfAJQA6dwr6/diz398K3V+wv8+r9rQFENdKGg375D1QJFlWjUUwC22S
47DtOyVqzGljlmmuZDK2IgG/nvCi/JgD88/LJet+iqFn0gdCChNHGFWZOhznGt0x
p2K9QWQs4HCNpr6AJPvzuOAX4BMGP85o5fnAt4LoVdOctbTht6KK7us16Z8A+DBR
NAcREvoQD2bFJ6CwQmWZ2ol1PjkxOucsnDCN6H9uK7AgLZzMigTM6c2izVs8pLHZ
7TdxYnayc0Jv9DWCGiKIafT79laTJ7QTSX1EzR8GcAu2Agb2RwUm23P8iKrc0JYx
BWVIdikJK90VQKrEheREqX+pxfSW94KOCbg4GOyTb1RmS9S5IdFolyE5ml4Boe4E
xxVkkyPSD35Lc1zx9MpG/9lHioGl458MEb90hk247lK3ZgwNvSLnASGf6BP/mZch
7YxFRi9C87bm0kC0miVO2KY+wJBkp0E411UTNGmVNGptthZk8daux1IVaLkcsBLL
gk8cddHgRgnYlE7LjMBOZ3A6oy6Uvq+OpTEqdUu62enDFFwzHQmXhSTJeSDMcDMl
tZIsLY5WqzD/z4xd2SZ/doR/3uXGemL6PZjaT1YE939I1XeqQu3G0SMcuLpzWzel
ppwhfYbZRsEpuz9Vgb29nrWgMclXtb+uLe5gjNVkrKoPnzNgs2LemzP6dagPmCj3
ryzQhysooZCc3V60iMsSgFXKgGR31o7gY9ncdmAZVlvGYVvy3UamzsI40+fwtW+q
+xY7FiZMEKwTvRNG+xzKnQvQGm4UzXq8Gjq30RMyba0Oy8p67+EjTurypgXLEGei
10eEUilm0hidxBLIphAKUkdWKNPGtCVZxB9FCNV/ai/LVO5wl1Dy5S4N1lg1VEdx
6UucBFulEFOrX7IiS8pZoyipBu2dXNJuynXcbdfC+z9266qW10dS0H85V+Ye1fuz
LuEKEAB3TALVwuQnjDdOKlJgmGgf/x0UD1dtyU637Fkb8F4y0tIx2wsd/CJOpylX
y3T+dLiHurEfPlCWRtCuBPt0t+ycEDrSJlgPbSbwgFjJjUp93qB+vOwIJ0s9uAUc
ZrGjmomtD/Yc/FfZ2dzQno53Nt0rGmPor8SeSHSAmCic7kCn9JiuWARJhpnFY1qU
XZfa9zI1VLaobo31W/oIPF/g7Pc3FDrKcDjDPbwkO4bTtLl9rFf/E4O1p4k1pxgx
cbt907umGsS8j/i1GYETpoQn0tZOe+Zo8Qm+53iG4D6GTZ13XTWdJyq02wqUJDLK
d8Wz+Q5v+xsclmPrIv5hN0PhhGuwjS0xHsZ1MkKCVLt5Roc4uqhvrJfUHunovoc5
3vXCQ1VNFVzk72cxn+vuWjEcXET7GahaDQvFSh/MoLXfR340H/OmnfNX7auCS+xC
7K6pH4mAcv8PM6ERMFL7tmSTnmc8AC9aaNPQwojuLlEy5FykYMYJBLkNUUzDMDkw
Zo+Ffb009fwp/mIiVDbtjrsR13+cqxa0KodC6i+zqYBq/B4CjdosQkPPl+SYpccg
O7VSwkfEnn8oPQIBCXLR9Nx1XGPyPO7xu8T/kwPuM60xJtGw6/8XpWaf05T5Hwb4
8LS/zWlhqJjRyIW+ToUEqM7+KwacvoZoNthfN0U1yhVBzyWs1tKIF3mTMr6gm5O7
7gBta217xix7tUz0h41bcL54KSLwAdjpL1V5ldrItTrD7mKdrlnxiThIndb4sg8T
jY7rvZlX/d53bzGZUJc1hhUoWPF+aMe18ednSB/pJQ4pzu/gjdrATLMK3J4reWGc
J9YWbfJia5g83AioaACv6lpbhGrvvvPhTLdBT8M/PsrJIhD/rngAFJtQ+9u6ICRq
gy/rJgh/V5LMXV08eA0v13+bKwyuxgRyeHlOKCI0sgc2s12o7JB+FHF9O8eQFQZA
KA6lyp2VSA+awqWgz2rqqbP6EX9f/wA96x0XJUrIAr90oJD8IUQup9HjYQakxWDw
b9esJvywT4hLb+wdZvXHGuvkRWW9aM0stDV5i9Dr783IK3Jd/w05nAf339Ru7uqC
FaSHwXdgDvsgO8m8pgmO9WOfXgmIlkWknzCjyku61mYCxTuIH7VPh4bQZegdBnw7
PW3VLyw0I5/wuqmYOkp7rMVJLuZYR7xhtNGWzh4twwfhl/VXy9Eyn6hLlT47tCAi
opNe6a9UAN6iyYY1CWwZtad0h9Qr0jlWgWWUIi+TkxfTjkWsj5L/q70ms+Nykeul
G9iXxwXjcPXC0YZTIFP2MENWyDxqCygJBYDIY6dOKIeEsgglTtM3r8O5Vd17qC/6
Y0dNCiJuio+x4ehVWC88UMlF1CwpBxfcF19ex6XlmL/BFYB6x9JxEUl6+DlGcuO7
YX1qlLZ8Dtx+zwEUegQRLU3i5UDgpwpxbOsdIv5lO82Aq/BmgBcdE+r45HPyb8J1
MA6m8IryWTWqMDxU78mpiWKhrawlnB+vXmAqNy2E+3ZRSFkoO3HX6BVXRTz4Li2q
zurLAQ25QpUoQBhJ/dLjruBOfx19mysHp2hP16KQCgtg/RF27HgD7bXtW+MjMKZl
6ilGL/iCCZIKsqwyFBmQ+7uICJTjGppqqWgi0oLvfC64VHIHnj2kek/kHu+RgBlF
T56G9FwvCywhzVrv2QUBIdHz4QHLI4Bv3dlvoqIN8Fkd+PZnIZ3xRPjAaOAghP4b
eGmDLDA2ncuKBWVeMD9rUDrZcmelzhd+Jqh9RjMVYpXym+dfH8rgamGKlTjH31zn
1pNnN1/euIufySA0hx5lQNMESXhaUXibuT26tRKH5kwQat4sjguFhY/bPGVmJjxL
xFaslEpfZUKlKqfES0lLLr3zbscAn9kSl4Hx4RRrFKE/qNa3qcG6nwg0O99m09Z2
isvQM0FIB4WxwRuXqHTmDH423PVu3T/Y/d8txetDHSPth5vZkP4BdIjYy1pOiK40
JsUesb2dIY42AmOd/8RBNcui88gxZ/OyKZ6kTpKfJ0xqfK+o7huy0olYN0xNBVs4
+0cZXt6e8eIJ/Pjlf3qvnfwsrOAXsAZ8XqJOUEI8Vt9GljP4UOuLFBnvPsXDZRsl
d0VW+RVPVgTXGTwhypTL+9eCGmoyxcaZg4zloN/xRgBFFguz5JkAjW1VrMICuegf
iE2xphi5Yi+4FD3d3EJtiF5VfouuVat9Ib1BCOxyQfj40cX5iTg9Xi+P9w+/uOTS
M7s1eFHr9WTdagnsDr3K1ob2jipRg9xeBjYAS/YsSe0H3K1h6GpF9T+fa9thqVjN
3Aks8hct9QAY6hCj+EYSsqTVXHdMeP5IObsw0x9g22/D7EEG80vxd3tm7aGH4yr6
CAqwCdgKDR6l4R7DhW86Vc6R3zABr5SSt4Nj0PQ4IvgzD9DhKKZnwFz0Y+K+DJdM
Hl2MUhoHFj2Rcx5ECYuSw/fe5PtAP1h50tKG3qfwZGRIXeiMTh4c7/c2iqU9Gw1Q
hOU3W1nTQedzDGUwOC8fS718LzhLy+A4SuVMyWqP1hUW878UbH3u0XLrreYIEnEO
I9tUem28N4b+jgxPpJa6dk7FK9LHsQAid1a2B6JZ4o8j26FOXdvVzEocVgkybkxf
3x/JW421rP/T8g8HQzRXOMpNXqQ1tpp3Yp3YSxAADHV2x+ImzO5YxeohyqvGLW6P
1fLJKLHB9lT3/0DWBkIa8BDmL5JZQ4pRBaa/bQJHIFuIPayMdzio/phXaa3EXT3p
gRkcJRIoxQC4kAO8o0jwahjUrsii0mqypdn5cDdSgeuF0B/caJ4JO+qFf3QDtnsa
97/eJKzHQ6bjDrVl0MWpGvmzXlSE8XOHfefWEpqQiIHvdi073y7gvgiXiAlptSMt
/UbuOkI+1tMeaxASJsWHgN2xZulHTjPxyRlORUXidTCmoxtAOLNAHFnKRyX5aY/A
6Lk14JTl5wqVQVvEoHY2tMjflRtFhg/3U5PjAB5fAOD+6BhIVrdBl65mXStCtk3+
8P40UKZBSZEz7JhKuFOM7E1VCnKMOVVi1TmwAveLONPZIR142g7EyEMlsTMzxIRq
5Z/5Yl0WKiGd3jgmWLx21xLgAA0YAzmHZPQWU8yallUzzfY/bJBbPEAumqAxIZsh
zWiFzdHlTo3TDbYIMXF34RmQ59tJWNC0+Lmh/zy0WbcSLIMgtOFG01ZUraQeiEOY
Gz+9rVp1hp47U3SBsZ2qPLg8x/CKxy+n7bqn/FnW/l9US+U9uJlbowYDztHnjuRV
IevCJrUa+9vANm99psskxaa1ko8jI/FHn5i07LkfeEvWow31Az9CetFeh0IHhTNH
SdtTY2zAFsQMERoU979OWPBhgE5mRBi1UC/2ijsBCMDiC6N/YtsfjQ05THjRXgNy
A+utc3QLjrCxKFXbM8dwa+wR8zOA0Pt4+XuEQwG6UBium6k0OyAM2CJopDFj2ovh
B4dip9NzfxwsblD8574Zb/qyHu0k0mNwlsnXMameVwSSRBWdKSr4DAUt0Wgm57Az
YYb3MfkOni6U7g5EKAPlWgXxuDlVNjyl4e8t5WmYdf8Oh8xrLyUQudieHrK2aZ6D
DjWWHxaH6kYgo+aym0/nCrUTXMdwXBQd33EAjehb94epGEztkpbSEbRVzGmear6Q
X3nb1OA/v3wOuLts9Y8AAHZnySDPttS2Rhw9hW3CQ/uQCdr1P2EGNfbC3RbGN0p0
6+FVGQLgvpx5uAYS5wSWrwmD1c5FuLKX3eJSHf5BsYXfZ1SV8Lg1kyhttD9ULwR6
77U7S5m7Z0dY/zOtXyRnhs+ZGtQ2oQEMYKpZRj65QUMZTZOyB+/JxLDQNXUxZ8C1
awBFQTg8gIyljt2WUUx13evQlaIAn/7R6gUGOiTAjg6J/bsR6IKZCy0dZRWyCwKs
82IDIvioeTGK5oXf3mYy8AqP+R5Nf2WTYAHgzMywZHihfgndnRzEeEk/y4AAenft
wGz/K1+NEgdbus+aoazqMBwzvkT30HFjuxpfrD+eqsoDZE60nFLWXWNxpqDfM1dO
p6xIEnYEWFcPr0hU/nZ2RpZgDlKBUUnhOBVfruijMDd1AjZBrx0cRWwtaQRCUvnP
eV0shn6InERr97IdCCoVSo3vdj7ew4wzYS6tPnf1Yrh37XgA8h+LIlTm4zlU7F2+
MdlHu8c8DICPJwQLwm1JxEldmXMGY0/3iA+2aV0DhbwRQC2d8Bi2bmuekogDFOG9
33qbSdt/J1ub2xr7VFNrxZ/fFYP5XP9v915JPiroG9W5BQDuvdODelQPYIDvAD7q
8HzhmCN10Q4kQIiPSym/9/wL/+iETOYm6hLCBJc9VJjTrWIY2Hfp6S2aDAeX4Ay7
jSwaUIh44GiNU1GzTxobkGUxy5xIKU/zRwKn6KLdITpwGjMy6tILkXKZ538yA25d
ZmWXSDClQx4UrvSQTSbZl3bwYWizW8ReHAs1F+wbF+jpDEZVUpIIQlrxhumBgAGz
bM7NXUndPUBLz98dgNoaDGSetN/g/NQHAqJQnbgZEx+o2G3Ik0Hgwmbq8Uti0Mce
mim/1YySvJEqNSb0yEsdoJrUWQ/7r9l3GT2+mdHzCyYMW6ZF2UHKOWFhZugNFonJ
5meCrfLMfLHUT7euVPnaqsjMBv4BfJ3+/ksCdtta/U+Bu1CyQKprXzqLujEMzdPs
dgPmqWKLpP2basGV9uCeooUzyl9SziASdzmLHOqQvCUH8tOlKJ7l5Nf9m+quENbp
+MHvStnoREiSPcBiD0+s5ibawWNbk0Bflt+vzVd0GSz+yeS5SIoHzJYj5i3Gex7m
OM04aHLsDuwSrW1GcC8EOCG3t9sDL+1aKoBQlaV5dXZI4jzxhxuCUMxlktsKkByw
4nzEThXjujXKNo4jwaUGRbRjHMIlaHs654GSibXyuwPTUaBeq1ArR7mTsxJygqHD
iyNXhPgnLHMCCiYxG06WABVeuZizEyalg+MARVH6pT69m7qrZkOwDlb7OBBp6RLc
31SiUpEAQd9DC7qXB/U6U/ChX6mt2NcT2N9Zvu6v/TRbPso7LEqBY0KS37GFwesK
EfdKD6UhrJzqzc5rf+0+tgd+Ybhos01+HvEFs71iL3mdE3tyTrD6MqrrAMKPRGtR
OR69CWR8yQkuvnOvGDR9RPFeNYX+KOVv9RGAr99Wiasstl/OqU+SnRlnscxJQiZY
rKQcfMtU1NZSdoUhkFWXwon9Wu1QRjx5IQ7OcI2DX+LDj9i8jkCW25p/38rJnjR0
B9pDGSyrnwiEz/2oCR7xdf0o4seJ4bsd3wG6RD3gio8SAPg4yDTv3Y7GSpwWKl9Y
pN65oiQT/7a1tb8KsyoNpXCCDjT/uovsQsiVMjcG49Z/Ss1Co3PKUL+cm93PDCSv
zSt5mhDuRwGA6VOxK+VhMSs6Y1mCbOO/0htwQkwy3UTYQgENBH6HiUaQktXJduXs
Wvn4QrIl0wbydEw1n7ybHJC+cGs114Xeu/Otyb2z0p6GjzLY/OzyaBdeEd6mdQes
2y/CcnsMMbu/1AEb63BjRDeT+dKQ6G1UDbv6NYFq8F2XamgrQzmYeLE6xBLkSa73
iTwbUk2WhpgQMyKvgx9qZStqSzM1p96MYDUhAkDpK434acqn85FKcJ8gguHj3dV3
yZ+wZ1EoHs8De69hrmkJEhbLE2ScdmKSYhTXclsZQa2KR0O/8v200sZMIt27a/fE
Crqh/uQSJfMyLDNyzK2O6mWjWf59cWZLHIadTGg9RI3DrS3bLsyrgh56dbPq5ExL
0fSjk9hMv55oG1+ZmTE0tlDlV4jrCGRCum9328C9oA4hC+nlEV6pDm4W9i59qp9n
TCoSzFN71uwdWI3SNxE5mqRgOekq/smJwqxIjHUs+NTRXLKCLcJxxZTC4wfmmsr3
qgGLHiSdvcWV5uFOF44MXA6XFaqqYgnyVr1jztkFcO70geWajPJjsIllw6OVkWs0
P4j7UzYE+72vtb0GsZfVfdyoX6fjfSgNNBMOQ4DLbl3d/UDL7lI2o7V9qtAc26W5
4dH3omYv0FE19FWb2yxhHzd0HiSFFd2Y5+7YlpMIhsBbRkZglg46bxLpnFs/5KcX
FUafFjtCRJ3ph0XONM/0Eopjh+/nwY/lY1q6KtFjP1LImTfF46VcJWLWT5MnyCwc
XNqFLC/jdcxue2v+7KCq7nTPEFS+9Na4iv0qpJ/gx0vnlqm5Qv4NwER0vsGJN0Og
vpIMA8eC5bXxpliuXkzZJjxyxjVwKj/s1olX+AmN2szTUSoOQ3tf3mTv0ZBKErYd
FAGsf/n17Vnres3aTQh73VV1QNkSzCibj6HvRxuyiqvG+5vGk4cBEhhKn5AtFFsH
lhjMez2RGp5iqZvBwdRPGtez+gY296U5RpGA8H6GtXnuDdzfEJspzhQlF4JrOHNw
cKo0E/wDjft2VDXXyswwfmGdQIvZNWWAqcxKgr6W0akugZaZi/rT8uKLcbuImAlN
1ku5/wJWJdprNV3hHsI/l3Y2eadElg7C4shzygzba9+sZ8yqFdmkFHTh6s2pAjU2
bnn8vtVojEKeoQIR0AH8ScAnPtU3WioUPq1I5tOdKrq9Il9+HwzoLcv79AVYJ0au
75R3isJS6hIrvh3Z4VWHGWxfDhukJmURnv+kV9B+SaxKozjLyb3CFP6dDfqDFSHw
1ZfYprasCKmm9m93kcV4+JGWR6DXabjDEgSvCxUi6eiI5xG7S8ed6+8QXKT/AIwV
9tCcQ+Q5Zj2TmDZBRNdkXFRvBNkHBbk6bkuEztdnirfXs2OPXC+jXrmYBwAQbSeW
50UJAp5JJO/jtjgl4/pLvFmMyAut9nN6+Ho/pHR6NRSphzMM7wK1l7H1aXDdxtdJ
VSlXRZBhjvcRNEe0weezaljlidFxN4W0u8QmNimOhXnbnyWv3kRaIeNLnQcJfWA+
plVGvq0IKF9LwNCqWxaje6T1FD14a9R9I6m0Y/jsgarl0ktu8m1yFnTtFwUhSM78
s5UsnxuNB2WMAj2KLKYXVWd960b/fwb0xHGK68saz5FjAQwpuKOXEY00fLzCCQE0
khuRMuXnX+xUSzy2nv0FadWs/PAtZ8zJ7T/Y9Bec78UgMFUjJ2dC2m6T0VEdBM/3
fUcJQ8eWIpegVfavubU4IVUb1KMU7bcIe1WAB9VPuyNZu10AJfvTDmTWRBeCZ0sg
+JFbo9t4KwD0a6OTI9hRF3yzF2T2WSHXmN8tvWHLIpJDDHIKFFel5b8QUNC36y+F
CykkCeGHZm8z3Symyfi6pt6T5iD8VNRoTaMwvaTMIr9pC90LCO7QS9x6SachEW9K
83gHIYvUQHuN6kkP6loVIGTvvbAwZcsHLN8ImOtjjn8+6D1VJbqPe+Km+PZtLC11
rLMdWMNqRqAZjzcK6dU+X6XAQwjPBfpGDIsDZZgHYShGfLgsQyd7Oq6SNgFZru7/
R2i3irJbAF58Um2VtimG3XuaOunG5rZHHDSmV3edkk92HAEgJNUtfL4f4XPci+Yl
M9JW4HjTXUkx8/El3KjaDr6kOsmbkgCLzhWYbbMjLueOsw7ifFwJpaDO/lDTIzO7
VuL1o8BIIWJBrQS4wr0ryO17aATvFXOauiY2GCgXBcnUm4QX39rAYZD2LqnnKaS4
nU6yhE8wJI1D8pxet9+wxMakEAYvJYE5Yh+N0vY6+Mq46ujh7mh6WKiec7vRInKw
JjGe59cTDNk29rRIdkVWoahczVgSiELKAQWih9kzC5y+x2WZ1rf7SzeXKU8avtCk
YKaakCdpJOgtqLLEjSXiHAEv9dz+WW+EdcX7Cg0xxGCdX7zaSWlTm1+3GNQb0Vhy
SS/lUxaC2lKCxTaIixh2U9Z1zaFs0EWQl+JZiBCLmFsnova0MXbCV5Wb0UJ8hpHO
kt7K3Dt9EXvVz+pOhcez7xVChtsqnMF5IAAEoGbsr4e1UvRAa62V7B0c6JC8LL4j
Z9dthhZf8bylzxlhxqof2COnQR3C/rFX73v/fItEzWWKdKg3lfIFF8W9LywlaaDl
WkwbD+Ihpw7MMWSr+pM1EFRsOjzjDGYGyJTVJ2gK+BnBD6Cg8GL1WEuuX4C/bsWg
/8uhWNRTTDsxT/SEi4drMF/FqD1N/uk05BIEvQaDMlYwsh5cli3inyXayFtRE/md
9CJIHOJuL70jPtkHHl+6fDo70JX3OMAuVCh35aBI1LpntpnB391wuGIo3EiaBu+q
0Gy7l/4GOSgiS7L8bTgqcLWc+HhjupC3JQRR3Bcp39cgUrgt4K6stIN99rmCdcHy
U3xM3H9xRPpMb6OCLmR69qC1GYdqL54uNWINYCg3H31A2FDC33mDP/8hBkrpJrOp
I+RHdhN8y5rK9Gjv/YvSSd93w+MDTHZAxeu0ePkygtC7p044wNdU2GXTT0QOhoUa
NvRFe4s4oYOvJnijznu/VCKlYxXKE/NK8C+YIvCCRnfCUcPPyz0qJCI78R79ZLF2
vDWary96fPDGzqY+GeD30L39y6TBvBh7GSO/louvRShmq2j989Y21fBgy9bc1ogn
nR7dRaUeDVCqpipyKckEZPHwpq61v7WiNJlY+KE3AltD0N9l+hBTDOYaaOaBUjrz
j46zILTXOLbgp/PbFgoKEa0Phojbzw6vPObbvH686FXKmY81WCDMvfcZZ1jKmWBJ
72Po3G3IlLBwhVT2GLAUMnUJBlrp+YjUxcM+3fuPNAyI1hmY8RuXd/iZiqt6EJkj
FzpnoP/qPkryNyLnLDeQomTSPNgdMnLKkSljnlEv3y27PfA1BD23JcMDeCrNlBUm
2Huq4x/fUmDMBppXCbIb05pH5kd8esdiaU+6I4rQyc4O6e+nCQoqv7WRUaDYO7LX
m+/ZpYINP4TkNvFIsny2zdHPmq9XmlFDWCrQfwW/d+MEwGi6M0Ov2JXrnEMniLon
oN4bFSNPs7ljEH6rKxIuNvNrqoRvuqJdlJ/iT+bZMgNwTP7W9HfzyKMgCRHz0OOM
lRAW3nImzyFDnGywd7hnZ54cFQagRJLrxRkc9LZj5Jk5aizj5XPR6S5FVevbxO32
89FLBzyOu3haJiKImrLwyfhjRv4mBjfq83F6aupbDjcZKN2I1HDoA/diPE1KRUnr
n7mxKmn4K217QgguOMKvm3nZXK/A/d6/PR6LZYBwnMU2VMOABkaNHNRonfzLalhl
hlny8g3YXFeKh5Jxm+1AvhjHhXjX3rSBBzCtm+1OucUIbaaGx4jXnQZ2s1sp/QZl
4anR+4rlObqIi4Ox26A7cNBJH9AIHJPUyKfoT8hlFZuQRzsGixvilvVoJbJaDQ6Z
fLCaaL1HfIkGH8JAeTTdhICpYD1BEKYHtWzwJoePtPJ196oND4ZiJ+SRnrVxatoG
q2V/vXEP1K6k51vUdqa6qnyWHdfxOG1SM4GEakN49+aXcoHWC3Yo6WbgpCxay1Fy
iqoJMwUQXyhMLo3+yRmZZoqEOOSBqCJYKlga5L62i+kicG8Gf9+CGbDxmmcGgX0s
4jgMX7ia+mGpNWXS+a5FiRi1DUznI3fUKaRz+1t8kq2ZLpC7pELOVyyQzFFRiaZ+
EP6+pGcGOuydfY9r9EhbNhCvGhe+c3Zr2nG3T2N3ooQDGq60DGkKvOHH/BbGihkn
Fv9gZCa2lAqT1uyCw6Wjj1DFljXv9IyScWmmtaNXsdK4Oz7bfs7SJweAdpBY15jc
p/gDwdN1ex2uvUKKvl3DH0S+9js6eXFKBfPCfRCWUPyj2RjWfcPRL5p1yjvQorCd
u76rGpKJ6fy54E51JliptR3dbhGI6E2FWyaLwu0RXNTgH8iC/3SjJh8Nghn6MNTt
CSOxFbfB2qvl53/iN5Mwuv0hMgRpwXRafaPq+ETS+kkN/87GaUKCS3xOzBHZWfmb
AyfLcnn1FjZYOiL6a7jW4En2FrAihY1ud9aLWObqs9SVkgXmuVZ/SR80mQqYSutQ
WRjJGD6SpfYqFu/zumW6GkRs16m62cxJ14qzznlHGnnrFU5cbUqvU+yXA2YAmURl
LnikZRYAmpSQdqIDJ/ght5kaoLE7TmbUDvwOc1EER+W0u7s1hSNvRZVGGo+ojf/j
fEXjfNRQMxbFWTxO/x/0HFCYs0uj9bs9evOAb680QcchmLTFmgqNn3imOnZgdRzd
FxU9x4DlF6nPwkEgw5PKnpGp7uJqE6ksEZ/reNFI323wMLGn12Hy/JDWuigS7UgD
NutiVrUiMj0A3/YBjbVWn1KI3JBamT8/3JLXSr0zt4lehkJkhJMvLObjWNbGbSZX
pAr6/IvQcKU99+2QoqprsZZwfdwnA/SBFMJ4Y6mYa68gBM9Sd9rmvP9aE+IqGeLh
ZVSaDDlShMgSM2iGMLPngSQqpqTHNXsrl0ecrri+dHZiiqH5RDg4kneyAKuniT5F
lQonaZ+rmY3kMPjdR8SG+ba2E6v4Wj2oNNo4g1HyiprOHTWFZeSY+5CjWnrJqJ3j
12eF/+/FWFAAx2voIgPYzrekElu2Zv/tn7YysDGAPMQTQltT5tXfEi6mAPF/RG05
QYg8OCC8QlBJpdim/P/nlNUKZCTVOjqRaMoCEileSySSLMViZoIPIO90BKX3shEk
kwjJayJRuVg/7F2weMGvb5CDLHfaWp+QKXv3qdUm6Py9ZO+uOFjrDlA42Ak29bLk
AYMSYpWG0hbMJIzffS8gBgGUzQ1Yqku6aitkS2n7AuoAG3BNAuCu0vPux/zjw89v
QzQPZB7QKmFPLbKYwiMXJgH7dESrdhwqomAk8pP2hQ6G4DG++SnBSbsXGvKdivNB
TB5KA9asIway9eqxZIqYVXC+GCrpsd11KFU5mxXtdL3bCPspQAfbY/z3CVRIYXz6
sZHnlR3tSsfRAZDgDi72p5gS3uEN/GClnnK5su6CeKvVcGae+fqnr6J9G6HuW5gk
E7AGHb4G9vd1YaBvIdl+WBHtTA1LT3GhkawBGZmw4BNeW3b9vvEXV8xZaHrcLU72
Bcf1prlzgzV3PEq8LAqeIbEMvl7nnGSI0ldRoB5xSe9uBR6ixm5IyUwfAp4HWUWq
YqUsG+KE5mOuOqx2LRjMcg4UcYhuTFXaSxo7WkMZKjHb4I6ZBdIMb4RUk1/fD7ww
724tRQ8QIcMHR1p0cyz8RslENywJw9mRpY1/x8BIw+vu/3No4NbZlZg6vXot4Qnq
j4WUTSHTegJjFWcKvRWaVMJtctWunMZz84zdET+Tn4NFSLozA/80VXBmShILD+Ji
63H5tSnHHynynp0sS2UiD9spnh7JNyfvy4NBZCtpRGReulLPKPuFk0UJVfsEw2Y4
n8+P5S+WQa8yfFkcbm2u3zbSy6JXLmPy/QVmZkq6xrr/M7tuGkPqvO5NNHCxVtbk
Nj7r36rVpaySpIKgCdugkXzTSIn6HKOGnUvaWV1xOV/ObnCvi0DaTBeOoWhQsd69
PSgOHBS11Enru7T/H8mNBRWdLoJWzDMes8uwU8d8LDe/lvUpqyP5Zk0QohoYYxDH
PVaduRqjYZ7sP5wpqmuSs9EVgLMFjdrpUvqCGvid7Wln4TZyz89XRvw4OSPCYBmP
wohZrccahJRcXlD7r2fPIqRNbk5uY7ipHpmR3liGw+Xhw8DarT73P/x4yo6S6Q/2
9/MRf68YRn9byy1ud0RqIOFFbpsVPSKSSjVACtqaiFYdVquXosNmJtr5u5gbwV2Q
JhHZ15iaXMEZUEmRcg2c7bGRL30u/68jFVdH9FALHAanWqmPAMrgM9sdRObbOEO/
j76Q7N28pzlIUN1nNH44Lt+Cv//h5tvBWNItaNFfSET9a5M9s1I+Je1Hjk9I5gy/
mXAqrXY+VmoRjv0oqt8Qfkxv9i9LeYtTpGZKqLAHXt3OACEnQ4zV4az/7Vv1+92Y
tkGA+Gmx+xkkocC1l0Xg6WioIzxRONxjoOMtH3GtVSVhmiuHu8dULUfyWU6eauej
3PAqEXg9eYEwoHPwBT6QMm+on+3wNFC27+uHLMEJmMov9ZETYcYDKkALL71WA/jQ
xO8I+twAASLnbuBUo5HDTHd5yRXp9kA8ivKVvOmE5VKld/oNtvAcPTJ/iEtMgqLg
EVxqfltyoCuN0htFqCUnatqOlsdSlWfsNpE15k75jGFJycJ6KlryOlVR/6BLqK13
gB1UQtvDR7N2LTucn3iujSZjZXhrJlJ0MiNuml/GaZmBW5DsWpuZKao3xYdOE7jX
/4DruY57YUajB6y7etn5w9wjZu5+UpEIMqyHTqGZ/dPb/Xxr5+DSYJZNj9+B6YCk
lnFdJnyVPQEoZG8w83OMDk2o1N0wTKHrlpQvQ5BSSlsTf+FOml4wg6Zfr6xtQreT
Q1OiOtUZQuEwwrPxKk3q+W/wlMroXSHunoUv1MOmuNJN4TsIOrv7LQfvcnqD7uzK
0mQqNfqRqlq8la2fPlxyf+6iltOfPMqBR6h6CYRob3FjE+E3Z6VYfmzA8yluTsDh
kBBmBMHSNTfrSRZh3pu91NRMy0/vYbmPSFA1SnyvWFeFRr0ivL+cRaIhjIMU+Ae4
FDv6Q2EqytMhKIJfXhcFd3V76qeIL9MxC7C4J+CUw/xcUC0Mj6gt6UAY+p3zM/Dg
NgV7tg1Jf8owl0X2NXheHdroF3X4VwLxHQmPVS7qFuXz3zdjW+dcXr8bJBcq/auU
KAqty/ocZoSCRs7818RvVG5NHfXos3RcCV4iFX1RKmf5yeLax13wyJjDntHCgY6d
XYQWL5gPqNVt/QMJ79N7DVG5bziXeeI+3lvihkBZ7UuLJzQ25q7n35ilUo7OlLti
zf4YuSTc/DHbnT4q92Z3HxP6wZkFETDwy4osp3+MvjrvsKDvxWqDmrmC1dTGvUNH
0mMrKE6MbqWgnprzLNMSfveTSFT9CzJGZH4BQyrhl/6zp+teb1vopwR9tSnpyZS/
39+5nELLUQPvjWJtSO/ZCIDQ4Uwk2v8SXceQmZ9PsdDPQg2ds3iORWWzPEAPmONI
coYyI1KBAyEdusIvyhkdo2qFj/fTEgymKAXdZRBre2BG/AhNB+ci58rAUHPbNQhs
vTOvovRq1I3TIcNQcLY1ksHnSguwvXeQhKJ3+7c5afpsGHHxHMuVOkmoMaVDe3a+
g+Vg1qzeY7aSmZVBcHWm/LBmLdP1MZG4ElKEFiPe8nR3nx2xmL6z1OD4uHB37yRr
PZsBp8yOA61Rb5wlysO1KvcXsAgnx89pywmpJUrGWd6HVpAETJGKnPBMN6nEiGY0
mUnClJwz7VMC1iErX86HQHsgJ5ec9FpLIVyUHMOADkUno/yv6oa4V6Q4VCGvIqva
CQ3LNEaKAjelHDM4eN56wlCkq7PWa/+DBlSXYSeRfWuezWxog8J+IyBC43dUcKat
pqlmHNCC21TmjJFXRg/ybgbOMDI/LInFrsJmrgBG/oJCjY9RwPYl5rYSN31E/s54
pnu/yYEaHwO3I/YmhAVcNm5iHhfhmsHNd92vTEQnMYRSkPLAq1vcI9TFCma1ygsQ
ZOLe0CqE7tKI060DmlSs8gaExPFW7ty/ZqS8RMsX9F1/3AGEFcb6LCfJioMBYq4l
e1RKfFr/eegGvMEYdrMDH7WQNqa4eSrBdWl/NWYTxEYIzoWbl2Hvv9rVGqZnObeh
aGC+gb/zHAHf1BriLtcCWDchfsQmykXXrmEzSypmF5w/xcx8lUxAFqhkCWkvfbtl
3X8vyTK80/08cwnB9y/kqxGnpfEoz3kNPk7tt8woPcwSgSZB43sqAXWWirtQ1lD3
+5mQaHgTljVxoJCOHBOCoLeWg/GC4TDUe8KXom6NaPaWdRNhtrTJ31kKfJT1cmXU
gK1SfEUOy9q/ERly2/ffNNzRSFwiBEHobIXe3nJUoONzsJWc2aFlXFEdZcG93RIr
a0My1TPqSni65X36sQdOFObdevTqoiEmnp24DDi30ncPZY3NhnxxFF5+/JdctW+u
pToPp62mEVow0JBMoPLSWCem9RESI1LkFIbFYPBLGzzvBIy+zAoLhpPYT73FTsl5
2BUvKoH/IFiRztppB9QWSt4VTkKhJqwB5Tc4lUUFCo39d0O0Ixbl2v8rjrxkdKa7
3eJzKFI/2CfOSfkQKSNZh4IT64QH1kKggPep4tRGcQydCdsbv57p1Zb84seN6ZEP
acNhA/2l3b1c80g8HHhce4anMU8wVnYxrXnlV6N0sInnEni8Vt/cuKSGHO9mP1My
GBvfcyQ7NoAcXwWHFNUoUHBcy10xsYh7D2/p6nlWujQW4O+CgfJcLocKDhz8sQtg
nhW99r0qNtYDJ+JC2A8tXNULTB7ivEXSMyroTsRLnM5oyxeDq5u+vwiB0MCUbRi5
LPdI5wTi8I/rrQ1GtedG61d70uzbTNWeZMy6E1uz+mOBe82o7l+daaNzXkmMRCtf
w3i+Aqpb77wY7qGR9nZFaYeVkP5Njr4Xa+HRmTG8yJ3WW9s/TSJCUlEedOCENWJL
KXAPsMHGbkJ7F24iqE8xkdWxI//MjagUU9minVMtEOOpi5v4TajX4+qjXdzUD6Lv
vFivilldO9lKxMKT79OeCZobHeEcROZmKkbOQa9GPYqQ3HGX+uBIAYVvk6VQrS0/
K14oBydgH+D+mGSZGk5eAY9dy64BF0h6kGESnaVVGSvZ498ppu5qvfCLyl6A3e/d
s9E5BUGakgddHsUcga53zTvh7Ag8HAM3In6BNfJSuDJyYJsXOf+qVENvas9oEP+t
h8dqvhZDojSk7JgC4M3pWf1y7+pa2aWFy1U39oFYY3tyEiHT2RZKgSGwEpaRm+ri
VNZZwspsSD7S3eqrvVN9t67VcSiGN5/4E83K9QlSHEdEKsAtkQXo4FESrN9J9CsI
JJMx/IUqPzP8CDArarVJhsrtPp3jcA9Y4azD8gf4uIw8YebOGyhmE7cmyU213m8B
IAH6qsfy6vNoTTMTVPDBTN0rzVKxFjY1xJhMbk/V2JeXJkRVrNNkoBSRRvnO4qMa
k/8xNDlESgwT2bIKpXY/2u1s1vnQm87dk6Nikm4ekqco7HfB0ipsbueU8+vjANd1
RzE/cyIt0XlP/gGNClhWGLiyih0sGEbyDLkcQmd4xnYZdm26gnFBIecmUX4nkm40
hJFriq6udE3qjOK+BkKKvgML9eiNnVEC4LwWaWxEIW0Y8yIsD/wXSTam7l/Ci8Nr
DGY1OZ20Ue3rf9MgPY68UTZgWTJWnMjyHFcDnJGKEBQvVAk9/2xtEzdsmfMeyf19
MJvUmjSddo8kCduM8/Ixsq18QgwZlEHERgaJ/cCtMomGDgJLmfjLyjPMBs8tQvMQ
JgSLlbO1MwzpJByaQ7E/DfaRpOexoWMvb4f1tOdAJzcmbGR6eeLYvYWbC3ueUyVD
mO4aA6Utf1/RlQPe6GCc6Nr1nL32QrbkqhAoRxKahwsRb4xGpb50GfVavSup89H3
ewZZThnLeC2VyGpGf4Gxcl73IuQumy2L8gm4z1HwbYC8psH3LfCeJvqgRC3DiVLX
+IA3D6iU/BhNDLFtv52kinOhC7W3zHa6ogpZk7+2nrMyHb5hg/x2qnyI6t3AO3U6
n2Nua+KJz6JMKmJEjbZ8vJGgUr907TlfQz7rlVwKf14JjEotnnwzACm2fWa9P5YJ
t2KGUFfac7N6b3uqOti4+BgZz540NjHrXQViindgsGbfktjOk+BOiKqEsEcpPOIg
IAmJBULns0UsPc9gsXQ5tLIKaXfq6TPwbU8Vi13suUI6b10TA7oJ09ddqE5Nc6+u
06L4xCzIxrVffgOJrQyokEmoHsct0m6FSj0hi2BcIiAvwhxxtgk+7PhfFIeeE5cG
8twBkZdYnh/0S8gznQ/xQCKH2bzViAkcytXMXNslCuGLt6LJ7zcXTLtnoufYj90v
u86Nc+e0iWAvJ9I6JDFR59S/EjxmB2jahZH2Lg5LUra40RSbfCrodDmmE/r4IpxH
+Z2qJhgkSiuZ6MNbkBo/J+c7dePXR+v/uIGM61cQCozQ1kVvWNfFvRGMbC854SWz
yOOnovMwSZ1w2Dr+MuIJUYGE9OQ2x1r+uubU/GykcqDNPTQwY5axaZNZHtEUzTYm
e6hOw3a7cdHel5cNybJCYdFW8OveYDkM7i1oc40v2a7ZgLIdWUPaAUJ2yQhleWoK
Uhaji9rD44d/90SldHUzvENtuc4MhEpXBfCDs5DEfvZOSO8eM9uUPCKy6W8R1gbM
rVFuti6Rv8d+yBo0StWnqRxrr/vos4JxKm5wYez8RsdZyKr0XqqzrNKvUJtX2xWK
TBgPuqNqz6M/HVnM3YQoXuRHg2ElE+HlHJMsyZxzsBGVpCY1lnw/VbkRd210gEWx
kkJFw5ZfEhMyiabWr0B1/SCYHMueO3k30u0+fO6M6oyLyje/XjmvxUqd5gxCGRnF
AWZl5JcrBoKVn872M6uEbsk1O+DNPVC3r+eV9Fwf0D8pbUHugf3xZORYUu64K11t
QyznxxAznQKDGMNwfdsVqlhug2S1FieN1U440DPj5itfyCYHGAbAMgoRDRmGRL5q
YUCl0TonV14izRhwyfd95naoYsb8ryulPGGZYNjsVDHv3nfbn991tacGV1seW/QB
nafFTsg0zIzttJA20ZBqyk2fJKLVMeLaeMuJ5QW8WBu+20Oy87UKRrL3yd/6H5+h
atJAZuZ3E68+b+c9a71YTs5rphywtWtbVgl3tKAoQ+BDBBUg6MXbNzfoKWAoRPn/
V/SCb4a4M3lbIqvnG4CcSnlGF2ZlLplMJFD+LzaErQdnL5xdwYNg+GuG2GUBWUr0
P1DrIdl/iPjVxaLbQARyYHpN/ONNIPmsI2q0xsaUKnbxw6+mh3FmIcS6nqi3HvL6
b90Cdzt5p09C5DuzLixukrTUQVyTH9EAjbDdRZZ0qheIWhSHtaAz0KV5ybDJCNaN
83mEwh8ix3FzcvyizgstMB/lBZZEF0wlCQjoBiKm8AEW0OxloajcRmvvmji+HDOU
hUYuHsvf4h1G1DO0WavDoSoYlk2bmV2yW4zlUgL3+1OT9jMU+JC0rPx4SIiYDbC1
+dxlfYGGiZXcqZPHdkwbMa6+GoCJbJUmU9S1W0kvSmSV27eNMTN3oPieUJZaDiuD
KjarlawWnUR2lkn42UHcfNTM3EOsfpE8kzF1HBOyHjXRakpZwSDVnxmFDVBuZus0
x1U0kU/jA731Hk4JOLOzdkS8XktNNtSETjwGFIA3jOCW5Pi9JR+Nu1uBb/YhB7J3
eVNrzjLgEq9FxcHvteFGcywWtdAecUUx8punE2Oc7/bOp8I95EUOmsQosUwwXi6B
+gDfeqMLDBDfBdga4OksR2cl/rFpwaUa002HMeM2mHicDZpnm1wcB0R44wePTASn
OMBd16xNSUhQxdNv2N0/ODN93+rY1M5k38HUlUfpXYhwT2qukt9aq+BKeDCwdG55
Vr2DCb/unJ6NAu3iHhn2EcAWYEPYpgb2szKv/8tKkwFNRVxinJVLA2D5HF5yzsli
2MsGiSaKbbycX9xzo0zjBZzyvZTEAJ863pfKeBxC+YdWmdIDhbg1aWjfCOU5pAGC
GNIsZl2ixLVGL0vSzUaWJzX0Ua4oAkJIOGE/uVJUNpqi9bVlbPOfgfcXkj3+xLvM
GOP2FN60Pi98qRHHu9JILDCqwBX8MfI/KGWyMLbUipqFx/tL0NXQMaDVw2Sex0Og
kb0zsjfQ9/fFyLcMbz6Lo/lYjrAGNxppvJ8joIM6Mx35LdGijTh7wSna3v1/V7Re
+DUATdypLAlb1yanWko5ZBbPMsU4wxcucivmdLaPyVhCFWK8eTqOO42W90A2L5ql
0Xwif/D0oIuatvKAqXfzhoQ61EhpGrA34NqIB1SN7mWHZwCXGwAsoABi04WBXYcW
X8ywAOkQ1UzHO+R8ZQFB7WaGWUnqp6UP6nEruEgc42CDCEGAXHTNxzjF6kaAvFr3
kMN2/7Mj6+kilRCRfsRCjNiz7sEQgxUxKgiGX8sw1IIi6dy5Lb2woSCQknRIJGcD
mqOuguyk/ww0pLPSJYFEkGiW3ZqzyGwV/WDCeCBvTDZiqAa7otAzXFbTwjNytkIF
a79lg1dd/cYOmZlGSJ9rTu5WlYQAu5O1uJabum4lp5g/oRGfLCHj4pBpjuWccRl1
ivqPdbblUF7Y1wGm115vO6BGsuKVvIBTPJSQKQhLg7Gr/poCRuUJUJrkb/hXMIgh
+U6+dYWDfZ/FCwXvQysTOC3e/H9cjc7s611ohBwhP0rf7BvO2i1aPerCIRuDUXMS
11AoZBTar3cnzfsrSeh/gwX+9ENWUVKcHstelYp868ebYTULoCrcOiWRMdu3Bvn4
G6FflMQvUlGaPbR9+tEvbmLLamiKojrc2YCYeA4eFLgFH0brhKoo5jOOHKJCKp9T
nQ1DUVDmKOn9YKQG098XNbkdUNAkPb9cJmHkX2wMvxEUM/Onf5zZKDyvViV9F2ut
9IPzw15uo1snlggdtMGv0QcdLfToSPqVWTCDM3ZpmXMpW6elmQ9/oIiX1zByFEvj
4LRJKu3DmPbN7VtrtDsVN5uDY4bLi+objgkiJOUe52y2uJ9zJmxXSTfhh5xRAzMx
9XKx8w4DlPMmw7IZogL7rzO4Szl0JXJUrP48vRRHpdK9I/pieBWXyCMF9mBUU3cS
jHe31rXloiofdXAuzEfjYWGVbWEh9dEWelhdaiGv8q5OOQxs5mvEX5YbeRqjyytq
wUtPFk/sBpjIt6tBDqmu+Qp++kwBWV5muY0iif46Api4fEVl0w8XyfqfCQUxve2p
pHQdQgs6JsrJjxxmiUkd0DLdiLyfVFvjISzMhYO9HI9zV/jC8FYpOJIv3sPLqjTV
oe+T8sWuD9h7NFiqtDXttCl9y+5rsdeLjGwP8U+Pjo8KOTefS7f2m6ZtWfwQqWNN
Stay7HQVlgdEQbS4nQngx1lRd6Wab4Gm0Y/FmAzkU+pd6QYeBILgXtBuEng9r0sM
C0AtsFWjcSigZYNK9ctFloYx8jVY0n+SKmsmxAHo4Vz+b1tTnVfVO2eBX/QniNy5
LQyky6kLFhpIUS+UMMjvjqWSJc7aI3hJArzCe8G0N50k0S21DJTgNIrmWBJlP08N
1vyQGzeM1sS+HudQvGVp7SiNtxyAkJwPpn6TZR2dP27rZBigIMDYyGCigOM8xKOV
jz1yFRHkHfD81TWvq8GwAJJWLOTdI1KVup2+hYiRKKx2TaDGXobqnDbmqX9YOC2e
jA8QNVIgx8ekomxewU0UQne1vqwbSCGa7wNsMvYCfQDOQb2q27Y2A1VJENhM1hau
8UdrE1x3c9/KaBN2A72AtTuvb3m2TdIbFFxir/f69h7Uu+RodC9GprMyJ8c03ZAN
1+mSBw5FHnhBKejcTKomj1C2hFsgt30MLLnk1ZqlkprNiTjobo25Svs5n66bVTuB
KHOvM3efTpK8vjLQOhmViqK1fSDSaKWEbesbZeIstzaeUdkv0x+nbFkWfd+x6AYA
ndc/GEsdQRguQTnAgZoHv+FQpsd7cHpIrW/UcnO+eGlO5XKaL2c7eyznO7vlKJ+O
mzCO+yqMNUzK2/zvSL349l3ljtAB/ebMi5bARsnIA6dUE18OeZYQUAkWAD40RVwh
vVViFRp6DP5NXf5l9CvpsnxsH0kkmb0EUkKXfNLXYeC7jlQHqTty+eWrGIyqaW7B
eWVJiU3+11SSCg3HZlvc5yF2pBni0RMYW+xk5bwYgApkkLKEniy3hkmAo3ZiGuFN
x4aze4smgkXSeDvxk9OzdcmpG8z/TkB1qtf14e/sc3SlwSMczrQaSvWqLYP0p22K
954F9ra8xY/hQfwaMsPvqvuecRVd1poZkzw9Hoz5kpeEA4nGO49x3OPHI0EtkR33
bAjuICxmZ0rO9V2zjtZxqaviVCxg5vHQMiU8zX56VNK7Qy6bF8Fi2Fg4EnaYY2QN
WRtNhNm7PaxCFgF/uPLNyok+pwS956DUw55qzoLdq6JADUH8npr30FM0XkIWbYLP
oCnQaaTCwexqVEw7s25p7iItVepMoYYQN3LT1OmpB25kkersaRPUxeMjq2ccOqL3
8JECW3TDWc5+DmKg5/gPDUIWVMrJjOK7nR5UXUm/6Or9sb8TCukBbAAwMhcGKZPU
5y6llChumQRB8aIjtwqKsugvzeYDuRwSMDGboS7UxQgh5oXsApeTXHMR+mKMq1Rq
y3bO0/oHhavo4LUAlbhYSa/AgGfvmp4OagVyKfP5ak5EGTcRKB1qgJHAKmIB0Wlw
ez7IowgjWApqCZQPLi8GVXOSwm3f5mHGUq9NNcV0g1SC3+Tqt3W/D8TYxXj9ZPKJ
w+KSTA4em79AAU1fOyY1BDabrNSLYGEzXXQmd0dBmYGbpVE3ahFxvFwABrShHeAP
T00IfYSaw6Y395ivx4BpOPJKWNfRkNGzJMg7Uonk7trMFnx2jMXV1JFysCxa9F6e
kEiPqWtFxHiTt89UnN9TVgGBJYJCBtWWYA2TMUScARkiuzZQZNcXyrQ2mahqCaKT
a/X3xswsFuwPghfuLNGFlL/vFaS4bY6zQU1wgEcK18VVrlPFSAYDpYAxB/iVaabv
V+sM0XSCBx2KD8RJYawRpXfV0g/adTITm3W1IIuuEfk9BhsNBtbpqaAsN06yLgh7
dOdg1/Mc1Ezonx3RAWZZdtTwv+E5qnFdimdCPtH4mqanyZS9wmMpj7CnAk45o9E2
N/vcvqXsIfTY4Zq8kIT3vLkfCN6NfSCmpjotTXsoZdRxulxGqIjhvwaIbdKbeG5F
7B8D0va/Zbx1tkub0BOuaOmYP2uLQ7Jn62ZqN/0FerjmiAQlDr2It6HRmy1bz/HB
IjKXX+YpLudkuOpo95TmCOUXDZq/F/7kOD6csrCwwzqV5XA5i6OSRPXjrBcRsuVb
FSXIq93uNJP3Z8TMCD+g6+hXyQypAKcX0X6BLnEkQXei7bEDhS0zd2/fCmxn2wks
1zzh8Ow00sARLFuLmdEaJdjB6UKwHjVWj9yQ38n4LYXZyT+cVnVTMcMZ23ge9ncS
RQ3d15myX9osVR9nXyzm8QYj0ZRDfqc6BP8Uc0tk0s9OgNaoxuVNf/lvAT6aSKyI
16HdxFznC3zfMSWXjvXR8kc8f9YQWA5TeX1ZVSoXy8ulKEYwZybFsDUbz0LyYz6g
0c85g0/d+X8dCkJkqcSQ/44oJOU04uQnEBXMDLPXGeGlQEP/xPVYGv/j6XfFF9lE
h+Te4cLL7hpE9+5estwNFBDamRaCyvvVA4GzrOGuXLJo4FdzsuRO1txubqYMh6NE
IgwzXh/s8sM2zvi3iXdJnx2ESVtsppzqQviztMsfCs6BlOFGz+yCJnIXlpj0qWFJ
Mv7jDDCZRqFhQJyvt/2CCbj5CTvvdI99ICGfjQGOeIkOnniRZKOVAt+0KF7TWRQj
VfLQR8HNddngNIfaV4Zwx0Q8gfV5TgkFOIzUxoxeqPl4C5Dg5rWiqoySwm9eRlaa
cW4jk9tyexXnuteHPaW+sx3KlXibbvK2LL81GUxBFBdg7I/ceeKQ+0y5wJbdN/Ga
IvQc0yHacTeHtZ7WoBgl8N1aQJOeUJCNh5PDcnrVHMICO7UClZDpPwQbp1hDEtOS
jz1AvK77bn/GigTnZAZXnVc8Zwk4C2XkI/sh2vv/DEPWQiAIX7kyhZsEq+UMmDGc
MLpj1Flnllo7rD9FSScRiXRH3yTcXV4feqEtLoGEJ7QePI96O+WUTcGu7MKrNGvD
eLrD2qD55ZiGjU8mfPdfYJJ/EJU16iHLngeAg5YZ8z4EVFm8e//7VhNF+bacmbVo
XqOIJ1BjkJRT8K8z5RG0fnXzpkQ28bzHaOGLADzNNYgfTq47XL8j7eXrNTH8YwxG
yk23G3J6vMQrmqxsNgwmgjKJjIW5o7cxu+ih2fOYa9oafewYhBAxzBSBLnLCMu9D
+L/kSNDXHFf6karHiKJmtcOD+NyVEGWW4O+2TsQ12M/9Zd/W0zCHwpGHd2r4Ay+l
wcfPt1ZdgBHhDs3nBAmdTTEmYxALY1+EfC5cKWDjWIQlk6/QXjrr3iM8Z+awrp/c
v+MdHum6GMpffwXA0uQ6w9wGhFNfzN6SRoTWKF0YyyzaE7CpWTQa5MDJlTuN9xLu
pvmukb8xdoYMevw5NgqmOpunwBCBw9AI0ArGJ6iAXSjmqCJ4nQg2jxm2RAz0uTQp
y6Cv5CMgMuVKmNJRGRb8kxD6OWFXitAY5BKTwjZBxIQimNJJwjZwwciSY4V1jN9d
Wg9gCHxxUrqmSNMo0BhvZPLMZ5HoJhhl/3ZE7Ad9f4bF9GXbJ8G2p3bqWTMIXUpE
s03LDzhJBZECjzRMGqQkxoMQaKfqhfHHVoffWRxoKR3o6f/aVYdgyqyiNrcIHOpQ
8hp+Ys4FbfHHZJf+ROUi+q+v+MnUEOIs77DW8cNMiLE8CPV2aKsCZ8ecDJCesMko
ng6UfRE1jCYYU/Jgj2ce8eCNup/VBx8gYpJfhvfKGiEYnGh7hCcIrsNaaJTFQMMp
ESQe4a6Q8SVIFZQ+UjJaUS0rzAqwa6acBdQi8FKmlyaVxlz4KCk5LTxc7Buv7+pd
tWurkbvTEdHrILtj1Cd7AumIZ/iVuPLQ43H3oaMwY5FtGvKK4BoLQkQ2dKcq7ptU
/pUsE5hPWtSCZ0PjIjA7b4I3q7687dpvv9dtHokiqUlL41Ewr1qOn0zt7LK3zx4N
dK6p6j7BqqiKtn5iUkakeczNPZlv6lKSlCNYlIdihIWteg075QAz9hlS767qfP2B
xjvRQw+4u3evskksdi9oAnqx6oF9/zxvmpDJz3xUNsep7hXPJ8pMcLZx22dODQcC
rEUoQWVzP3V/GTZ1EEIT1tFtxr+a+NOYC79r2Sz76PrG+XU7BDuOazkpcF7EcjMz
OVmhsLTnqCrDdOjUoGdZLui5Yu6hasKprBsFycVsEWdytA8Jz+LhURm3p+QvgBCu
sbl8O5ddOSKcrB/5n/gNLIibNs7bq7w8PnACRE60FWYL0X3eAH3hKjWabZB5FuXJ
T3uT4SaJ7lnSW2ofhHlYmx7NWaVWK8ajrSkwVPV/idAYcmklTxr0HqUIpWrFGjE9
rIhxiTDmn6dnE1ZQDNIpEi+RKyuJYiSe1jm6+jEcUtatSANyx0pv4ayZJxmTA5kO
NfoyBKIzaNPuF7jmRT9m9/50TX7Zufo7crhnFAyxV6L3ivcNseLGk1ugT5egF/TW
gW2OoWRavfTw7Y2dOoNp9TYdZxvApiqCj3CDwvZEtil+l3zfaBQVKti5pJGwIiFL
5O6agBYefodYhYb3MczXKSAkXL9JJzkIWublU5Tt8RZ82ocHzYrQLaNqHW3m15oB
rBLca4g1C++sDFdwGG/Go8V90i1aIn4IZEkAfpXEPJFOO93v4cZiVAcFa/yYQkXa
F4XiREzUJookc3jRw3UI8FHEZ6HqO+OrOCAgA1xXpZ/tcO3fCP4DhFCDxkbOvyeq
WonXT5+nKjTTI2uDGUnpoXqapBjn7v0nTCgUeSHsin5l9nbbnprn0puK9QJv5oCt
6zC9kchIRmvNnFHfJTgjlcrVQsOn1nASRse7vaTZhfTBu+JaqU68zbv5aGoFf3wZ
Erj9KiCbJcFfXQxDnMFbigDauLrh7GRuPgnVoIZZ2lcPOjlXiJN0bUgeN4m9mu7h
+3gPbMXDsKPwXS7T9zB3UpCpicAdaBMvhjf48KNkmaBYzIM3BYjawFxZ57CdQtoY
nBZLXVKwM56R3WHaRUbwZfe+XyYoFX3pFSr90OnxNvlxwwUfj2TutbVVcdTSbbUf
v8VrEU0EtB26yit0XFqnm1OrRKAMMkBXTE9bnoi/K7F7dexe2bWAuqnEw6/OZnK1
MOvwMpWyc9zMhMHwGBO7PxFxHVK98okuxhqi+7H/boPFMyZ3stYxsQ//KcTPlkIP
NrVbpaIcH1fqw1dxZ33UzTqf4sXJo6jSLoNIu+2h2K3kgUGzd2s6GaUsTmZvZKSg
4FX4G6/ezy9NDyDHrtlfrRvzm6j+p6KUHeIlSl04wnZNu/8zuurO1vNDj4g+dPJj
ftW4ogpzkHye1hDJxqqK3BOFwcDLS2WImXL5B3JndsxxcDD30wbMs6NpPEBwxQst
1ljAuPMxBng+U3TfHSwn9H6ntoy1BxMrBPt0vQl1U0IK8GY5QBh0loCuh5MY+i3D
mU3XTH8/5Pckol85wIoT99Zja77bxQM3cOFQNpt3wdTX6ScC1bIgZXhzNz9+Poa8
99sXp1n8tqI921WQUlBK0n6WHZT05lmObF4Sm7te+3mci0BTs+0krwrTSgSsyavo
labt/P5l0qhBLtbfABj3P2V4ZBSE1E4iSJ1Kj686jgF3BJonL6+/Ydbc5nKHdzlg
nm/JuqcW4Ophx8X35kYihQkBfY1k+EDleVr3bpGxKDCa6KzcMqZdZpGixLsnI+b7
ocXZ5xRRrfcyHVVeCEfkUee9UB91E79ZN7H+1y+t+SoWrmEP5Bpy41UT1Cagin6q
aY/XLAMkYyi1WL9ZpwQzg+6GRZYcDA8VoWKlA1pPMN4KkNkelKJIhnZARpn88IMp
6s7+B0cqwcsRUqkm1yuSbltFUFpYQucno0jr+hzHuUieG355/YFGLxiyJLaLvqpE
Jlw88yUW5Z/E2qrk0/q4N2wSbKv8Q9EOP03awbql0BWhQFicxZn1FWaZrsu3z/YP
xaY17v6TQs60fQ7GxkHB9UUit84NEP/FGxF5Fmvc+QwFarbWOsYvIiZ1oDtvApoP
O74qgEvgDQuROHVrPUGKRUrAvhe9PahmtjINVDBAHn1OJ5Rarttt4wtfT9ROpULz
JRYEzb6u8r9StgrxuIcJPo3TBBJWxcBTeXluuYvJfhikRAq9cbG9HrDcb40ICUDy
S9D90r+AHjevXyLUslj1vQTeHzdAG7ajo7dtybtk9wqA6X8kgdEhOfbnbKyv42er
IwN37vh60rq7Tt1pM/2bC6D7Tm4Nc0wgeSIY4SHdXADNS+CN+eos71fR9cItV56C
xSQmFkzZ2E5Ef+plDtmFGtjGM/yp1anETI+a3pa44i+3p7cwn2SctoVVGwp+/aXO
++Gtuj4cSvR693sYvfVQCGQS8sEow+qj9952jbr8IRmSi0xZfDrPcz/XaAn/4tTE
07VERUWr72Xf90TubGi9ShVeoDL4ghw/rm1qeye7XJJhok0VFVjdPG4V9KXyPv0/
IDJjPy41UTfx5/F2bR0sFFF1c4Js76jZFIVoJKIgDQBdRC5s/DTioyCuURHzLZIL
6Reim5IssD54oe+Us81czS0fR8eBLrsp+g8Y9vnHDbO9/HAUg8NUvn00A02KUjHb
tGg5l19ZgIuP+adrCauDofyxZGbNZpuo/f+p8UgvJU3rpWC23BZOW3U5ow9I0VrD
L/o4WCLNuTGu3NLEN0W4kUK3prQ9AfyVNiDXUhIeSm7lhmcKCzCyeBvz4JHBLh4e
dsGmz1d7jhYVDe3Xw3NslpTFhq3twN8gSxz5xmQdNvtS0rIrIBl2BMquQK+PhU27
TImpyDtE59Tb2McHm6fVBNn2IJRt474eB/ugoQn0+O2LZYwnLjKtfuc1VvmSzbRs
6IqyCFreJx5HJzGUJcsVYsmK4z5gCIXimXMo5ek34F9tZhDhxaVsUynNkfltgHHr
5Ruc72reSgkFYgJ82iTAOdiQx9pCbMrV4p8ihZJXYKovYyMgm6sSwaaHJDi5aOFW
IMSxfv+4BMSAJlT7J3XFr0wzQmdM1J5c1oiiw12hxmGLOGl7+cgtjBb9SHxOqYIa
uEJrJdCvpX+AriO6HfkwqCsCyM8KZmnRZx9oAxn2HmbUIRdoNW6XbptXMTzU5fpU
HfAQSpd5GR3DxC0N6KD8hH8apAPYM/xCbWyV8yiUl8YbSgoDOBnPBy4icahII7/o
FtaF1mkrlWWPL5R0kjRdw7lCYul0Ob27h/ZdWXqvzV/CK619U4C4k7jVe48SYC39
dsgYmzOHUvSmSBWC4GltKadQZW99NJLGpWRiedj2t3RwN8zl4Cn2MimzRefoukpu
0ukzmxCyMeXQwkGzrC+Yc7qVJyDkXLfLJzmb8EpJD6invvWJnpn4YHFpZ0vRReBf
EzvAGjHs2RxIOqgU26+Dl5t5thKWsLDJitzmP2CtKXuq5qMzXXNEo+s45uMV6+vY
1jzM5whqo2TXxz9rhDGidGuVxF+U4iCN2y7mmlAafFKj2E2Z/+Ovubwb3tMzMsSx
S4aPENqEK7p7D8KW8LetmJ1PUuV0A+wEGPQT5qx5j9z4gW7EJddZrr5rMTR6X6xf
65rns+LxF/HcBFnl6SITqtpkg5OoF0BjHhUrUTIY6oiEuVH49FBFb8CrkbhkRdwT
P0aDJjAsAkLcoXOpxGk2PPiFYQwlGdYj2beP8N96ORogxmGZYpYuOhK22pU8AfAW
gpiz6vjOf8LwaB/+pPepWcCGwz4iZ+vZf8fa7Lj0yot4seXUGu8gQak/w3/uCKdT
orO+yf/I5m+o2i38n5fpWeKxtqJnsRBKt9xwloEwRafaix8W9dp3lWNO4ZGXkgu1
4qc/GW0FXWLdSZndjrcE98UXiuj7ma7B8BvS6neJyEfhTR9w0kxzPsQC3X7u4qFS
MT4dald0Xv9nXdX7DE2awcw9KLN2gcGZgAnUqlLD7azwHLgPPi5qWbE/g90m53KN
zr5Q14OcJS9nfQWbKeewk9f+UAOpHNc/XETurBlkGMP/vpMT3BDL723/pgEtbhDQ
kED11uTGLsLQzvLBgfsbQTmdAD+A0BfChjlkQwK9C6vyAbh7YHFR3wzl0H2wGcf8
vILTWVm/83P5hbDe0ZaLkJ1og4DmmJr4m1H2Ct80vHnbu+cbke2B4hpGHoN32Q8Z
vKU37roRkUk/r+h31YPSM36KTocKlYNv3Ce8GJuaRyXxJBnjHt9XnDVjeWgRUEVl
s5UWBsAVxhXW22hGlhcSWeegrjDFuHf9/gS0Dx4ehYJkeTGH4amVT5JNJSP3sO5g
Aw9/ofShGGhS+Ws3jA+XXRGwQ+DOoJ7eRdlAkKppUhyNaaDMUpOE3Rjrb69F3pR5
//OdQfrJceSjmpCxmJWl8hdGl8ZOxXrm8phCLfvpRY6QVeQr/O0l4ahDddYwEM8b
hL/kfyvBfmDcNnPPzHNuLDt1iarNHtMF4u9Dv+e4o2mMe2EYHDmzsGbXj2DhKAd7
D+C1B+OpYgZiNASekqudj/u3g1JpTRqyFblURAovQrBOHk2RIcz+d7ILbXy0VZbD
6MB7O0j2Wh6aKNdH2yCmydTtwz+T3PLE6MZmvkPKTuHCBQKi3JCtbS3qM0A4Ys8t
lNCX6eH2kf4EFj2ln4xfIOygyn+1jqHoOnDp0kXX7aXyGb+lzNB5ar8Zo1ZGlMM+
YDfdqEMLJ+5xDXmfnoDWg0n7ZcQDJszj7wj/KZk5yKPLWm0Q4YDUHaAs73TDoSS4
+9S5S2TTzdPv6v9Tz+9N+y6ydqDq4Hk4t58g5zNbcGFqAXVP4NynWUWQIJ7P0ccq
pJVyyzOIUa+owBDgl0Gk4omYQhKWA342q++Oc5ZSigTseIZCIVNZuo342cY/8Ois
1SSqgm/qWMUWzu1E32cRzEYHOcCnXUOmi65QWFMHFuSorqIzeTdbEXFxhlmxv4Qm
qU46eMEb+BWbHg5zV/xnZee3NTNd/dhnrjC4e4SnW3tqoC7YNKUHmTG6WDktwv+K
HxVEzrkXwipfQZv6w2p8EGezOgIt4n2PQG4cLM01ANg14CSqJ+3ZedTDFschseh4
fcfFwwKEmz69enKavYyS2YE5celWR1z4SbplMH6ccF2dNUg11ECa0Mt9RC5KrjTe
WJc2830G+9glJ3eTHjd/dq906nYqSYt7YT8tUdaI4yUBJYxgwTe3iIf4oEUuabln
Xhz0NtAsdkpfhi4HRAAwq3MBw9tMJOVNP/5SRFW7jDeBQOtsdqiKLtyYpPWZFaDy
7PsGVxAjAXazM4e158r2Z9l99OjNNI86KubH5V0gXov7OkVDRn0Zam7EJZox8MNs
CvygOP/7fRoJ27XlcRz8rprOrPHDLuwURJvUfmmEeqziDOxEjMt3ryuuJ2JGSS3T
A1mRTP09q1+8PSmt3yuAkcDHhq7jm2m689meFdb4YoB5yXuTU/45nElmSMxBxn70
1wmXi6hdm9/D5tdbUb05xHQS7uLMkZmqs2QrHayRguZSLCfsezK2XTOE5STf+66y
yGIS/0LOlFY/l407Ns5eWHrFNhyAogrLQZh1ray0wr+AMEUmlmHayVYezsre/B9c
NWO0RXnVAgOPZRbmZGZM0waFKAKntGpXViJn/Q1m5PVAfwo3sdcVMM4BgL/LxWUd
L1sOfakmdlhX9PP83QIoPHCRPTGwR0DZVfEFgqMpn0SRvJ+ATgfKExquw5dwIURh
VhrCZKlqNj1Y+pXzYLjr/E4Q9RXWi9Z6klBUd2BZSfn+5XquViICoNUx5RMZqcyH
MCyZWmWoikVux1T7dk6tmtrW06i5RIpYXDAKtG0BBHp27uXwJ7GHY9T5SdyspvvS
aHt50AENNAvG1qrltDBQsbiq4PrzhygPCfnZI2TJjaMfaatqrkypRU7Axfpnt9m9
+1rNO0uXAjxlrRorQFgl+tcBn6Zwm5c9NjPM37HHTHLv6Jivq/BJSTPQ58gH8hm6
VGbFNfRnbhf6CT3+olgcEDPdSwO5XPTC0R+nAVC79FknT5QmbqioulQcWqG7H865
QD31NQ0aAi6AF6mvHSku+KmlIAVS/SY3uK8TP1s99+OGAcZrgHWtU+YcRDnib13/
OeaZjxG/a1Q82HfZdJljkw8lM0ycjer+lEnQ22+7Z+EVFnQYTTQZ7UmrdVUMXaSd
3PAje6mGfBpZ99fv0pcmTheO1nzObuGFvWFUl65se2zVdBa7NqtiIflULfOPPkui
eCJqM8OT1UHQqDV3JXpTuAOaDaFOJvolIPEKDELmWiS5XIzpJE26PM+G2GBwljqh
k7AdqclAdhkbSTLLaVZvZ+eom40RwSBf3p7UIpXuU2qgiKBPTPyLZYZLiOHf2Ljk
CFqZqYo/ps5ysNIoXwHBh7lOsalmm6aa5wJCCFKDzA2E42zWl4oTMqtSWVEoDQOm
IxzlSpj8saR5QIhJ6GbRyNDQbjccBZeG48rmf4If8Pt1lGjFq5LfV6gPJBfbEWo+
ewlj+dAyQMuRro8NKlgSdUq7yvuDbzEMa84j2Gjg9cHlLVt8JQTSQIfzLc5k9blc
MQSKBga7Ve5flbpB88A/9n0x8GpznLh/S06Xpz4YpAu7mLRsbDjUKnIdV4pagszA
QG7tvQL/7escJ7sDBMb6uB5S5M0r99rb4q0dIaIMQdxdCcooxZm9ITYYmf74qdcH
VLQnNZRznSSWCr70ms3XYb5Jzs+W3jUoEpfib0WQWdFkOa3fz+UItGxe7YnsoB2X
IfHLpw3k0Byv0VAp56fiPrTO2gNCxT3/zXYrE5S6zlS4EBGQe6mWrVHnMCqmhTEG
Q9N/VNm2m4C8fRnwhopz1sjRrP2fjCRoCwf4fRkdsUQ6RkznsdECbiVq0kC9UFE6
OQLHILWA4ppf3vtsXWzO7lZqHoBU3cqCct5hnIW+/3TGF/WBH5Ahh+dLIMgPyfNo
3ijDemYvHsz5+x2En0bbddy7zYdWHB0ifLmaWg0Jl41tWyiVBBKmLSyhTQfQGz1M
8vFLlSN6GTLKqx/2MERZKDdR0Dm1o4tObK6Dyt9XmLlm2wPgbx4pPSF0eOn16IL+
xsoCD5eakYoX9/unkpDNqPpXuDbxFrKgYqhfRBqUtVTMlQtlEBisi70ixktC8XaB
0N/YOawTbERSz4sBjm7HcaaveyYNaplMe6LnmWUPO0cXSflztjJE0UObkGGhS5Fg
Zr3ulC17RliBiI0SLErw9SaO16lLAH0uF0X9tii5BRJnSavwk5MDOxSJ0M4HW6Pe
YMlqiRJYtu7Bp13aiI+Dp482/tQcw1iClKOq5fa4/kTPdsLkXnRmUTvMGQ4geaQ+
Uh/OD5ZDiLdl6l013MVviD/+2ee+82RuACmlXfb0MSquGj7IxhO8KdM5cKNmjjOX
L6dzMotryOmmY7fpctufYMWG1k3gQhqPwNO72/bBxgO1WFt5PnmPaCS9a59OYnxP
fncpbHKtHc4Q13gt61Zb5e20YHq8bIkFBGGF8mD6CnSO9gGZ7Gau9WMVwwYmdrYP
UxUynXNjc2Z6uKRLYClBtwGDgzwcI8Gw04EYeh3VTrS+pm1Fb1IHnhTwsnZth0TY
LxhOmP0Xp4r2OSlFDCP93kaNpqK6S5ppNuYm8BP7ll6skBeiqfi9DG7ayZ7dfFTo
/RRisdLfuBx4XG99YX938M71XkKhA5EuIYlBt6oXtRdxs31dup4wa/UNIuQGHy7d
naSpDXVn7XvBR18FvLyZhMiuvo1yMlCvnvncDOnAWi9341thBxBwyGNGlrh/vO8r
EqDkFKd0cIF6Fud1wPj2XMF1li9Hyh40UfXjgjlsJ2omiFjSAetENi//1pMoTq3A
OCPKDGEvk/Hlaw/64vxeaB/rAmZKtoApEiX93/e6Eq4FOKz58sbLPfOeZ5Bk0EmD
w6H0akSM0RUrYeh83yRgJcUeDKfKTqDq0I2H+ma2LnBGCzJUgT1vVuaCbSvEW/ZB
yDeAJYibFMdTbujbNEBaDZ5scSkKY6vudug3GyyC2B1Hm/UkME8bjvFYD4h8qwbf
MJ6QSR1vsBvAKohRzDWH/GRZ+wdUxbr4DSjfqRkmjo2kFsKfcokj1QwI6xWrxNh6
fcC2GXU4BFicWg+muikdZ0sURWL4Ke9gMRPEa+O23a+cGAljILZQNPTatLA0Cljh
95NM0yBUUs7DEX3UDP5/15YuBfVdUPtbKltRbNZM/YYsqjJ6etX4RVzUOONSCBKT
dCe1g5EfND8eUCbWXJLGggYIjGuOYlQYG0AyLmcQ72r4jkHLWce5PKHWOkaY7SKc
lz4yIhqG1EndRe88U2YF9UWamIzhVEhbp66FLS3YF9KG+OSe13yd1OttM89eoFCP
KYboa+h6z8UKzUWkS3SB32hm75HSehTsemuEr1B8opSVgQ0Bd5PR/WCon2f/HfCi
PK5bBxa9fKkqNOOUXBzFeqCl/bJzBIMLSi7TnWTQ9Nv0TwG/j35KBIKl/EhMd5RW
1IYLlGOGeoO/NBEa7Y242+g6tKL9kJ1GKf2/dFMRi+R0pX0P7ZMo+0q4O19Nqa0i
uj6/8eoJiY+1fHvcsa8h1Wips1Iqgt8q5H8OkPxjztpd/kRYLPOnAiDq5dK3Rua1
xlFx6Bnf69P7CEGLeqxhLpENeW3J62DUG6k8fXY2oqyr3Yynx3e3T+phJ5EOeupG
xsGzF+tmjSNmuvrjsGAjciRsc9bpnQtJEY2KyLxUOW3I4TegAHEOWj0HzInaBsoI
KhStZCoSe02SDRnJD0ULsDxhLBuh7sXJJJ+dDl+lmK9JS1JuRjiRl4dP9QrHAMAW
TlBuuhayrDfYHwUbEBNqhmaNhoqpfHOFcR//FeTMKtUg3+5TwSiILvy0CuES+cje
yj0z40pHln+M2tCc/s5UHglk3YFRjcTlBUvflpVY+83IzCORt8uDZi4yqK3TF6qb
m/xRGxdva5LV/Az5ckaiRTO7kyJaPt+QXMSJskIV0Y0X0ghFsX0QH7pmf+KQHfN8
RS6QmL3PyRW26nMN1bqFk1tHGS8i16Z3JbvhInvU8ayN/18VqdKfQXq/hBoc9Wwf
lrP8fg67d0NLlqr/+6u3IlpuYLsT5uTBZWyuAmPISnRRaSr6Wqym0ml+SWRIhZ4a
UV3e9ZKqHpmqysaxdksDZwUGPGEOS450c7LI+Y0SMX+iXbWdc+92ghEDu5TCMA+Z
cR6uwQDbf+t1gD+h5f2fmTHCBwuIP9nyIQQhnR6L5arN+SXk4BERF5hOIo29v4av
xEs91iyUtUJXikd/+j4lUYt/6FIcnKR3ZThB3wtLSgKui1wUND2KfvrXi2jQFtpV
ggS98OvUf9NIaYcU0e4Z7tcITkWkLy988fnvgY8yO7kK3okIW/ndFCzuE91W04ya
AsNcGPeDQQr7aQOZtzNguObnQUAmhf6T6MSZzZOLYcIdSuRZHNggn//5O+Jranx4
F2G9WAaGbkRle2XYm3sf+97xiIUxLqfG5nr0Td5Jyav7tNISVgxnzHQJFOXEVNoo
gq9CndINuPelv+RhHmXNAgilWvjWmJicZ9xQe1dCHGLXOiz1BcBpm7/qVfkgSbNJ
mINu/crTiOqcCIell6RuTuTpO96c+q88pZLaSl5y7yFqt1FqVHMdJrw9FOlpq0+j
OT/t4OuFpoA/y/drfSRyK7NHeM/dfTp5ELlLGrOCG/I3YLLlHxiO7jC92JnYUaRX
J3AbnjWmLfL8jjDyXL8CJm3c12N2exGum9T5hWpVnGQ8tDBP0JmfArIK3Opg2Diq
GYtr1/yPlpyCPa8K0QXmlDUxvYVfCKnerInLMZ8O/P/A26o3DqSZTdW3DKdzXh4m
+UOq4v1Hf76EmDIJNpdfLvAcBJTkVFwrVhG+K+Q2gyz3wiUdxbbtRz2ZoJIdMvk4
NvyI6aYzxCDv11K06KfryoVbijRqF37zbjrKsso2U40Bh4jA0WAa63O8x8fZ5yf4
3T6rR/pID6aQouAwi7VNk85K7NeSi90G5tKSdJ2PHW3p8R8AY7/lh2Ap5w3rt4BP
9A9l2/LnENBNrKJIqAx/XHShC6ljRAKy03LFHfnOSWaoItLlg2c+OzXtTH+llSvM
q/5rNbNq1XOrEtA/MirdcpULtyvm56eq5A0ZR1I4w79jDYrGOxQegJ6gTh97VRU4
/EeBYNP9Sp0ALGqYRKKTHer7/ENmsGNPmdN1Wdv22as8lJIm3kvMHYU9gq6qP9Fu
HWDdUAiY3/oSqOCdFnXp2a8XJKl00w+5P8GxM5xneJ2vYhnEhhv5kh6XDbNtIDr+
rNsjoKG63uDtaI8Frc7sRnH+5czQMZDAqzlecHp7v0z0zccpFVlt5ycTmEXdn8Un
RpttjpgzBaxiinmF5P4xn7XKzy7Iq7Hh81mnC4ut5Tlg7gqvVQ5wCTQmrtGsfXme
kh+1jfKz6sfxr4molGw8CSsVJ1X9diLUKkYQTGv57E2EBtyKSwpZfx2uAhD262Hu
Tw/pselh2h38se/1lM+ECgCvF51IDo9F/g3ck7fOGXFw8cOZGbKdDsO56nkX3+Vb
ecUycbGbMTg4UxeJqRIyHFsZRAswe290t05lFXw+r0ZvKuOburpep7szXcY9ppGn
PQZaQnAgA2bH+6Jx5SwQ7T/4Ui3uxtSIC2J3xHss8COBVyeoDOfuotfYHrMiKOfb
CZMHmrmmuMXC9BeFEjgBnQOn8wL0YjZaoEE4oRcBRyTy+BJTbg3aL4H34F8/EwFb
mbL1cYtpzMQ9dyc9o5YJyugCzhh+pnrQFkClzn+zx8As3puN5Zpr3Sp4F4qUnk2c
xi5+tsBGq6eOzhRTGlEdJfJf+zVi/PlMV7l9B0UgCbmLdqlE8MHN48baTF8sK6f1
zY4Q3sBidk1NrPn5JndvRJAIz/BMQz9qJpJw1YWNbbS81txG1+bLe80c/IpVuq7Y
1XdFe0LNJQ3BcEpw6TX3rZuXoUObTjUOl4kusllIaeBM1JXS+YU4EOtM5mk3Eqo2
vOlIUVf1XHq81i6FbWqRBcYi5QD6EtWqrs/+FybDjw42D8I7eT/a4zVOMsaDl3Qr
Gqnq/h/F4sl/vJNdAB5oIOzAib608eOfC54vE6czOvunXFxspLco2eZ68fBpQBpH
BlcWP9iCTSKGkHCT8YjeMeQ2tjqNUTzZv5vVU+WmRJCxzL5rFGmNY/Zsg5p2c7qC
Au752wWUkRMXMeN86XPC/Z8fpy9gxUvtDrlqeUckVU2oW8ls9K51oJKNtRHvcwrv
g5XbARqtfRxP0WGZzQ1ZWQtjtBxXm+/kn7j0IwAUHtJ0T8QhotvDs33Xu3pF2u2+
yOmokNL+th85JVkLpCnIYmyR6yNBjhoSNjFZjmk3As4wkv6DIs2TRzvzEv1oTEcW
Hv1SYk9CpNO+erGqv8t7o6L2lpZ9Ur5uUf1kqB5HypZxFIUyq9GjEU3D3p4ul7+n
JuEfwJdvh4a9KyrtASlmZYVzsf9Ky9tC5wC2UECyZVP44e0FwlPLD8Re1W2Hk1ZD
g+QDneqWQU0LrJPdQcqdwPxYtHms9fi4y90g8qblwcj+k43Iun5T4BKF06qrdjBL
U/4+ZsKYLyN3cdQniT7NjJhb57rgBJ7twb4W7Owv0t3Kt1CnDq5Elq30+YAgxWUw
xPjAMZptZ0u53C5cC+utcMN+E/Z6UwK5O6SvWDrO10IVOy3sEMGDd5t/RGh7wJCH
XXjwxo6A5JPcMwyfskp2i901o6XRZTU1zmy93hcaRQ58tm01AP8y4ozw0QNZJd09
uaqzetBbtHalBOLuUIlMZs1z6dJ2lcmHAM2WV4P2Ek0LrC8OPGH/ZqySTAT/KVi5
LAeecDiM/VH0Db7BlBIgo4CpLQi2jmoQ2NfbheZ3iRXcM2Nb2HyOvPv5T6O26kKd
66ZhLVauboGjjEhSljoebbaQOxVHO7AT7PRGbBISpEczEuzx68pQREixkgFeKGPc
K93g5+xO7jSeutWCvNjX7JGTu0saVDxCYRCQP1RyA/CyHCqfW8Z7A5AIwYxp77BA
rsazDmk+NmyC0lyQ4gbEueTuaeu3ehwEkJclWvPNIAFXxUCUn+UPF65TyhztqtYA
lIhAyoKaS7RmcyUjEBNWm2aLUInuePHY5NGNBFhPqZ8q/jS+PfZm5A3WBdW/MSmL
MqTifJ34M7t6sHSxUDSy2xBQXtRVPF7unzVzJGbqwjz/ELWzaQuzGLzz33fXUgBF
+f725KUt5Ot2cB1t7RIUqQZLf1D/3MsqyJGHqeBrv1GSr91TO8qbIaHf2KNcjIHe
OpPOW28FzAMNw5mDBkt7TEMn2OoSAQ/iH16h1TC2m5SxnprValtFwiBfITI/KZyv
BcTMYOzQLQQzkl6jbmEQvRR7QAD3ZrowTe3Me91zmHT8DqGTbz4lVkBlARJFp6XR
fcIHgp9AQ1jqoclcmnqI4Owgdn/QrPvnuc7F31U+g8cqSVyikdJxP+FktuhUOWL2
UF59146R5UCaOsPDNlbBMz5QHkDazF2DJOMNz7TkpkClbbu9R7zSxVorhyT7mGD5
fJaJpev2Cl2HWveL7iO87LejrWcrWQP/QPRvj4bNamXC+x1glGYfbI/+88quvaix
E88wE8cv+7AcAAEjqIsp3bXf6ckaKBxM6iJD9HiOnYoU7OcetRbYn7H9jDhTVXUI
0J0c2qN8dp5wUZwKouj7qwLDWQWbA0RcLAeRD7iEheu6VAk8ostCG/+lp+E96M5s
Kp6KlkUKakQf7iH5HyN+7hDu1/ah3fEpWnDdaBcm4ym7VN/8rAc6qlO5iaVIyRBC
4YNRhkusQ1eIW87xC2uZZ4H+jxcRg4TvuaQ6kT9sOliqmsuJ2fgAAL+bGmeefgGq
fSf+UFqpovC5eXZpEKroNBD1Wp/8QMUGqrYgdzpDvU+t9uggQJwpfU0wFHSRaXOB
FOwAdjhFnL1LwPZPrXlmDCgKp8jqw+9WlfJJTMWqiJjTYLU/kirYW4MOZqCR5U8t
N/cUIfmNIppP9pU+dI7DhnshUjTcBxaELav6rA9/0jCc/ujR/0VE1TeKw0zKoFZ1
uGSwmfIai5qRYeRZCziDG2yED64ls+4EQ7bVZoflD4a4eMePmGvsXKpueqTllMDD
RRxCr54Vv6zzTGpDix35XAk14zZdueovxJ7yOW6z6h+YksXIFWYTaxo4eskU1zlA
lT1IdLgG0555lQA4yrERUCf6NIXVNmUIHnCojwdd8ClUQN2fWQZrXGaXB9rwyb6L
2gwcWQ2FzFq0ZIDCKk+p8jcNVO6tGUkQnN4S5EeCGgCyumeW/pWmWgzYYjzOqfS5
WaBv8SSwpYy8cHVQYLFSnfewaxvvt+LAEE9lr1jgTk6U6jA0yg6mOUnZsDMqE6ZH
gSxWFH5oVhxs02yb136ubzXcH2nskaH71bx9gRZ/ItZO1RrgBflGw7IyOITeAqwo
anurTP2HGdvRMLYZZEgPRgwJeUqfz6qaKdgZU3cTGP0eaHP2XieMVSAlpMA1uhAJ
GUufUObVxioaBRs+JoU5usKU2/pgUw0Ppm979MwGeriNVbIra9+WVSqYOF58BVzo
Jrhs8JIys8CmXS4ThcGrd3GUaxXE+HnVsXV3N5UMfGtnIbHIR6AIlCWUX8hX3Qlw
xIiBmEjTe8NjYp1pnRmYubdvWbpIlMoGDjJIQADatduah+xL2tPrvWu3dXq1PdsX
D9tNGKOZxTBKeOrTVDshdez9CLDReXfrhuwOc+ZnavwDUrTvyBuRMYXBVNAbLfoH
XU80Q2B+iRhT2Ly3D8CcujykOSCA7ZX4qPZ8b+OT9Ag/xfF9Q1xzRpfq8QCk5k+M
8EwMHT8eVdrLqk+5ZfjdF76Ld08Qb+OakyOA+wE9dG1H7SU6ZHE0gcq0MaPGXblz
/r3yt3Xkn589W+fE4qKlYnRI25AmQFXOjjE0WW3YuCSKvPezSo61n5w8djbSzfE6
rKDFoBpOomK0Av3JWDgew0geyGDEhLWSBcOg1TPXT99pAwGz5CWwpoTTEUONN7hl
I7w3ICLf4eHXZbV+9JbaocDncfa4K88ZSu3Wych+dwwhkKOmJ+/J0udVMUz0w2uQ
5rF1Oee7FGMCPEB3dhg1xEgHILqE6Q3b/OWzexgrKF6Xm0XOcwvsVUMcKttTBDec
Z1i5Rq747w1iPs2NQV47ZUzWff79xkNiPn7Lq4ETukpeSuH2MiDbJW36O91AyY0W
qJtGvSEG3GxDhdw4tX/429ToFe1fXYEHdzXc3Drktu6CbvYqXbRcNMFMB0302Kwy
besL1djyQNyy3kwq+rDlXDN3Y9Qpou2Nr4NBBEE1ritot63sfPIVdlxDWHWOaUmA
VBBY+2EwzHw+MD3aUcapDdU6qmAhzzogvwlEQlzc5TPI2r/jjNYAnX2EnvwV8IxV
Dc0gz+eJUMmitHS/OUeHJ9GYfUnih1kvcWPKSlzeKAK4KbT7dDyx35+NDIEdOd0h
nZeuFhUtvxDXzf0VH65Y/9t5jhRVejqMILfakC5O1kvKrvkoB58EMYs7N2EBM/q2
50FLBb6m0F/xv2ngZzadhKuycXs7HanZVl9AYMratzxHuJEnwpAxNTI+N+vQLlJp
q49k6qUc2BHTOovq/KQBuzzsLsTAYhQmSabdWIa0Py4cfrrS7jArKA0Emm35U4xo
8fKRW2Wme9erGE+hgrPx8e00zxQcdzg8GCHINnffcRIYFBQV7fSu2+AsEB+4UWV+
MeiVwY62a8do9v2boV0uKf8M74QcULL+J0zUszpI4NqSI6nZPmaCp4rNTr9YPxFG
stN8sSL99WPy9jhI1GKJLNCRcE918azi9SUK+fwvvdnvRY4wvgtQAtd2BT2J3RB4
YIHGbzcAHwEWRIIhW1SRipdIsDJpOzud3erDl/A0pRh28Acj7NV0paT6GT7h+xPj
fMHAHitildKRSthF3iDDEPrzAeF9orR6zRXYlHVwz1FXkAiyqr1BEmdtB2D5n3kU
hmw3tIBQUAJxwjZsdaSotluJT4btjvstFYEU0ZhYn1eQ2m4xyevfmm/AiMOeGt3H
Vcdr45zMqxXPut+uYXcHfzG7brZ+F99YVxAhHeFZugIFZF91tg8Cte5GyyIJO9hA
yRhnSbCWLJsMcuZuBdwHjSPFyVGAWTngwRN42+jv4uTxqz22f2XMhRCDkGlL7P9e
S6myf+4wABq4beu+x8W6YkSlvTemVbnjGhvriYc50ttYKBL4BQ+M/0glOgBVqMfY
b1a0x4W9e3i0TjdUPMlJaeGPUJLbepmSRxijuifjbvlCcYzlnpNUcqm7Mf3XTaRk
DVxpHrQUOpPQ9OxokhAsrVZZ+fH1RtTOa/Y9r2rZaL8hc5OwqQg4gQZvle01vPQ8
hUzhuFtJtQgoAOzJW/QrjmE/Xydnr05MEhD1zdHrxivZ+e4Ia3he33NVhFoS5nWM
HEgulllUpYIHrgTn8vKN1WMabo5tXmegSXFWJdRtxzahxPliM3KHkog18eUNHwkV
r/iDcDLGw3bxrujzRxvCqEkcTxZVVtteO4CzlO/ECw9MMzjhSbp6uCEeXq7Socjv
21yqhu5JBp3bWWk18qODN5OZ1yIMbyJkOAviyfmT4ZHBFZCTke1waQtuJt5czZUL
koUFgybcRU7rrE8FjV8egnuU4MS6LNLsUEw3VaL6MUtLwAkU2FarxFmEIzSSc6c1
shovkUfU0l3NgijUW1nyu2WYfMywHsUu/LHhV5e/1tE1nP5uQj0vrtK7hxPoXZwx
4QhmEY2lSy1aU7zdspe9htOBx+ZZyNAYmsWePbr/xKLzy4dsfnKDCfv+lZ+rtStS
9L3q/5inXN6AfmtJSyPrsf9dq4sThW9KhSjX6NvLEfbNn2wRQ3+No4jhbFWlLx0Z
xOGiyrs2vvTApwwylb0UsAhqk7rl6nCEUwjZ3mEh6IPiWvO5Uc6fBu3lMXwh6+i0
EvVzJC8QuBmDQnDVoDuPK3Z3q5PA+NsD1skHux85ZCeunOOkrpfXdo6kr25h26cP
xVFtuiODD/hR5aXb7Azp0eS2Iw7sKt8rrkVXbXCVqXXHGNsKN7Sbd/gDc4fjs+vv
UOpGR7mQdydQD2fwVKECTB5j6bFPHkeHFTeerUnP/dhuNl995qZ/DWQz9iFdeuDD
y7QFJu7WwwZmqylt3t0YWg+vx4HB6MVi9fqh8NStRcJGR1upHTFucm87lAqxnK6U
VbrLIDQ2VxtP30JasfZ6FjhAPAXhrK1VbbCJoBjnSf555UmUkaGzs7zfdD18PR/2
fb8d3EmAEchC4S63dbbl728TVDOQtCeht0zk++2rUQn4yJ3K+KG0F9RQ7w4qiKrS
PmdSwM+Dhg/nudv95lbWghLmB2LIT+WskHRTo2MJNNTHb2F8DJCmAZXPfr3VwPfs
Uau6xPeMRrRxE0jEAdPsA7HauF5g/+i1aZXFt8m+nM0u1YnmV3IVqSaYKVBaH+XN
/HsR+kZhfJ+OYrmZhtZDrc2ksMV/ted7QsP3HXb3ojLn2OmbZ2aIsvY6vrzQhI3B
5iOi6ulH1YizxIhcQfoNj5PZe0LOYj1fJGrTkVY6qrnoc9n+mFExKrFHukdcD0S4
NwoiT5rMXmsWJ029dJdC4g7kS4Jj8cGOPx+EOKOaHpZeGHT/kkOZ1yCMh/eqoBrQ
L1nnfU2KLG5mxxRagWtYh1FnA3Alyb5OevUUQn4sGhI6aEN4mRoWpJaEHmW+2H4J
pg+WtY48nYtfhG7tklnV8cOgJUQM31sQsxr4yFT3uxxhufndox7Sqlk5bAL4FazJ
bWVPk4eX+Br4U4IYUHDuKjCaXJ+C+MjaNgJ0CKUBr+/vMT80PPGhfPjUxsXTj9gR
2RUbQbpE9OI3fZhFDBBB5uzH2k8aHicqooxup0Su2aYM+2MBbe6oUToyY0XZXEKC
0GZz2qYZg5YknKDuuIuBqePElCop72i1GOVAcXeRufkCXciErnZb6yvesrjmoMeu
dEqZbx7WKh7M7zbshBgkcslYveE8m56ZrPRW0RABbbCJ8ZxM/fHICk4NMXWaAwJi
rQdaooEX5nCW4Wj4e9jK7ud6CXv+Bw3dhPeWK0hJuhcMi70Ge1UBNMVxVkZ5kZxu
TlhiCb/wWsHPwgPnNH4cZlCp4JcXgAhuSt/WVmuZ5cro2g+ogYskVk9Wj2N1Klkd
anP1X9+AtpLdbRFJKJPvVtJ8AX7SCjiyqswpGntJH9bSiF6cod1T7l9VOEWyB248
U+yh830TxFXSbeNsetaETrN4+C6GWxvsacCNFg1YnPNuEn9ZH7APuHKwQKKQwWAN
IYQfPbnfhFLNaaSLjNwZLPOo8Wmtjsn4iDR26QVKdojCL04Gjgzc8BuPnEKTQFeK
J2FNeu4/M6bxlvPOFsylhqk2t1kf+VW5wIO8HW1hrZnfAj/3CibtAGwKpoajIvK8
7RcH/snnMyCwlj1pMKhiYfsI6AYNcTnYixsM8NXnNiHJ+lBPQ3l8rZaPlN1+TywM
EPdAgO3gZWBa/OKwMGMQFmSCO7vvb0C9U77BwgS2cpJnpTgu+INzJw8/QSMXFjDm
87NEgCj32xyQfZrnkNyaPBdvU3GbLL2GZlkx9hT7dt7aD+Jy2kxngoRTpX4KIzB8
tqhsau86b3Pr58YkIiYvJTjr048Ao+BJgq7VmJQoRdmqDGIdPpdJDnCc7oLFLqgH
d+HLz6m2aES+KXtQOJ2HMWic1OV88eJln7xntdbe1VjTB4YFqAkmoZDau+JXlrpr
d1rNdE4mlWyySmj/7ATbOsAXR3gdz7TTCsOYugs8grZWtm/Uuo709feZ9UdAT8OS
1LIh4PhcIhGYfVu80+Q1OEGOsIrcmqQgitjjjmFVMwgD2yPIcqoCdkW3w/lB7CvU
PSsGGtcBzaSAngQ2XbNy0+fwOfbLl6/TJEGJZi39pVcQ+9+WqDIV/rn08DHW1Si+
QWDTx94bK5ph8Vss06zMPEOwPiUYQW/+b7wzfbBiP4gM+ozacrJZT44vkykzgpgY
9CG1Bxmu4ny+EpppmqXjSZMTnNt6AoWM5nSuqpBCuS+sVCtolZkuNUTngJFZ9DjR
xz+LTI5y6RUA/fHYLvcEBvAHjSDFdVXCv8c06iXR95E7RxBFdF5KlFfwCG+PzwEl
tq5PjpnitmxL+15Vd1wvJfMiS3/Lk0S5hveDNWjpROHd8Yn/z/7gi6AK9nkEeUEJ
7+EEx9X+4a+/c2Rl90Voe6kivWfjU3HWmxAaOo2UM+shqVrAKQqU/8mPiRy0n4ZK
NCjWydYFu2A2eSr8PycWLw7Q1StvLNqp6UlDukgtLwCpZ8IPWcV/WKdupMdkzhEb
qaS0gDLrhYPpxwNwx/rDn2LNt90JWmFonjnrqw7tZLZfx81rnvD704YvOk00a7aP
LC4Y+Zl+PSTau3eypQ658jS/J4QO5OVIw2Zx8kaWwyLyPc4Q6QLtv+TLyHCsOWBx
tBhIZcOhfvxbQCkBgHHrVkkeeaIeA/GQtsBm5XuZrIdhtxyt/TQD9T8D/bU5yiFl
rZbj+sZddQoBdny9gnTwz7LZUSJZjexLQ2mlVw68dLXoeC+fcpU8io2H4sil1sNj
2TuG9Ow/M+MesxrlG6aFclNbAeoxfdHiktScNPuDRT6fa1dd9LS6GaK3ACcGwdK9
eqQe3YzOFx8YTrri1i4RWvKYtdmZzZVTP++Q/2cSwqwK3F/bI8H9oEilLVfeXsJV
/vUO3hZrLaxu7mJzWnGs8pmudIrU66+Kl33Mep9jEL2ZulKL2lHid89rQbhjUlpT
aAV3qNyF03fmRwYNDLAPwmvonyyPMSCBLJCDyh/GIfNinIJWQKYqjgdqxPIA75Oe
h2Yv17Pm419UGcPJ6HUgQYGrS7Z7Rc8cKnDtL3x7Itf75oJwfF9Js9p9A6ouYves
TRpBCH1bJi9gu2P61sPjld18FAxNqBDobZittcQmReR/z/zpBNElwNcsbWew9Tvm
M8gPh6zIN4jHp0u2AfbMKjUZkkkNFtUGgjx1K7WKPlK6Q6VVqpTUnXRcbGgaYrxA
wUCTM4uwJBfnrfEZ1HhXNvIySJ/yFkYe5H2/ujw327TawVnr6BFlGbp4VSsI4S+L
YI3bRGApURh3NBquhCgYsHhbASJdWFl0E7X/AJzVl+aqj+GrhXx7Hf/lU4ahvpr2
j6Tan6gOaTd4S4q1cESjriycKuhr4zdqmlhCwdH9GABYKW/YvdIHPpDVGR+W35fX
saVIwFqOkdh8N2EmzM1dvYJIeO0doFqDypx2VWG7yc4ciDAfzPHCkxQdSR+uuYKg
yQQZsmvosOD83lBlO7tn/5SqTXk6RUkPBWKBze5FQmArRFbIg/O1XFE5WdmnY2M+
CQg03dgRl2GvCC//siprrD0n0wktMnmqRBTcjL6zWACqp9N9a+Buxlpgd5v9274I
Qi1PrmkXop99VLpm33OHagRVR5uw/Dibjz3j1lIzgDh8/5E4xNkxt5xJeAXVdLFr
aDvNlgo5Cnzlc8YY+2qMp4jSkjGIEDRVTwzoUWOXZWD5bcVrLATUiKxlgDhC1sTy
6oLbS8/OvvYdQZEhbbOX2Fzl9nPTY1wTYckljCn6dW5D4UqagDtODhtONUQ+RlNY
fjiP7xTJArZQzYJmyqoPj06URDgJTrjdQhs1Rd1KsC0Ocjw7wM2qC3YDYPabPZq2
HAfGKHK7dv6B+XL30vhi8NtSfGhthqrOicrhJQJCgsH6IZDJLcMEKhSusiF0L8aZ
/cavy3iLJWPoeDmER1lS0+sO0TwlROS22tJY7UwikTO0AtJulFkNOyRhG1U9XYiU
QDRECPvHJ8HYh3R/QbT1jyXXzE2Xf4Wr+ZfEXXqZ39k83h+RsH3OatkalY96muhw
GA9CJzfeCiKtfaahp1/nISYJcRN2h7DlV9KfJQpGBUND6xgM2DDnpmt6iruHJ4xp
8J4nqMF8xsmCdgxdU6P7KGTbDLPjZhuER3a+pchqmAJqrs7IprNxXJxU4RZ1x7On
PObL31og3giPg52bzCylQJWBJ5sJK2+IDgfP+Y7abr6gK50kg7tpmgZAg0IoHA7b
kjQcC025t1+aEj8rr+2ntOEkm6CxudLF8/MbkmOZuGnLvrxRn8cP0dJIfUfi8IA8
bRnF3HW3D9nnfh9YmbyeXtBtSHX3CScRZLuVMHx333puBb0tlL9qR3OohEREhySR
1Fn9kVNro1xyMYRe5BAI9h+VKrrM/a4Hzfx4SN9joRteguHeCi0JS1SfQyNqZ5UW
HtGA/X3eUS0//looyGIVDY0OtU51srpynAXJ5zmvUhPZtPyFNsA26NJlhtGcfa2s
sQs9h8ek5OFuL+Dhj5xOHEZFaxOcaypGHueCDX29yU7AlwJ/s+gbAcCMcm0C0IKm
ybdRchyIlou5RlAbAHIMrZbbLKDBDURs2EnZtz7d0M9NJ72gzsggbD2cz2cF0j6g
fSJpqZGuaLguG2CaPsMhvE4lX1xpVLLIU21izvedP5OPVZDSwJ4AOtB4MRYDoY6O
49wujMvAALWLm72DY5fqZeuhzpVwn0aX+kzLrglOAPzxlqKlXnh1frtkkSahl58T
WSH5uGX5vFL0CZNKrFGY2i+OP4qwhPHgvjxglqh1i+jQ00KQsPEUbEzvR2sd/jRU
ZI0Zh2PqJYEOomLurrKcvgWK8+9W46Cgr21LOn+co2FzgbyfijJYBmBznfEfvQPU
t3ckOO21jxnGWNC/xgyitl98GSuPtFxEg1LxpM5TWh5bc92PCLvS5Z2Vv1rsbzG0
KInbFFvGNC4JM4oqHbys4U5QX6GTUiiJyJgjCIYS7JBDEVy76vMrY5vB9+GT/n1T
iOuPKyyvkUrxoc0UPiZEbbw4M1yRHMeOIYZtAwfesqMppB1aE0u+1xtdwapOpk1U
ZlPrHNSV/oDF+0miMJY4BA6YCl8TkpZqm+ay76bHwKkgzmk3VNcV6JDKcyCu8uOD
mtyVv5Y1Q9q+C7r4vX6Qny6ALTKJmOiqC34s7Yc231dMEm8qxjzEGuIASK8tm1GL
RpiWG6/Enr7HxhIQ3DzQ9C3y8bwbmFQk7MF/jdk+z1ENu5z2ap8/jB6nOrvtGtfw
hnTiWkrkH7FzeiIiKH9UvTl1IoJoK7l1Eu4oz3RxR73maYUVfHxhRpEC4opAI7g7
PfvV3P5vQ+XKyya0u3gvXev2E09u4mr+Lk+j2xeuRIr+V6XRJIAiI00LZdAbJpn4
g7OgMoIMyR0GPmmBW5ebRS3Ach6CCZzh8bBqY+bRRXpshZrzBq4NG1p/RNcsR2fe
q3E69yP6ZR7ot7mrpfdB2RZMpqcOr7v/iGeSfJQTzAvK4xim/v4gYge7Owpr80Z/
p40jg0a5cXBaF/voF58Qtx0qdgDrVp7XGIie3cs4dBw3hVHHyxOilUjLVnd6h0+v
67c/3jy1ne0rPHFuZSqljc40uSJyGy5gaYQk8o7QI8oTP/PP4Ry8RDiiWNC8ZxNy
o1vcGYY1OG9mWkkJANIIgP+K7QNMjNE6nrMfS05RWIjxT6yrk0nMBB/6A6ZqjiaD
g2acQrJtEj5ud+RwZzvQQqNioiN/svv99GqFIZEDzUbOIb7F72nhr64/1Fz9aN6T
WZfQ3bzCpBGD5/xaKbWVxxrj4aTEPjT7Kw9PnFf0sfRv7tDt51pRpQAYawuYk38k
xdGNHCyExn0GiFTLXhmBL5Yrhqbv6ZVekfnTxDKkAiJeGijSC2vK2yyY65NgQrnm
/nMKkAl13FWU3HHN2Bw2OSQflQME/W2g15vQvWNs+2f3wwbXk2UwQFHB1kZIQ6zB
Dpqwx5wWWKkqeOIHT//Y3HueNuaPKzb3Md5bSn16kVQsd+jiEaG0qdpI+FOfiT7F
/xKsN2c520Wf+SyY05Vryv4X1dBIJ0x7vfJoNmUcvAVNaiMA9rgxr5aqlliWaLim
ogZQylY2Kf60xRU0ZO+1oUF+bN4lK9usx8lre0lOI2tRrL8ghJ8lVb5CXUAldbkQ
s+oAXaEHM0MVm61s6gwfO8Atw5kIzKYuvwcpDSrH36VuajyLaHR2IM2Zb8GplKO7
sbNhYgjNCzeMK4k0Blkm2Affy18gxyC+riBvtpGhAseQpPUcY1eGt3eXLm6wiDGr
sI21ZcbMgcdemxUZWQ/2kJsz6VqsVzo/wMHE/7zagg7TLI9zUf79YnPLWHj0vgam
pVxKOJe5RoT84z6xql3aOOop8JDNsKRwh+kXcjOMvq8iZKiZk51d2Q6Xy5rgB3Pg
wUw4sQWvvGwa4lJEl4Dx3RM5+pvbLbbroUUQ1g2Mnki7BSAoWGviTzbaYHFizUXT
5GH5ISkwDsWwcTcgQd+ijemgNTNHYmi12R4022/PxvdKVaQzHT5Bsi/6i6UGo2dA
/XTD7v8AwfgTcJIx+ffoZKDhA2dl0uxxYZTAOhM+gwoJl7MCGZ8fbjisArqQT4Je
MvS14uxyB/t1SNcEHGeWi8En5RY2+EBFU7MaZAKy7lXIEkbwifTY/VXL/XIendg6
SAOwy1t7uRbgi4DdvsmKDCb+by1bt0HN2IYwKZdKY2e380PqFiO8PVGzZ9Qx1W89
b1bJ0sw4u0tNs0s3qIqHxxq3Rxmq5nS7Dk6VeZAsf01NrdSYLUbBRG2kuoltPDLy
mMVeZCEepdPL0EOZmxlYhywOR1Rvu6hTFNviuDFPu1AAms5edTSO+1Rkuh9lMaEW
HtWEN8jezaELbsqblhi8Wf6b1bVinkr4qQfw68U7NNaPsUlv9bwhV6hO+4R92UML
cPQUzE70Ap+XVstBtBlsp2Gd64hBQQlwNYqdA0oxPV6Q8EB8yYU0/EpVmsMtJtdu
YeMwSRJKiWhA0Z4f98n5zmnhO11CaJWRT8TMtKwjSgoqFkRIe0U+UiosroZ5W3/N
yg30uLWGLB7usyXBQZAdB185pBUCKA0RTyRO99cmPE6KMUjGToLod7vlx1wHIUO8
w/UtR1wNgvdEjZImyerAchSJWtQZCOIerLqYjn+V4QMUEZa7fz9agFp6NvCnm/cP
KTJmKsvygoVgFuZXlDQ0c87hzPsOdSe1861RXl3wmjpDPOlwyxhLmt1C1dq2clIP
+x3YmRzsibfFFANBOvc7qOjJsvjUkgOim1yUL6l+a4Ty1XaEBzax3zqiTYQMw/Fd
kQBLKHlB3l38QCXGL1ZzMCVgTJHrNUs72SGDw0mfYZZifT9fxHqjUKqpJrractPf
NtJ79s5wgMzY+8PNrs1nWDJxtkzcK1bQIuwSohwDTxsW034yvK32WNOb5rolte7/
tEZRLu7aKxJLT4YrQ0fnNpXpEo7qyxr4DKQgqXHCgMY6Xmj1aGYtKNSBwwFISOm+
Nnokb8DKBq1tU2ADUwrwKx+Vj82A5RHQcDo960WHWnkMg7M+cSqtvJNDy/ShvbGe
iunkLQas2t6gXe8Ny5Ad29DTJ50a9/o5YAILpVXBj4a3NMA10Lb/WDoUt4pF4Q3b
3KkCOVwL6VlBHvCy6Oh+AFBIbJB4sn+PjvWEuqQoOOT+2hYsufj7O56S/VJQ8egt
rA8RpjbWjP7YkHpTW1EFNrenMy/1Q86HN1LoajVrSEcaFG0nPA0UQlFnNLHTYPHF
f44WShGizNHb5+krP413Z3azF6QyJoJn5mR7tbJ+USCxZ3AWcgm2rKVkHMeispsL
0AI5oQ9IIxUF7DfOHfT6rUEc370id3C3ld4U4/VPJKPwWj3esctCWVfOmHbCtKpe
pP4IR348HchpGZ6UNJquPYE4qRiC52UnZT8ZrRAIsqR/NKsu47+UPdx58gvcnWdX
vmq0L42IY6VTlR5fmxckfGFNMKXRzNSfM/Kb6lzHC8Jd11CFwNfuIEj7e2d9kPZD
phyu886Kzmx5htU5KcZqbb6J5eOq76GOnTWzhQBiVrP5Flu43bL27ZeBkojHtN/N
Jcjlt7pLgZfOXceOPQHNhxAhkgwgLvnwD9AdMqb78eLxpRqCpIINkn0wj+vBQIyu
eVqOH8vEHW7q62HeQHWFk+ReVWUJRisomWVnp6FyB7UfoeFevBJO7CHTAfKdW1t4
QDiCQN7C8lC3+LMg3fAp4N5DNhcO6V9CR9wbf+Xasqbf3Q531nkeGeCiqC6RHdxt
w19DuvhZUL9BN0oxoB4KHa4Sc825+mr8R6scgAsZvethgrZ9IZE9wwlTg+F1xfgF
jjsObrZjDDy92qJzFuEvhLj6PAWeVwk47BeQ5DMsUtNe5DfngWU70vaoYQ2A+VcY
rvXXpcd+eQn6yechCBhKpJ0kGw5YgoYuHiRsvQ7WXRuHKjWgh5cvENQG0DIvz4BL
nE3ZhYpdc+9Aj9T2D2UMnzM2eocRpCFXxuF20WGD4oFzw1wMznL4iJOqm2tLceLk
P77dqiQlH/rB8dZKF1AdIM7r1rnr+3GYApaAX0kFPlBuAKXBM8ZNq8W+MZ8YZaGh
OGb45KprdMOs6LcGXnQ+DKq6mZdE6O6rEaSoTNoD4QQAYyRVJNzYKzh2mA6wTyqA
PFiuzaGsY4oTrebm14AGJmOJSPZoQsiH2XuvgtcBLhSlJ4ELlPz8HP+gPPX1jEeu
uv6mB6cM2XTHL2IWE6qr+D0fXO1kPYvxDGeA2xZgK481++mU7CmHfuHXy2IR352l
fArcqj6rbx1/eby21F6ue4jqfOSrNNg8fgsFEBqnKeGQA8rSk/HESq5IP/1b9HaC
ucLRdxSW/xr0Jk7j42e0lJzIuU5PTRrVqKksHsCNyrHZVNtl5E418NaiQ7Yly9Ds
AJx38GEhIlF5DWFjuLwpDMtbPV+eZzs3VcxOzpXkfmmRoCv9+VKJVSnZyjJE1COH
N0lbASjDZb9HCmE31UCAXEiLt080NWQFhuKTlwChzwcQjUuoA3+lbng/gAWgt0Oe
PhQlP064jcIsq2NFMUvBJAIH9p64YjB7StV02KoEgGB7rb6kGiIaAlRLZgnITYUB
YEGj3hOhimjO5Z5nhm1wWqtDUSBi171kr1ReF5H4Jl0IHfWO4Kfn6BIc5iIY1Jnq
OkKPP2MFdSmZb4fZ94uE7zn6TnwygDiJraAgVbKctbmZFUo8GPizjEr4rrRR0jUG
Jdk9f/KAxlTOewC16wsakhFdizeSraZVcRptzInhRWoIFYp8Oo9ZQJMNcy2osoKa
jBqs7fpQoSAyzdTVOpOAInEC/UJ1vYpjK4HNWYXD8b07TR34nz1DtqbmrH6uqJKk
5Z515o2DijgCUw+1x+p/UPAmx/3xRkXplhBCVJObj6tn8GqlnuRMerzjGlTXJUkZ
zSIeD9r9WvV9EBEi8Q/2Q9sHlwkYy8FntWpB7YRsT3ZHbf+Vzsjw4XFohjHI9suu
SJeB1/VXBDxkOVjz59+uK4YEEM1opmOgxKCPGnWozhhRNwaVyuCOeHllWWgZT7sU
5lqYFWw90fY6BSt6uSSR1YNOzm+2T9f1rem1nXrQd0tTbEt1OySkCvf15bb5PhFS
pnuHhOCFz6+pWphG8mNzYyHiD3b5CQ5FaQEzBcu2inumU1L3aRd1QL52fpfCEnPn
13laRzHelMJ5BqCJnsScBvsiuHo/SvrSYBVsXVwfYZ007Tdu6nXDB2WngqQfp4BZ
z/PT477bp7vlZQNjBSdO3hZ7TRHGESnQnuiLZDmDNX44W6llKLtwPq/pBC+eQKgY
DGH/dtE+CPCV0gAqba+9YUGBtUic7LsJYrN6xyAhaRLVUaD94lJ/+zQMajxt4Lwp
6yScwA9i8H+yutUfldaiTGlLQXpmkEkOXfgEOaIiNiMW2DlE7ICLq0P+xVe6drex
4vIiUilLr45VXEXXvQdLj6Y+l/KI4f09v+IsmAwqNr5xPGAZCbl4uhQPqKZ1zwJC
LeZTNkfPb74b0Mi02piUrLW1u2qBcwD7Xkg0lEMAZ3TcVfzRgZ/pR0ioHN1KQSGl
FulFE4P0YQ5hTPcQufWMsobvvQQx+4RLIAULaqOnrrIlpHSyNqwKMnPyNX2nQBiI
1vgIZQWblTeqGD7TIS7QSfhpmJNR0pwwjSocX0ox/jVHBktc9KqH7ouFsDLqV23P
SyQz6LwZFbLXXMvDWyw45g8P/SdxWpDxZx6KproWOIcUZ5Qo6CDvHwQQ/wZNRv9w
DAZlwVk3hHlq+FLwdwy0z6uYo99or499kDkRUPGFNwrxZkU+iSDXE2IsUmRC02sC
jTVeoRJeqnUPAHpsEmJEhNCU4rNQIzfwvcvCsdJ8Qkvs4tqSq8CIb/Ui1c8YYYpD
J8IyoxGe6yU1Xt/luFgzSXSXNd4HaH83FxME7Asy+Dj+vhLoliPQggqw8+xjfLEV
Usbu3T2j7fL5Pi9Ymb1R+z8WOaIuBg9R5dCKDa5Y2s1KPInXtPSlBPn8nv7lddpN
/gM88fGT2/HprBuS1TFZz4/S0SGEfH/5yU9+phHO3kpUEge22wL+5PKjEQ2wfviI
TYHhLwPPTQfAOpZXwCllN0xR0AxKIuYkTpjNQb89OWrAd3kR0mPdL0T6Ikuw0PqI
/I+hdJwmBLfrgXYHupogPTQti0RSES8W6IkIYVmrdOoBXX7REGZsgptKJG0IfR4I
Q/PNTpuUX9Bs7/PKCvjMadlJ0uHNqMp8AVflWuR/sEg5bwcjDldvaz81M433q1TB
EtEEqAu0JPo1bBZ3jMYgheJMHoep5Udd6SrKZ4NDa2h3yzV5AzCqRvO4hR9Bonag
a42PwyE6Te4Wwe8At/94AIyoOrPlwN8bct7J8s7i2TGL90E1CNCrBn5NsGbSnFXo
G7ZqlxGWt9VhQG7ub/o5fmt00fI76hP/+EGNoIt09w1qtv4LWSdib8dlSgpFnUjW
9bE3NJD7KSdx6zGmz8c5Zx7MfBZssZIf7vdge3C2V5Q+SGvkkieSVGHVfOU5TvPB
xqO7LF1LE6tfrZYQd7U1S8pbcj02Yu937YC9pooUZoU6q6CKeZpFH6QwWyTk1pxD
KvS6T2fPDRjEvhIRmbeLR4bWCtbe1cfxrl6aogBlivrAMYZLh7vFQqtnGa4zVCAy
QpoUXmys44IZtoVYT4yjm3PusYUWxZXGuYUPsi4Lu4IQnTXYokkUsHGWu30MUNPJ
VkLJrtE1vCvC0BPWrEJ/a4Dd9483AothoS84+eZ60HbWGCD58OCb62yB9h+3IaIM
7MtyVGfdT7mPkwQzoHETgpceLozvor0u+7yK6EOT47X5+/XHrruwtsjOdfVjnvVU
CVsn1bdkfV7GPZ18xdIYz8wCm/8l2yPMnASjlf6Q/GYgnUthZaTYxy3OtM1YMovy
DbCE5bQNbpyw85DryTilanEhSjoGPdWgxEyObfKAujXCWa9+wYnSCboyZEhV3ln9
ZkMtmY+7B7jccqM8PwBW0dmAZoMOD4f6Q+dAlnYqDGouwFurT7xHHBQXNLcGVWAE
eIIfSw6j0j2Yp6rY0IUqELmTnyy2wLVB30s7g2NlUI6d28o/5XGLBCJmx7vl4nnF
3xfCckyTDdTbwhKEM3YzBx0YeOST5OQe+qSOc6N4pllcPdACbbN7YVekVXc3l8/w
KUPJg7EWcM7uAu07iArHd2y/Sf4z8R78gzRwvJFLGGj0+Quuz5CpPFPFhouM+Inn
D2rLN23qYvY2LPPYbVRTfmRx2GMsg+x4Nx6SX8RYdShYAMULITcKLsHSrt/evrNB
MBgn22AoxbIjZ/fBTXxc2rV6HJKd2tcGZiV3ddIjecv8bxHuJLVzNqa0COIS6i9k
n5bWCtVNJyaTJXPaniEon+khWDESyu63nMeCDmrlKHWqZezy11m2x2JRbgHXMe8K
gPCH4W06Bl9zvy19L0/6EsbSLVQFmG1VY3z2HLRwW7ETRkdohj45IQJeUwOQ74WU
rmgDQjVm46hlEGmiWvnRBrAJU2tlr+HBMPwpiO94jXm4n2MqzjmGcmX0kVeoYp09
pTX6yno/5yaD5BMOM8FtTkSydCCHYXVmwKJm7GxSe4wLnzaUa1qOsCVLUvEsSO7R
eGj0br0zGiEPGuEOttCdrvvBAPrrg3OSpRST3dFIGKAXxVXY79WvbvfE1Emq/3Ni
1LZ5cBeOjS+JR+EFBYusHnrV8iAV7O8OlD/AfDqqVdSDsFY75uCcJfKnMGV7PpUu
QBFvIet3XTk/vAZxc6CfQulE/agwG/bUp69uz4mMauIFz+/kyiRQU/3jSkacpPn5
a0VdxvmAjqUd1u7/WKIg8G73mqOi1WBC+uV+kc/Pz5qTKGZWcwjdjTRwGp1MC0sm
vjZSlRSdnhEGjjHcKBtD3p8tCnjt5DntDGa+oul8icQR+q1PAdH+VURwhpAru+Ob
urDhkFOK5qhB6pRz5MQ1lCEro1u96su1qSKXyIhurtNy/aOi6JpowCcx+7qoW6dS
OhHmD2cIsP4qOvTGwBlDNHqsJESnKWIHB3ibGsKU1CcGmcSI6nvO1xvxhatriqhT
RhB5i5SGrCVf/yKBuf/QUbOT7mHlXHBFfSqrCrMmQrJJG18whgHlcJdC0BfB6t39
mAs2xCTEgdA3m3kr0q3X8yT0B4GJB3+GmhyCYlvo9tr2I9ZSQmSjD9c1saNyYR7D
r/jR9vWDZ8lWgSS4G6Hk38KcoB/wimMCV0oaeO1KxGV8zLDzEvVlg/i8q3/oKQwg
M865rPzSBtpRnNmXJ2q86p1enS+IrJheYIxkPm6nxdyaYruOuoPu5pLt8iNkA0KQ
qzBYt8p4JmRKEq71LYcoGW4pa9vr1plN75SjPKP07IXoFpb+rf9UZrY1izyH7s6z
w8v1qMx5rjKS43esEIS7ApMr9rdkZgBR3hg6MGMjRc9uoiYuzxwUGoHAcyU0SDlB
XDcSZY1VtRbxiz55daLxBNigdEtZE5gyZ3YGXU/lEJFEWK3S32AwNuMU/eznlZe5
0tab2ydzeOYSi0GJOMI/TXB2Z3uKX39vRwBDlX4WY0xzZuzZxD9MppboP6SBVaOT
j/Y3XZpsQenfmbZXeGWnIR6w/eKMZhfMZxmGwgCKn/9jgiSsozzpz4yS8uOe3SRX
OX0P2KOCw67I3R/487+elUdJ+88weyrNYRNjkBTg8WYt6j6LoqFYXe1mw96GdeuJ
fIniMYgzJVAPCPDHcjxmzVS9KlhkPsNGrj+yCO+6pO19Cyvmba5ZKnZED8bTGhZF
nH3KZ/AajwRbeOcTpURagZJo2qiJegPtiiGbpEusGkNcmMgQFDx//zj4Xsvi/GcV
7I5th19OmuCFixJROIvL9KkJ3hec9KD+ZL2IoNkiukcbUhLOND2K4wVkD8miTjHC
nhUFu4LxzgBTfx8M/zVzK4e4FSpUJezGkLftol1otHjwPKT8Gj53RaiHTjYo1SC/
JXsESfJhGC5c4xpCm+bicfuT6wpF6HFYksbDWvMd4E+IOF2WABxiUMciENBfUAZf
TVC0oCEb2wcyetFO4aEk62FuAek/crflWh9xGGVOYy+Ai18nuODEflsNhYWplfrY
12wHv9JjCqMZm+G4o5aVfhb9PC6+0aNx+ZrxtnPheLZqjtIeBaQrA+OZOiqx5b/a
FX1oy3bWgICZ1P4Wcc24gL7hDvZHUDZ3JeIoV3yoogIJb1kJ7yRCS16WAbJYz8sm
bgIYZlWvBZjLxz/7CG0sE7Dk0tVwFbWGAgGyclzOsjWHcdctxy+tZwKomGOqoU0j
93AyQCeXMAjg8A8/OFDmQsaND/nTCBHJWEPZbC214ZPbkBeme7NhW6HGZsmLp/jR
iIas7ej31GqWLdHsN0mSvpezSg4ObRqG4wlMrW6EcDIhAZhUkRYYBvE0Ahobr9lY
NPhFrbFyRIMKLX3mD5VdXZsPtvobi5kiXl4XGqQIpZtj8l2A8lcsjLIW2UjT7I1I
/ozI0EIMuNzfTbCNMp7eH9Cj/hNr0NGJo2HMl5P+m++sVWfK51sUBEZhxTSm/0KC
yKz8y4di6KkEkSK7lOo/POvE8MBBAl5K9NCwyijH5UulEqD8Q9MqOFPdTzEdLPCS
VqmSwxh3d/KUwbOOZswon9PSMdBuGMMecH2ZR9Sho7OKb+xrbAXFIhTdaWgSZOPq
RV3vawICKVV6zRBJaGUY0u+ReXgOj58FzrwCvb2jpImfnvlAgkmCub9dnBwRbOXK
7a3BIwStpz0Qdvc5RwKP0pTZyTDGhBpFYpz/m9v/7HoWnyVU5tmkIEIIvlLFwT+6
ZPCaYnobE2fn/4SkA8FRs8gwNhgg0uEcIPSI0g4B3L4C6GiD/1lmHHf7ccypIDax
/mSYhZYavrs6utZZOJdclTHiCM5AUwKcV8eMmlJeP/GdqTP0MoQDHmuFiJC+q9jM
Onia4r2UilRLBTZCL2w/JG95qyksTUJHPMnOz0NdM0VMbvmPKQhW/0sAqwknzz9w
lHAgaqhgs/KmEV0jMLvyui8wNvRT19i+u3b+Ku1EsPq41PhTXePZYZ/vw/ktoUla
WNdNce7U+Npr1gHgiX2SssHzjGfc38mRGW4dB9LSlEnJBbwUNb/wNRs+hiIp6DG+
YSgcDCax/ASLPA/V22McWfvLZ4c68t57W8UsRTDPAa/v4E0Orel90xnhdnGnsNYf
Lohp+F40zZzk9eAqUDYlp3QEMxN9QiYx9tkzDL3pPMDHQFapOcoUIGi0Tub3N/0z
WVkRfI9Qwm/74dnoU0fnYxCklu/+1lWfqPARiZimv+waRQt7kyoOhhs2Xrp2fmJg
LSxO8UjOXWOw50qHlZLM9JDdUe/wpp+fp1y7tHHES65lCDgpZlpUF3le41DMoceS
8xS/Pqkob99kF7xpM1NrMe3z0y41HTdDSVnSoVn1Z0vzUGTt7tNh9l5M/YnuWCpt
iVtqGrsQN5G8kBXWO1PJB44oTGQlX5dprI1wwJ9bs6/FAoRecTHP1iWzI5ojqgQg
L+HVJEbyWhitNGqVvlq6bAOC4WVDkwXHVuPmbmUQmS9sCTu2oU6vUyvWfcXeA295
vCZLphmW4jnBMAwi4+DSqyCfSMW5sX5R5ohjwAOjOdKfW6uWzK3UCZuWca4AtKLh
c7zsL31vsn7AqjjSLnH1z15EBWOwSpdSid52831ycY94vyScqsfgaeJ9tv1eGVAf
k0fU3wFAZ2AUudcrdXzcuO9KR342QjcDgzgdUo+nWzmMSeDgEEf2T1scR1mNnCSG
xwP2ZLqtQenWU0VkibOD9K5lHN8vsqZiF06fH0u19DW+rttWFC7XxbVWzT5vTjyQ
cQhi7hVdq04pF1N+D5tTSBNUC1G/dxALKniw/MMDVK2en2N7ROYrr1hDsgj6Ymp0
sy2F1GgkrBNiweoX+iHfFhuefF3CfzGEnru9mmoE2/GjyQqjggonDlsM5AZo1zS0
xG9G1K7afpABtQeJOsNJZWqEK2552TJf13B2OutiRZxRH5yTok/MkdyvzvWkHFXt
udJNuZvqqHR8grmbFW75clzG8LnjAubz5pcErt6ECBsq6GfY7X1+ZUv40LBRYxhh
fyQENcrQj5soxigKlfECl6Xz5DjqfQjYTHZKYruoSQjkL2MGmLGTom65qExM+9i/
it/PwU72yfgnJJYrV+uQ1gO9j/6qP5HXuIBv8pBZm1MqVxYQiBJtcug0gC3N38kt
W0rBKDBTP/AvJsR/vDMsUlUTsHZdfhhDc0dvfruh+jT7NZbuWw/Y5G5/TMxMxSmE
lVC7Wv5PdT2Vw/Hb7shipYfIxR6H42Qlw70MMEtGCv+4joRgTApifsQCoavQfheL
yXJb0fQdkt+ZPxj1TbBvyWejoqfcSbLMOOGmPOtu14sGLGRK0Raz6jRDcvhgZPvS
SOteb9WlMSZeWjS0+XOOyL4aqDa6PsZIpD9m9hv0LT/62TZ/fyfYMx6dqtQYVT/5
2lcsNJPD+h45ACDwq0VKwqiFyaIhwEfYZceYyznnigOkTMThzBkNMFWS/QUaABNQ
I6D6szCMN/B/wukCzS1JUr0N3ny9DdanvCMn0wH6vc0a1Z4JRErMvEsA/9azTWbj
ANWyp6auTHyJFC6QL3gws4IhEyn4Zbsr0OhKWa6vognOfVcj1SLjVVjuRf7fUC1L
4fyvqMLJnY2Kz9H5gBJ1XVMZXl2K7C7O0TpafN/KN0OcfAEzogjQ0/AUTs7akhpU
5r+YcDHZVlACdjTorDPcNyLhbWjlOX39lYHFQxLAgvqjQVhPjTetwifV8TGbRqh6
W2UlOS2+HrGSqBNS1ozOLl5ofwY+oOumysBGiUImx3KwhNJpftG5i533SKu0PsiO
FbsKxP43M0hPZ54imAx/hUTla374y7pHWcAsV3Q0C5Vqx/hqAA8wxyyFh9C76GTm
G2fnCatLHS6/uWmUbAKtnCz5UYxT+SrmSxhoI07nsPSzxRTkAoj9dy10D6aXtXul
X01mNN307MH7NRQfZjEabicOGIHrVblFzOhXa/nksxRw7C+PeuiaL8VdAR0lq6GQ
7iKJ0JsW8lW2rB5/kMQeLsHvYnxPRhuIJRYO/8VRlDr2Ur4AyLHIjo14ex/hWKi6
8zsKP7bOAdT2C6MJRkXk/57F3XBMcnTWplC45/oiVPovkMvW0ekiRXVOK9PsUyX0
W6Utxo0JneDUhiU8rafow5X61x6m9f2tC2R4u6GFHs6tUb4OU2ECFVHiS1QlGwfd
B1bi81grG3pCe8C19tPkq02sMHEH3eyJWOecf8DUPObCuRP1fJCmqVlyYmC3WKEp
h533p8HlmbYlZbxKzevZ96tIALlronAx5I+uzrvuH/HkpCYQd4GCpjxEniWXgxzB
5TU1J8i/lu4+P4zKXOqA15o39Ym4/ofPlNzW3RRfrG6klm8NtOG1LXmdNLQZybz5
+n/pcpUxfGH2NAjAks0TC6mUttjWS2Ubh9VSSrnSq8pFCYpEdiMkZ4Bd8+6kpIUp
+BXW88MNe5n6In3wxxAqbBfIzcxQbXm6Im/6D80PjlP2vy+NrlAjzBKXvXB8HSEE
9y55dfE2YOR0pkUBoLZ876KYxN9uc6apADYg3EbGC7AdVVX+e7QxjV2UtBzB86ZE
4bZbT3D3b+X25wpN/NZfckgpCyHPnKb/WfhnFfoBMJ6+Y/XbSg6CrdmexY5As8q2
KdZAOf3kZaxeskHwNASJZpaI2nzQcpNOPwhGXbpdmq0KApHfLUfpuKIXZxWEwiyv
X1+6x/VBf8q9S80p9gc60OFtMZ48bxqooORlspCavFWWl10QvMuOIPSPgfHlQI+E
3KPaIH8yce2hqgpR9H7WawyL5diC+XIwe6cEr6ExWebSvMAOc4w4NDNor1VMvY1X
lF+LnoUmyaZpwPPe38BmTQZzeTUCZahH37nLW7wdJV+mNbcBpjRZnjgi0yNcijq2
R3VYwfOzfIzVx+3QiIIDepaFqjr93cHdfMPEcXFWguAT1VqIIubJwzOb5td+F5BZ
sANLqKwvMUZ+AvkF1IoomSU1G+1UYG9L8xxWpeOCOauGHzjc2ZO3dFk63Gp1F8ns
85UIRljPcj6IQbF/iurWg53K3qReya28sVsNyXEHUslo0qiicmCVxlKPWVQfl6Sd
ECj0XfFVcv/JUk710Jv+PowWdwgV0jLcixyTwW6XQpUp34gSulDNh1lL434Zlw5d
+WVEFRfo3Umr8FZyCXwLNxTSL/WGFdjKXUxSLesrYatDHdFJK9jom/aDbuQdbqxd
X75tPIFNyYGAhb4uXUtEyuWglFaBtKGICz3fjEtJR75Cv7MhFnzf9nZTuNotny86
+hRHydom69o+2ZyqZJxMJ4ozZ6F80xdzNNYY/EFB9CvxsQK2EqBLfTr0+rEbEZNv
yqAXlzEzI1VYi1YRFpGSgLubPkvRXMvsrsrt44OqLdycGCrppWz1n4iknpgKeF40
TBOqjysiHbl37zCJ7CJKXiagHDyxlX7w0vJ9Bl/yGeDLuVZiUhXQ8M8Ca6w48EDK
wwzlXlVMUcTNjFEaMTapjK+U9E6DwMzhPfCSicZ2cpC6VGaJSkH8l2M5I+J2mAG0
eQLm23wj2oVNNRvyHagW3JHlHwLc/VG9C78yv/qUBPH6X+bhNZquTGsBVpdN7A61
81toj988erMcOnyKHRKyA+i5DHlvhMZUP+soPrOpecdqXm7DiYLSU3HYnZL0y5Et
03QDm17bmwlDWfSSc4J+N4JptUgpcvoB4ddOqAIpDAX85z0RIZa7WFXPNz/RplvU
YjsoDGNuwNi/id0C5govIfO0ekfWDZI95vEyu45rO6rcIDq9ubXEIBrJK5pj61Zl
k8s1H/Di8ait2iii8plf4c8N05jYa8FWB70CQ35Ce6TQZHCXxRt9YESb0VgskAI6
UmY5ElnGHoCw5Krm4x3ZMOdV2XazY38NAu/EkdMGr67pEO/6g7evV6ch9o+vTIM0
R1qarMoBprNAhiXL6GJKWh+QMg4M8MerKir2CZn/NPoitL5L/BOIQLyQsbzEUc1S
+aI6hVhbT/bo5HfhLqJFLlny5rlBOK6iETQfzwgJ7CuXI7lxTweaYiNI7id+Sa4x
SSCXoHIaXPQl2tZVzIPPDU8Q/ExAZsF4pq5gity/PkNUD8H+OQEsD7jd24puh7z/
+VqLUPPOdYNHs7FeVZ8J3dLJu0NBDalCHw3CBL6Cl/eFfb7hea3EO7tULG+xC5Me
Aasck5sQcfSOTBmPphSDuylPnD09li+Vaynlid3WGqvwkstUM7qhPWFXAsXKp3t7
0OzPiik9l+jb9Ir3pqjphFfyvJsriNyZicqGBMri1FBz2kFnTYewlvmeFt5L7dyS
xuDsfosQ1PLfUXPpRupTZYa/zYJ0IEXW24cK5oqaDkEoF5bdVPTRau0oGYKxPDNq
ZtaDM9Pb6lpj16bfDTDWFRaXo0hWhoVqGy3x37imRvx5FuQsrs70UJz0K4xhx2/x
IA0NtNHD8mCrkdvtqzL0+I08N5fMWvELoscCogGw3IfXAZcjBfkjRbtkWGKZUtTr
jr5pWjzI2L2timsI6LrSbzHJwwhJ6BbrI5SXw/r5fqeqe38yNuiCd8m6fblrUE4Y
3Hb2bi4YuGxi3hkKnYgev+rqpgc07OfmjRPAR9WFnWj6PqAYFcHFvFjHn48sAQib
aU3T7UwpUszXUppxZO+SeUoliSAsYuDiJYcLjoC6SV232F1DYznGL8pmXQ1Qqv0n
PRDj9x619LH5fvXC0VDDaaKUacI+iCGQrhkD6SSsqNRiY9wyGBqzXPgpVp1AQYvy
91CGUnPPb4KsMrzKz/NkdF4tJSkuZ5cxOqddmO2mlBVjyC4wIVGitNvq7nl64mnv
CkfpnB6u09GOGtbY95+Cjq1Y1A0vSwljyTIgjBH4NYtPfWoanoSqU//6Z+r7aC+1
zzNqyBMYepC8Gdl3L+jRY35+HJFDAkwX+N6Ctyf2VC4Vim4Gs3D0OcPjE/ouJCm0
FHC1UPEL/CpsvfYfuaIxUtC5xuhYtFIMnVkJiX+JrMEIFZyH6UETovJWs795HZ1p
pa16wMxW8g9/hj6HurGI8kWg5dK9v5Q+e+L/wk9QcFTk2i4+L1zQ5jE9GKjUeDtz
zowd2Nxv9r4pL73QQJIeorhh3aIZLcRbIKuhTFUkkvPk3n5Or+qQJOUliAPWJ2Z6
cvDAZNqWRo4Z0pwxs+mr0r89B0pJeQRJpVq3lu+VpgMkEhBlYQLsL9wVHftTzh/e
EAnRKIyLO/mshptfD31XjUd6pUGw79QctlMlQcHdlQPZKj2GXFExailIDrXmMSnS
ScElC691ncvQHtI/ZpoHTi41KpX+CKGOZXTeQvjsLMHDS/iUHoOvzvouw8cSbDyI
QSMAVTM1J3f3PXC7KsEqK5HQXTC45YddaQ6J8O2yO87hbyVPm2b4yHAxngYG8CCI
gqNvDTWz8Iz0PjPCbX1PcUzhdu/RChpGxjaQDA55axXfBlunE3d7E5j/mGomnXDK
xQehEPzQlVxsq4xTiemWAy+zFwMfWYtqpHzUFYlVN1F7hSTEB38hsTJlaco2n/F2
Jkxrv25LQGQMWQa4JZBAQSIdqlhTFyaW9u6jlUGqqAXolKlzEbngtDIMkTfZDLRp
HGTng/Kki/ndfP3eCyIQReB89lXMGZ84xbps7STA8PvQV+WJGsMi5Oz7z63EguxM
WQ/p5lrWkZWeQhmPvXQ1YsH8RPjS9j4n5N7ZnxfQoY3DNZ42dji1NYyUqwHuBSZY
wgBn/MIqyfLl4/RiyZXxU4FJRv5Qp+Q9mYTL7Dh7eO/W037jwk+4S+Mb0rQYWdNI
mGfM4JlvTyomObq5Jkfy6BwY4GZkEbGJuka0+WBDUHcvPINGM5rgVvXvUEbNZBX/
CnOJ027Ft0rF897vSg5M4crX5S9Ra90eZf3F6yIpE169zafA8tBkYcBKU2nxInf1
oFqug7A+J18SJ6Plq0ZAKpRm730dd9v2Z609HqzrGkd9RPU51fEpN5RnNfUvPRdn
OxlHtD1Hwov47UkMSiYJGt4oO/GzvY0L/2rOh5j+NPD6gRc9bhYVEuap289B2Vgo
CiIYQbdU4/EVQvzuDpUcmyTb0sBd3VJACOD28AtU5kHktW5ge/h5cyCAgNLvdlPz
+pyov3kiWgQZsGcCPK//FAzKMQ4GHmoFflL+ICm+4oBu4mM+LKrJMSn4kttdvU7T
lShznM+R/rQSkW3auSHZmGFcyY8ChvvviSJKAyyjTpBk067HPkvzWqJ2Ued/dnLv
gFVCRHRNcrndcbwt5ycWP4pc6VKczV3TuXCRl5YTxcGGhVabfQqwY9DwMr0p9bba
lGnPQesyLd6SKDVa61+9oMlHnVNyLe8aLDrOWEHVlOWrCFYahZsEHHNIzaQ3nIRY
eGsfeN1OY8fWlYMYlFBqkRbO7598mWLAhQT0qYdSJgl6H5fbrvCaVI4PwSL1/ljE
2G3V6z9F95ixYwmc4+tGBhSyWm/5Gtvz3YmY0vceIEpwjOjoU9FXeHJQhunKzXiB
d/eMsho9bqt8l4ATv0SlrRbvkj6uF5fWGpM7NTG/AFHF+hEAWx53iX6cAiZqatEe
Jt6LPphLqXFUMoy3+G3oCNXkYOttOhBZRjqSM4Mz5EE9XjkETHpftXGi1dBqTfMF
WgqWVB3/NoM5SgmU4NmmOHZvatHL03az5hYqW9QEQho98QtnbTeK0+BvBrUwFujk
GAoZr2O6OKIurbiX98tdLcMRtP4sJALkRSQ5JvvGeuD9Fi2H2hZAi7k0L+yp8/W3
Z88X1VUSwVnvZVVueG5B6nzUfcIwUgcaIjmQWvmcCFs7eJxFiBsl93Ss+LENm4zc
3k3EPJ4WzRrMT5bOZKaKrcQtJioIbPYaX+LGqNcKuWhjvZHJ4c9WFqQ0nTeqsRKt
XTP2DwUPDPVk4EXHr7rSwAVr2NJZmrhtwGq3GSHJY96Q/3VlFcxV8/8fTr5E1Nc0
ZT2krRfuC+Qf2zSoVpH0H0skFUGD2rrPWM/VmEnUEpoDYTrc0KK6XU+pzg+5Jd0X
BBqPoPvsYhMFjmGWjZbR1Y5EqrZflKQMXpDYvEV+v3yQ2RJj//2cJ9R/hRW8Az/r
hyRiGLutEyXDp0FG638XpzgJ5tfIIwSE9LYsw2hQlOGPQgxgVBqqrKa4O0NZVlWR
T+z8O/51ETfX2yO9DSZBFOHtE94ZA0EZSRV7HsiSa1lrdKSTATvHkEUmUpGZqIoK
zUwr01f1fhnukHK9Nnq5C9JmWoCOrMGBqCri64j52aUiryuedRsbT4szchY5dlvB
vHB087HDZiEH2Wjm+HPMtFcc6U6kwV8Ud0146GQkJToOl+/bk9A8AoLf2HRXnZag
mTai+cRgZgDugXK5jfaaqiwJxM5bkfql0aJg6APIMKlYcZYd8C3lA/8EULOIbB8S
p2j1Qjgdfkvgov3/O9ljJxw0G+wlwYwlkWxosZwbZCdRAJ01T6T66TYixJ4gsPnK
icyex8JeyvtTXSU9IKil2PuakR9/DN6zz4uDvqb1pSniO/WQFiLpOBxrC6yLHb6l
U0zrFIefg1v00SiSA9iimyBEC6uLOv6CPabxHVGcuEb0tAwkOWH0zoGYWvfBLLQZ
vS86lTUcw1FobO1NfZjo+z+oOm7Q+EAlBwSOWzHVouWYp2FLALiFkemfRgq83rAJ
FqFcFodCFJYMu36UbGsK9nypJC2+lcbfgZOjBqU5wiGrmXElcIHzxGDG0sNHAjvV
LmBFSDAVTE3+b9D2kP78c5W3MVVrEHEGzY6SbujzppVn/0jfM9aOzc3h3bwxrXOo
o+jbqkyNLKMsnl1m+AW3sYjmekVs/0MlF5wygsQBpRhNdVtZv/Bq4UGmkp7Yy2hn
iH0iH1AG8wzCpv2lVcjZsnYrNWL0e7xNSoV8kQL3yrv28aXaQgeKPVbs4dxekJC/
tsIuLfrSDWeRkkxfP8/pOjgBFN3w/t0wiPrJBL5EhSTE2a8Ez6mwZbVDUjCKSbnO
6pNiFKAWWcV7muTF6mip2i9XYiP8cGFqSMY8lVRQGeCM8sFK5ecxwJHv22N2beIQ
YDXLxtJD5pZCqCw+lXDssiUsAguZZVcibj3pBbMKBdR7dyYcdiyitFIbZ3hB3AWh
kqo268aAYP+w2qzvravQ1ONkUl9blueStZ2Brjre91gQy7pK9YmuEc9aeYHogNJ8
Z4ecrlqUdQYh2WmVbuxHrAxQQQyjN3YN6Cz9fyalkbVSX0aYWJmlLW+RapkNiZWo
CIF886inBxCx4BGAtwpb003yaihXVYnwBcyvQIdHRD4DkO6/HapcLgZg17FzInOZ
1Wh+EjBqhRa9ZRukMjLs7PVhby24XcIypJXPm374pXFKuUKRX9dbq5TgIvMm2CC9
aFih/qKNxAnHcNI2+eoPn9SSpSONQoi+M6mxN/Ho7TBqs5uoR+nxrGluUfhMQYmm
nq2R8SEVbkYjwMBp54rL+4lveRcqNZDgPG4alctzXpTEqcYJdtK3JWjqDXTtMsHk
VivfWFYBz1hGcXHgDaEEQXkRKkUDJEeKEy5xtgIwXY2787jSZDsJiXcmDzaS61DE
u6rFAAPGj2MqSn4aq/IscXGbLIIDdD5cQSStKQStl/fzE9LMO6hEEL9xg7J2Kf4Y
rTYpaj850rDj5PTrszD0sXCEunVqEE3TwVdswqmCtTt/HJUEET+b0+p9rvcyIDUJ
43u2ZjjOBbMlY/b0noR8C8jbwF5adiMcyIUARHfDXherJ8rBCEra2HPoHDdnX0Pi
yHYeWTvuopWEYxMyiZJacs8Fkf/1Ozd6w7pWEAJ4DRCtggCZnJh4CuBEafbdy0Pl
Ru23T/TsZQC/6ZCN4xMOb1pFBke26xmBafGUxlLSyVQspy1Q9YDnGDcXozAocUXf
V7KkA/vJaY11wOnklOCcvZzuej+PVOTlPXG6c1grDaSyfRltsgHnNq8rr0EfF9+I
koavz3nTxDgtbyLN6qouS5aoEMRJlpA/1UlGyoCPsB4RN3fDXaEktO6oYZVCHatq
8PEmV/HYhNj9muDRBAtAEwVxhH3bhVWySpNPQX4vlvUK32Fu1PqjzaAFZtPI9dhL
DV19zurupIMt6XTgShCOQjhawsBPt7g68HSVksiXlbF3ZTG32W2EZsgvjdUEK8Z+
i1/N7G1yCKP1HKfZJTa5+mqxZIhsIN6Y3PdXe1f/7VErFVwOE7e4BP46qVlrtIEn
HmmEsJF8P8rqrQvtU8qKXSdwCEz/Eq/RLnduQ2lmBIK1LwJI5F8LondXhKAZfQhE
49jMYZHO82Ytnqnp1TVk2ikHkbj5fIXDni24B2lsyz5rJ/UaCReoGBxV+iUR6lb3
vAWB+SWd8EFcJUNv5Pk2mHUGHuIl+RrJblKG8cCdE9Etk+7R7P5eI4+t4a1ziRHQ
04LZyKLZyAbKagns0H3QEshBr8n6nrF/UDEHEfEKyzuEDO+PzH1yxGYwl6rJD3Ej
bsObWhHp2I2FQ+3Rr+xqVsZR5eIQZPFGGAzD8K2tt/sJ98VARfpuk0H2i+Yghi72
MXf8gMO60OnO5tY4wv2AGixmLiZjQ5wdKEqiSOiQ1ZipS00Vy8NyS8co8UZT4l9G
K+IbA67MhqI/8+RoIHc3IjUE0fHWUOWDcGTL0kQBtjAXm4fVc2W/OOu/q/cKgHTY
36sAxWRrCSAxJ4QNlM0CA0NehPn+ojJBJY56jqYjHAnKaR+wNm+tOtOYVYGisxVc
ywlHlB3Sisry8t5kveUvioJrVzpXFJbqVDF8esrn1tyelAM/9JTKfe23q9QCyMqo
U9zSFgUiWPexLLfT9n5GSSYTkigs9y1Ps2yEUdLJlZRTEnh1ohKcdeLEU0AAvJPu
qtBt8/pzuhaxH801ukTyO01UjhJl3I49rAKPi/OYaNd6GBFcBQRFbBZlRQ1Gela2
PRRNvjnaDr4qD1QRqXgpHbTZ+Sl4rIPwckX4LCCaJoKVZ95KURVmqWII8lyy5N+w
14vANSYezCGcEje+DHNcWf0O8oSPcCSA0jUapREgYz9jjim0TEPi/X+A9l1EbDQf
p4Pilickmt4dfJtRDPmrTmTltcfyfU3L5gqVlqyG8jxdEuUg0zbsEkKqp8TUUnIZ
FviiPPCq3m1jYArnpGCDxqWxBoEE8pcpyg6+dfQduLhs3HhznoLpEMw/Bogopm5/
HkVZT2a717D3wk+JmOum7P+shr/sBdN7B2mYjw/v2rUs3Fl6a8eKJv8Dq/EmXWL3
hTh7+4OhayhwbklMAvdtJUAM1axsY8uounonIc4yWyUFfMNJBD0UvQYGIaKbprfF
DG7LceWHGmDCCSGVv+eY1jJPZVW4/Ky0PhvuCXa0T0qHIeZmv8HQdDSNFg8bppCp
B7osZmytV4d3KjPFUyv4Dlr0ORrkJ35yBwqm7rv7zfvYfN6ANnGBygRRdN5G17FT
HgomGXZ4/MXpRYRkXR6oz2vIiDNZ/fNLkyWgOz+facmqe9m7zMjyJ90VEQwDkZQQ
ullt+0fdxT4PxZx54ZM+XxkVVBFmNd7U0oIVwnz467LLK3/DEoNAi745VvVmkOcm
CKTJo3/y6U8uJ5vHkLvJRag/Tb+tfX7CJWj0UO+f4JdGemu9NsjUkdruArETjMqK
LZxekH6TLXKmiMiGRB1eudkvyuEoTYluY6NFeck9A6hFR5cF8j9P8zUyLa+p5Oni
zLh6jxfhNM60NlFuXdIkUWTqAIruyqDCUDl0pjU9grGBljDXguUXGZuWIfEQlrO6
X4ixjUXYhxLlKmj4d0LtF8HzE7JrNCXXr5mP2EaW+tgLOnsEKWuEP5moLxrQk2aw
uylTwc2rRGiLQFuE0r1u8vOfwsTTeXx5b0yxfp5bLzpw3eqbZ11bL19aBajF6HOl
4iaeZ/Kma9SOj5dQh4KnHsGv+Ag4xiHqc6sGrYRUoRrKIGP9s5Z8STop0ldcpIYI
MydgFhOlGRJdTY8JGtbYNVt5X3dJzap61hCPS3tc310eDAKsM+tEdD94AyhmGsgy
HgeJKPctHiBv+IYB4i0FrjTSLWdQJkQXoy2pPvC94qnFWGBAkPFnQWOzxTzhq2K7
rQXD+hoh4gWRag2JP9oBSfE96zLDwusSKT7KrQnsCyonqTSS3Nm5jwdSRD3HR6Iy
v/u4uiL//soKXmSM9yQj5pUFazzQLBsQXS+HMkvgvjsFm0opmylgWfjkbZeUjRot
4AuDlTUv0O+MJ43khBIUuGBaieoukw47ju6K6m7lyQQVtJo74JuGJp/hLePnWvcj
iC3kdwnkOpgSgxqDI8Ujsp1DsOOfjj7Rd4WprnOPhmMRMKsgIOPHOgDyiBWYkV8W
HUY79F4nG6VJ+Ewj5UwGggNvapEHgQhu7NjDXglJtFL9AS2/PLqWIT6yFqUT12+x
2nNSS2MVQyCd45SsR0ZAJWxLxek9zHUDrGcQod8H7Q+eeBJFt2Sleo9DDvdZ+/id
7qSgaPknfIrfiJyMcmMkjiuTygT/QOvQzI7RvjfDCcse4jHjclKq8OBUgMjNuxBK
HcSCKn3BghyeCEQrqg52DGFTp85fIzrrNrMxxhtTfGDTokpdRfAIWQ7ylApOGTfi
gYZwPZeUP3yjz4dF9QQbsvXJzSSoIVg1ZwE7F5s2JNcVewYzX/IxhsqUlfbQRtqO
OCjmSiZr5RdvKkzDmKfPlnl9NKC5iA0I7j5K+K5i95zySViJNOREfIomnUjrwx7X
Ffv5Jwp3Dcgo71/EzU/FRRPRkza6xbjs2wvw4ckbt3GvfCw8vHmUhs1ziDTlbwMJ
coWAAgC9IZfHfY25RAD/gnSu2edgDCwaJcL6KuRD3Uwzkf9oUEKUGWsYzd5RqUy0
TXXeAN27acLKAOYRLZOBqxRvVId681ZUZEr/h7pr7Q0o2aicYBCLk1FY9SKwXG3L
8BVKJkazVQTrRrdze6eiuiRKfNnNiJDn48Mn7AbqQaYK74PZ9NfkQol9UZZJqQtI
h4VGF1xklnYps556gTqJ4EiKkx1YSgjXX55sGrxoMchGffTkIuebM3vTE+zIEC3n
Yq8UrlGiU3mmEt65ByGd9LpUZ3+F1Mkjp7wIh+z5gCueN59dlgvkpAcofAayHNT2
yuA025UsFf9DtxZD67ukFNWahPBvQG4yrKsii7EtXQLKQdLwrnrZgXw/QG5FcGbk
8zRv4N2WSahvOqOeQn/Nn8wtRXDu+foG9YrV6X9C1nxIn8ibdNO24hIM0YLXeXzM
GYlwzp6kmF7PP66mDxPE9rS8fcc6ofInymViPwhqktEg9k3BmUIAsK+gCLj2BToj
/xRxC82btKPwNbetx6uEdTSJulispHs2Bus3xykseOXtZOH4GOAF0oR+shanEA6l
kfPclxQ6ItOG29XpB7woS8gwXNXxm5G6rbK8cVMZ4HHYZuPSdxr0+iCijUhDARNE
hiDtHoJ+gwz4jRE7F/U0mNeTYCxHlKhk1QqB/12xrWkuyKwqWKrazpszr7PA004Y
B9JflhKRM2GaneVFoAWRLb7OiQG9zBXZBcovW+OzdPInTBv7HEm7VtEznLntZpF9
IIxzxA0ZbHlTSm9PFq15q07YFje/PevWSAXOdktkLNZzbtVGT5EaB/gf9pEC2GnP
N1ax0n4r9peiQ2Tzb4cRzV0RnW/ouP2NXjb/ehFHMJlnVUL9qMa+eER1TpCXLfV+
F02+lnJRkCSknZ+fSbX8QowcPXPCW66yzdIVXVBOSy7va9yeqzJcLVTtxUACbcO0
YRWcbLE9E3ie+E/oS7VqIzNDTZIsdZ7r2UAq6JxA6ueyD5ha/7zfh1Kh/qHUVV/Y
gkgy1NKW4EoyWzzJqzCnow8MTrQ5U5gxmzCSEDxOC63Vhg2AzGo4XqPO+JowU4E5
tKB3ZsT0bBZk8RB/nIw2RCd8iR1S8yJfmjWNlViFDDSuHyTaHZ8NHpSIrVqc2MfB
ASo+6HT0blTupICVrsRgl0cnRs4ZMkQWCA9SuJdyJSS3bq05vyWLVqG+vDdN+fNj
iVtKNk3yig3qQaKrrosOVmZz0gbZKumemYoAez6ReXFmS/+GDljFvZ6vmaE0Bd5a
b+ItQHD20/dWwuPuaVorWOVukmPR6Mgjn6zi+s9APYTP0roWk6EYOq4Sr8NIlRKk
DY4ulTz9BVD7LeUm2EGpYgkLvGuhiWr7nnZVNUzowVZkbTHfe2paevjYfixxMrJe
kJDfwByfF3hxlRWDEQ+KaH3Y3x1sHqmUgH5HnlQ/barPxM15d2jL5B0URxspvkuy
Wl5H2YJ7Sa/zGroOW3JLUxgkIzcKDqemreuEtvl8vte9dNv/QSD3k3mW/mG8Cjp4
8R1ximOenYsnXwdwZKbR7TnCcRBpX4Vp6CxmOy11ijJrRhaMacMVMWaNQP8h3xeG
jyCpMU5VWfSYQa3lnWFqW0I1Xx3dlp+iW6iGlExEPvfTWnheTPvaYmhSlAmf8fxF
QrkTJmD0FMN09cDIr9+f+pYu8+3qwrAvR0d2GkNuBI2AFm2CunoMLwHORKGFfmik
dUsO/HQ3eU6YXhx0tfzLSEtXY/rnQI5vri1Hi4Cm4WLZxE1Kh7tO760z851aH2PI
j+weQzgDfHzoDB2mK3MSaJgc7mUKr2Cy3sk29/1E4qrIynS3kcJMiYhKG70ou+fj
hrZ5RtSQK8xOxysPy1LM+/rjAtuMq/L0vf3e7tCWNxAlplr00nGksqHPk6ZGwqWs
8FKi2XglWJwUuVFiSxqpy3A8SCv/GiuX4Dg/w2j5f2q8XNWNpTEPFt+9vWz5apCN
rGjlkhXgkThp1zEzs3oMRCgzEy+dulLzRuEDLN2Y6PnQchCRdzKQvVffiRirQbrG
EiVD+cgLx6y4C5xgJBJAp+9KT0jYSHw7H8cENKkjPf4bAa5twKEzt9XBseOnG1oo
AAkET79NvboP7Fu9ou9l6FZ6YoSss8b0toRtyQgKr/EzJzmZMTrfwrEEXFq5jfjH
ma8ZgPUFJPniqNaSHAHtQf4IRMrvxc7IpJWqtsIPAqp+K+4xVlafOshSrNMlQVCg
qmyHUHBTBv7xhOZFR2bmLgvUWayw6606aYGcYrM5F9Veve8FV9IMG9EJQFLmj/lR
zJSRBnnJTaTppeMWhpb4f6yzqYY/sP8BZMGtm85zvvrrnXMgYUeJVVmTlSuuu2q7
2ojdRUNlnoUS88MPLN73kXxbMnmundkcjvDU12tn/UyuSQAy4Wh62FKs2lHSdqzt
oVVJT9rsVmeHjs3W9AnxxHFZxWIpsGTvZ5c5q0V9qw0aCkUVy//qjl/grHj0rZ+g
ZmYSE8QQMi6rL+6EeS50rP2La0WjovAzU1TOmyJenxIe5J2TO7HzAB6kPx2LtBlo
T0SXrjmht9Hck55byOYRxFknN3G5l5vl5bzDJLozmVfz/R7DUp+n42Zgk9JwmVEi
IRYjKKURV7+R5T+MX3PKEDDVrqKTke0MS/DBFTLUjAxQuba7YlNasguOBkfjOnbq
7ds9ctxDfq9y6jGheHYHC9XIWym7gL/yYa13zzNylDseYQ78Vqk8JPTg/IKTUn8J
QQFTb6/E+3Dt4TLwSM3gh3AvIIwsEtxSwqIO5lEU/ob2cs6Iq3haxuWLrbrof6Ly
/rWbSU1vTCD/TbfwVTPXS4cEsIjM7nRc6Kn0o21RwxIZABXqOpZ3uSvNUHL/SmHl
eHl6/49DRAu9lflWOGZPvhiSu26qJiSlYk3Zu7z5T9lQLndIAnHCQTjqWFlvvkhP
xFijcfP09wlav2nF658PBg==
`pragma protect end_protected
