-- Copyright (C) 2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, the Intel Quartus Prime License Agreement, the Intel
-- MegaCore Function License Agreement, or other applicable 
-- license agreement, including, without limitation, that your
-- use is for the sole purpose of simulating designs for use 
-- exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- Quartus Prime 17.0.1 Build 598 06/07/2017
library IEEE;
use IEEE.std_logic_1164.all;
library work;
use work.TWENTYNM_HIP_COMPONENTS.all;

entity	twentynm_hssi_gen3_x8_pcie_hip	is
	generic (
		-- Entity parameters
		acknack_base	:	bit_vector	:=	B"0000000000000";
		acknack_set	:	string	:=	"false";
		advance_error_reporting	:	string	:=	"disable";
		app_interface_width	:	string	:=	"avst_64bit";
		arb_upfc_30us_counter	:	bit_vector	:=	B"0000";
		arb_upfc_30us_en	:	string	:=	"enable";
		aspm_config_management	:	string	:=	"true";
		aspm_patch_disable	:	string	:=	"enable_both";
		ast_width_rx	:	string	:=	"rx_64";
		ast_width_tx	:	string	:=	"tx_64";
		atomic_malformed	:	string	:=	"false";
		atomic_op_completer_32bit	:	string	:=	"false";
		atomic_op_completer_64bit	:	string	:=	"false";
		atomic_op_routing	:	string	:=	"false";
		auto_msg_drop_enable	:	string	:=	"false";
		avmm_cvp_inter_sel_csr_ctrl	:	string	:=	"disable";
		avmm_dprio_broadcast_en_csr_ctrl	:	string	:=	"disable";
		avmm_force_inter_sel_csr_ctrl	:	string	:=	"disable";
		avmm_power_iso_en_csr_ctrl	:	string	:=	"disable";
		bar0_size_mask	:	bit_vector	:=	B"1111111111111111111111111111";
		bar0_type	:	string	:=	"bar0_64bit_prefetch_mem";
		bar1_size_mask	:	bit_vector	:=	B"0000000000000000000000000000";
		bar1_type	:	string	:=	"bar1_disable";
		bar2_size_mask	:	bit_vector	:=	B"0000000000000000000000000000";
		bar2_type	:	string	:=	"bar2_disable";
		bar3_size_mask	:	bit_vector	:=	B"0000000000000000000000000000";
		bar3_type	:	string	:=	"bar3_disable";
		bar4_size_mask	:	bit_vector	:=	B"0000000000000000000000000000";
		bar4_type	:	string	:=	"bar4_disable";
		bar5_size_mask	:	bit_vector	:=	B"0000000000000000000000000000";
		bar5_type	:	string	:=	"bar5_disable";
		base_counter_sel	:	string	:=	"count_clk_62p5";
		bist_memory_settings	:	string	:=	"000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		bridge_port_ssid_support	:	string	:=	"false";
		bridge_port_vga_enable	:	string	:=	"false";
		bypass_cdc	:	string	:=	"false";
		bypass_clk_switch	:	string	:=	"false";
		bypass_tl	:	string	:=	"false";
		capab_rate_rxcfg_en	:	string	:=	"disable";
		cas_completer_128bit	:	string	:=	"false";
		cdc_clk_relation	:	string	:=	"plesiochronous";
		cdc_dummy_insert_limit	:	bit_vector	:=	B"1011";
		cfg_parchk_ena	:	string	:=	"disable";
		cfgbp_req_recov_disable	:	string	:=	"false";
		class_code	:	bit_vector	:=	B"111111110000000000000000";
		clock_pwr_management	:	string	:=	"false";
		completion_timeout	:	string	:=	"abcd";
		core_clk_divider	:	string	:=	"div_1";
		core_clk_freq_mhz	:	string	:=	"core_clk_250mhz";
		core_clk_out_sel	:	string	:=	"core_clk_out_div_1";
		core_clk_sel	:	string	:=	"pld_clk";
		core_clk_source	:	string	:=	"pll_fixed_clk";
		cseb_bar_match_checking	:	string	:=	"enable";
		cseb_config_bypass	:	string	:=	"disable";
		cseb_cpl_status_during_cvp	:	string	:=	"completer_abort";
		cseb_cpl_tag_checking	:	string	:=	"enable";
		cseb_disable_auto_crs	:	string	:=	"false";
		cseb_extend_pci	:	string	:=	"false";
		cseb_extend_pcie	:	string	:=	"false";
		cseb_min_error_checking	:	string	:=	"false";
		cseb_route_to_avl_rx_st	:	string	:=	"cseb";
		cseb_temp_busy_crs	:	string	:=	"completer_abort_tmp_busy";
		cvp_clk_reset	:	string	:=	"false";
		cvp_data_compressed	:	string	:=	"false";
		cvp_data_encrypted	:	string	:=	"false";
		cvp_enable	:	string	:=	"cvp_dis";
		cvp_mode_reset	:	string	:=	"false";
		cvp_rate_sel	:	string	:=	"full_rate";
		d0_pme	:	string	:=	"false";
		d1_pme	:	string	:=	"false";
		d1_support	:	string	:=	"false";
		d2_pme	:	string	:=	"false";
		d2_support	:	string	:=	"false";
		d3_cold_pme	:	string	:=	"false";
		d3_hot_pme	:	string	:=	"false";
		data_pack_rx	:	string	:=	"disable";
		deemphasis_enable	:	string	:=	"false";
		deskew_comma	:	string	:=	"skp_eieos_deskw";
		device_id	:	bit_vector	:=	B"1110000000000001";
		device_number	:	bit_vector	:=	B"00000";
		device_specific_init	:	string	:=	"false";
		dft_clock_obsrv_en	:	string	:=	"disable";
		dft_clock_obsrv_sel	:	string	:=	"dft_pclk";
		diffclock_nfts_count	:	bit_vector	:=	B"00000000";
		dis_cplovf	:	string	:=	"disable";
		dis_paritychk	:	string	:=	"enable";
		disable_link_x2_support	:	string	:=	"false";
		disable_snoop_packet	:	string	:=	"false";
		dl_tx_check_parity_edb	:	string	:=	"disable";
		dll_active_report_support	:	string	:=	"false";
		early_dl_up	:	string	:=	"true";
		eco_fb332688_dis	:	string	:=	"true";
		ecrc_check_capable	:	string	:=	"true";
		ecrc_gen_capable	:	string	:=	"true";
		egress_block_err_report_ena	:	string	:=	"false";
		ei_delay_powerdown_count	:	bit_vector	:=	B"00001010";
		eie_before_nfts_count	:	bit_vector	:=	B"0100";
		electromech_interlock	:	string	:=	"false";
		en_ieiupdatefc	:	string	:=	"false";
		en_lane_errchk	:	string	:=	"false";
		en_phystatus_dly	:	string	:=	"false";
		ena_ido_cpl	:	string	:=	"false";
		ena_ido_req	:	string	:=	"false";
		enable_adapter_half_rate_mode	:	string	:=	"false";
		enable_ch01_pclk_out	:	string	:=	"pclk_ch0";
		enable_ch0_pclk_out	:	string	:=	"pclk_ch01";
		enable_completion_timeout_disable	:	string	:=	"true";
		enable_directed_spd_chng	:	string	:=	"false";
		enable_function_msix_support	:	string	:=	"true";
		enable_l0s_aspm	:	string	:=	"false";
		enable_l1_aspm	:	string	:=	"false";
		enable_rx_buffer_checking	:	string	:=	"false";
		enable_rx_reordering	:	string	:=	"true";
		enable_slot_register	:	string	:=	"false";
		endpoint_l0_latency	:	bit_vector	:=	B"000";
		endpoint_l1_latency	:	bit_vector	:=	B"000";
		eql_rq_int_en_number	:	bit_vector	:=	B"000000";
		errmgt_fcpe_patch_dis	:	string	:=	"enable";
		errmgt_fep_patch_dis	:	string	:=	"enable";
		expansion_base_address_register	:	string	:=	"00000000000000000000000000000000";
		extend_tag_field	:	string	:=	"false";
		extended_format_field	:	string	:=	"true";
		extended_tag_reset	:	string	:=	"false";
		fc_init_timer	:	bit_vector	:=	B"10000000000";
		flow_control_timeout_count	:	bit_vector	:=	B"11001000";
		flow_control_update_count	:	bit_vector	:=	B"11110";
		flr_capability	:	string	:=	"true";
		force_dis_to_det	:	string	:=	"false";
		force_gen1_dis	:	string	:=	"false";
		force_tx_coeff_preset_lpbk	:	string	:=	"false";
		frame_err_patch_dis	:	string	:=	"enable";
		func_mode	:	string	:=	"disable";
		g3_bypass_equlz	:	string	:=	"false";
		g3_coeff_done_tmout	:	string	:=	"enable";
		g3_deskew_char	:	string	:=	"default_sdsos";
		g3_dis_be_frm_err	:	string	:=	"false";
		g3_dn_rx_hint_eqlz_0	:	bit_vector	:=	B"000";
		g3_dn_rx_hint_eqlz_1	:	bit_vector	:=	B"000";
		g3_dn_rx_hint_eqlz_2	:	bit_vector	:=	B"000";
		g3_dn_rx_hint_eqlz_3	:	bit_vector	:=	B"000";
		g3_dn_rx_hint_eqlz_4	:	bit_vector	:=	B"000";
		g3_dn_rx_hint_eqlz_5	:	bit_vector	:=	B"000";
		g3_dn_rx_hint_eqlz_6	:	bit_vector	:=	B"000";
		g3_dn_rx_hint_eqlz_7	:	bit_vector	:=	B"000";
		g3_dn_tx_preset_eqlz_0	:	bit_vector	:=	B"0000";
		g3_dn_tx_preset_eqlz_1	:	bit_vector	:=	B"0000";
		g3_dn_tx_preset_eqlz_2	:	bit_vector	:=	B"0000";
		g3_dn_tx_preset_eqlz_3	:	bit_vector	:=	B"0000";
		g3_dn_tx_preset_eqlz_4	:	bit_vector	:=	B"0000";
		g3_dn_tx_preset_eqlz_5	:	bit_vector	:=	B"0000";
		g3_dn_tx_preset_eqlz_6	:	bit_vector	:=	B"0000";
		g3_dn_tx_preset_eqlz_7	:	bit_vector	:=	B"0000";
		g3_force_ber_max	:	string	:=	"false";
		g3_force_ber_min	:	string	:=	"false";
		g3_lnk_trn_rx_ts	:	string	:=	"false";
		g3_ltssm_eq_dbg	:	string	:=	"false";
		g3_ltssm_rec_dbg	:	string	:=	"false";
		g3_pause_ltssm_rec_en	:	string	:=	"disable";
		g3_quiesce_guarant	:	string	:=	"false";
		g3_redo_equlz_dis	:	string	:=	"false";
		g3_redo_equlz_en	:	string	:=	"false";
		g3_up_rx_hint_eqlz_0	:	bit_vector	:=	B"000";
		g3_up_rx_hint_eqlz_1	:	bit_vector	:=	B"000";
		g3_up_rx_hint_eqlz_2	:	bit_vector	:=	B"000";
		g3_up_rx_hint_eqlz_3	:	bit_vector	:=	B"000";
		g3_up_rx_hint_eqlz_4	:	bit_vector	:=	B"000";
		g3_up_rx_hint_eqlz_5	:	bit_vector	:=	B"000";
		g3_up_rx_hint_eqlz_6	:	bit_vector	:=	B"000";
		g3_up_rx_hint_eqlz_7	:	bit_vector	:=	B"000";
		g3_up_tx_preset_eqlz_0	:	bit_vector	:=	B"0000";
		g3_up_tx_preset_eqlz_1	:	bit_vector	:=	B"0000";
		g3_up_tx_preset_eqlz_2	:	bit_vector	:=	B"0000";
		g3_up_tx_preset_eqlz_3	:	bit_vector	:=	B"0000";
		g3_up_tx_preset_eqlz_4	:	bit_vector	:=	B"0000";
		g3_up_tx_preset_eqlz_5	:	bit_vector	:=	B"0000";
		g3_up_tx_preset_eqlz_6	:	bit_vector	:=	B"0000";
		g3_up_tx_preset_eqlz_7	:	bit_vector	:=	B"0000";
		gen123_lane_rate_mode	:	string	:=	"gen1_rate";
		gen2_diffclock_nfts_count	:	bit_vector	:=	B"11111111";
		gen2_pma_pll_usage	:	string	:=	"not_applicaple";
		gen2_sameclock_nfts_count	:	bit_vector	:=	B"11111111";
		gen3_coeff_1	:	bit_vector	:=	B"000000000000000100";
		gen3_coeff_10	:	bit_vector	:=	B"000000000000000111";
		gen3_coeff_10_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_10_nxtber_less	:	bit_vector	:=	B"1111";
		gen3_coeff_10_nxtber_more	:	bit_vector	:=	B"1010";
		gen3_coeff_10_preset_hint	:	bit_vector	:=	B"011";
		gen3_coeff_10_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_10_sel	:	string	:=	"preset_10";
		gen3_coeff_11	:	bit_vector	:=	B"000000000000000111";
		gen3_coeff_11_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_11_nxtber_less	:	bit_vector	:=	B"1111";
		gen3_coeff_11_nxtber_more	:	bit_vector	:=	B"1111";
		gen3_coeff_11_preset_hint	:	bit_vector	:=	B"100";
		gen3_coeff_11_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_11_sel	:	string	:=	"preset_11";
		gen3_coeff_12	:	bit_vector	:=	B"000000000000000111";
		gen3_coeff_12_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_12_nxtber_less	:	bit_vector	:=	B"1111";
		gen3_coeff_12_nxtber_more	:	bit_vector	:=	B"1111";
		gen3_coeff_12_preset_hint	:	bit_vector	:=	B"010";
		gen3_coeff_12_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_12_sel	:	string	:=	"preset_12";
		gen3_coeff_13	:	bit_vector	:=	B"000000000000000100";
		gen3_coeff_13_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_13_nxtber_less	:	bit_vector	:=	B"1101";
		gen3_coeff_13_nxtber_more	:	bit_vector	:=	B"0001";
		gen3_coeff_13_preset_hint	:	bit_vector	:=	B"100";
		gen3_coeff_13_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_13_sel	:	string	:=	"preset_13";
		gen3_coeff_14	:	bit_vector	:=	B"000000000000000100";
		gen3_coeff_14_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_14_nxtber_less	:	bit_vector	:=	B"1111";
		gen3_coeff_14_nxtber_more	:	bit_vector	:=	B"0010";
		gen3_coeff_14_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_14_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_14_sel	:	string	:=	"preset_14";
		gen3_coeff_15	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_15_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_15_nxtber_less	:	bit_vector	:=	B"0000";
		gen3_coeff_15_nxtber_more	:	bit_vector	:=	B"0000";
		gen3_coeff_15_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_15_reqber	:	bit_vector	:=	B"00000";
		gen3_coeff_15_sel	:	string	:=	"coeff_15";
		gen3_coeff_16	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_16_ber_meas	:	bit_vector	:=	B"000000";
		gen3_coeff_16_nxtber_less	:	bit_vector	:=	B"0000";
		gen3_coeff_16_nxtber_more	:	bit_vector	:=	B"0000";
		gen3_coeff_16_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_16_reqber	:	bit_vector	:=	B"00000";
		gen3_coeff_16_sel	:	string	:=	"coeff_16";
		gen3_coeff_17	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_17_ber_meas	:	bit_vector	:=	B"000000";
		gen3_coeff_17_nxtber_less	:	bit_vector	:=	B"0000";
		gen3_coeff_17_nxtber_more	:	bit_vector	:=	B"0000";
		gen3_coeff_17_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_17_reqber	:	bit_vector	:=	B"00000";
		gen3_coeff_17_sel	:	string	:=	"coeff_17";
		gen3_coeff_18	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_18_ber_meas	:	bit_vector	:=	B"000000";
		gen3_coeff_18_nxtber_less	:	bit_vector	:=	B"0000";
		gen3_coeff_18_nxtber_more	:	bit_vector	:=	B"0000";
		gen3_coeff_18_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_18_reqber	:	bit_vector	:=	B"00000";
		gen3_coeff_18_sel	:	string	:=	"coeff_18";
		gen3_coeff_19	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_19_ber_meas	:	bit_vector	:=	B"000000";
		gen3_coeff_19_nxtber_less	:	bit_vector	:=	B"0000";
		gen3_coeff_19_nxtber_more	:	bit_vector	:=	B"0000";
		gen3_coeff_19_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_19_reqber	:	bit_vector	:=	B"00000";
		gen3_coeff_19_sel	:	string	:=	"coeff_19";
		gen3_coeff_1_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_1_nxtber_less	:	bit_vector	:=	B"1100";
		gen3_coeff_1_nxtber_more	:	bit_vector	:=	B"0110";
		gen3_coeff_1_preset_hint	:	bit_vector	:=	B"010";
		gen3_coeff_1_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_1_sel	:	string	:=	"preset_1";
		gen3_coeff_2	:	bit_vector	:=	B"000000000000000001";
		gen3_coeff_20	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_20_ber_meas	:	bit_vector	:=	B"000000";
		gen3_coeff_20_nxtber_less	:	bit_vector	:=	B"0000";
		gen3_coeff_20_nxtber_more	:	bit_vector	:=	B"0000";
		gen3_coeff_20_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_20_reqber	:	bit_vector	:=	B"00000";
		gen3_coeff_20_sel	:	string	:=	"coeff_20";
		gen3_coeff_21	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_21_ber_meas	:	bit_vector	:=	B"000000";
		gen3_coeff_21_nxtber_less	:	bit_vector	:=	B"0000";
		gen3_coeff_21_nxtber_more	:	bit_vector	:=	B"0000";
		gen3_coeff_21_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_21_reqber	:	bit_vector	:=	B"00000";
		gen3_coeff_21_sel	:	string	:=	"coeff_21";
		gen3_coeff_22	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_22_ber_meas	:	bit_vector	:=	B"000000";
		gen3_coeff_22_nxtber_less	:	bit_vector	:=	B"0000";
		gen3_coeff_22_nxtber_more	:	bit_vector	:=	B"0000";
		gen3_coeff_22_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_22_reqber	:	bit_vector	:=	B"00000";
		gen3_coeff_22_sel	:	string	:=	"coeff_22";
		gen3_coeff_23	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_23_ber_meas	:	bit_vector	:=	B"000000";
		gen3_coeff_23_nxtber_less	:	bit_vector	:=	B"0000";
		gen3_coeff_23_nxtber_more	:	bit_vector	:=	B"0000";
		gen3_coeff_23_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_23_reqber	:	bit_vector	:=	B"00000";
		gen3_coeff_23_sel	:	string	:=	"coeff_23";
		gen3_coeff_24	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_24_ber_meas	:	bit_vector	:=	B"000000";
		gen3_coeff_24_nxtber_less	:	bit_vector	:=	B"0000";
		gen3_coeff_24_nxtber_more	:	bit_vector	:=	B"0000";
		gen3_coeff_24_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_24_reqber	:	bit_vector	:=	B"00000";
		gen3_coeff_24_sel	:	string	:=	"coeff_24";
		gen3_coeff_2_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_2_nxtber_less	:	bit_vector	:=	B"0010";
		gen3_coeff_2_nxtber_more	:	bit_vector	:=	B"0100";
		gen3_coeff_2_preset_hint	:	bit_vector	:=	B"100";
		gen3_coeff_2_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_2_sel	:	string	:=	"preset_2";
		gen3_coeff_3	:	bit_vector	:=	B"000000000000000001";
		gen3_coeff_3_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_3_nxtber_less	:	bit_vector	:=	B"1111";
		gen3_coeff_3_nxtber_more	:	bit_vector	:=	B"0011";
		gen3_coeff_3_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_3_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_3_sel	:	string	:=	"preset_3";
		gen3_coeff_4	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_4_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_4_nxtber_less	:	bit_vector	:=	B"1111";
		gen3_coeff_4_nxtber_more	:	bit_vector	:=	B"0100";
		gen3_coeff_4_preset_hint	:	bit_vector	:=	B"000";
		gen3_coeff_4_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_4_sel	:	string	:=	"preset_4";
		gen3_coeff_5	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_5_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_5_nxtber_less	:	bit_vector	:=	B"1111";
		gen3_coeff_5_nxtber_more	:	bit_vector	:=	B"0101";
		gen3_coeff_5_preset_hint	:	bit_vector	:=	B"100";
		gen3_coeff_5_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_5_sel	:	string	:=	"preset_5";
		gen3_coeff_6	:	bit_vector	:=	B"000000000000000111";
		gen3_coeff_6_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_6_nxtber_less	:	bit_vector	:=	B"1111";
		gen3_coeff_6_nxtber_more	:	bit_vector	:=	B"1111";
		gen3_coeff_6_preset_hint	:	bit_vector	:=	B"100";
		gen3_coeff_6_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_6_sel	:	string	:=	"preset_6";
		gen3_coeff_7	:	bit_vector	:=	B"000000000000000001";
		gen3_coeff_7_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_7_nxtber_less	:	bit_vector	:=	B"0001";
		gen3_coeff_7_nxtber_more	:	bit_vector	:=	B"0111";
		gen3_coeff_7_preset_hint	:	bit_vector	:=	B"010";
		gen3_coeff_7_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_7_sel	:	string	:=	"preset_7";
		gen3_coeff_8	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_8_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_8_nxtber_less	:	bit_vector	:=	B"0100";
		gen3_coeff_8_nxtber_more	:	bit_vector	:=	B"1000";
		gen3_coeff_8_preset_hint	:	bit_vector	:=	B"010";
		gen3_coeff_8_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_8_sel	:	string	:=	"preset_8";
		gen3_coeff_9	:	bit_vector	:=	B"000000000000000000";
		gen3_coeff_9_ber_meas	:	bit_vector	:=	B"000010";
		gen3_coeff_9_nxtber_less	:	bit_vector	:=	B"1011";
		gen3_coeff_9_nxtber_more	:	bit_vector	:=	B"1001";
		gen3_coeff_9_preset_hint	:	bit_vector	:=	B"011";
		gen3_coeff_9_reqber	:	bit_vector	:=	B"01000";
		gen3_coeff_9_sel	:	string	:=	"preset_9";
		gen3_coeff_delay_count	:	bit_vector	:=	B"1111101";
		gen3_coeff_errchk	:	string	:=	"enable";
		gen3_dcbal_en	:	string	:=	"true";
		gen3_diffclock_nfts_count	:	bit_vector	:=	B"10000000";
		gen3_force_local_coeff	:	string	:=	"false";
		gen3_full_swing	:	bit_vector	:=	B"111111";
		gen3_half_swing	:	string	:=	"false";
		gen3_low_freq	:	bit_vector	:=	B"000001";
		gen3_paritychk	:	string	:=	"enable";
		gen3_pl_framing_err_dis	:	string	:=	"enable";
		gen3_preset_coeff_1	:	bit_vector	:=	B"000000110101001010";
		gen3_preset_coeff_10	:	bit_vector	:=	B"001011110100000000";
		gen3_preset_coeff_11	:	bit_vector	:=	B"011110100001000000";
		gen3_preset_coeff_2	:	bit_vector	:=	B"000000110100001011";
		gen3_preset_coeff_3	:	bit_vector	:=	B"000000110010001101";
		gen3_preset_coeff_4	:	bit_vector	:=	B"000000110111001000";
		gen3_preset_coeff_5	:	bit_vector	:=	B"000000111111000000";
		gen3_preset_coeff_6	:	bit_vector	:=	B"000110111001000000";
		gen3_preset_coeff_7	:	bit_vector	:=	B"001000110111000000";
		gen3_preset_coeff_8	:	bit_vector	:=	B"000110101100001101";
		gen3_preset_coeff_9	:	bit_vector	:=	B"001000101111001000";
		gen3_reset_eieos_cnt_bit	:	string	:=	"false";
		gen3_rxfreqlock_counter	:	bit_vector	:=	B"00000000000000000000";
		gen3_sameclock_nfts_count	:	bit_vector	:=	B"10000000";
		gen3_scrdscr_bypass	:	string	:=	"false";
		gen3_skip_ph2_ph3	:	string	:=	"false";
		hard_reset_bypass	:	string	:=	"false";
		hard_rst_sig_chnl_en	:	string	:=	"disable_hrc_sig";
		hard_rst_tx_pll_rst_chnl_en	:	string	:=	"disable_hrc_txpll_rst";
		hip_ac_pwr_clk_freq_in_hz	:	bit_vector	:=	B"000000000000000000000000000000";
		hip_ac_pwr_uw_per_mhz	:	bit_vector	:=	B"000000000000000000000000000000";
		hip_base_address	:	bit_vector	:=	B"0000000000";
		hip_clock_dis	:	string	:=	"enable_hip_clk";
		hip_hard_reset	:	string	:=	"enable";
		hip_pcs_sig_chnl_en	:	string	:=	"disable_hip_pcs_sig";
		hot_plug_support	:	bit_vector	:=	B"0000000";
		hrc_chnl_txpll_master_cgb_rst_select	:	string	:=	"disable_master_cgb_sel";
		hrdrstctrl_en	:	string	:=	"hrdrstctrl_dis";
		iei_enable_settings	:	string	:=	"gen3gen2_infei_infsd_gen1_infei_sd";
		indicator	:	bit_vector	:=	B"111";
		intel_id_access	:	string	:=	"false";
		interrupt_pin	:	string	:=	"inta";
		io_window_addr_width	:	string	:=	"window_32_bit";
		jtag_id	:	string	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		ko_compl_data	:	bit_vector	:=	B"000000000000";
		ko_compl_header	:	bit_vector	:=	B"000000000000";
		l01_entry_latency	:	bit_vector	:=	B"11111";
		l0_exit_latency_diffclock	:	bit_vector	:=	B"110";
		l0_exit_latency_sameclock	:	bit_vector	:=	B"110";
		l0s_adj_rply_timer_dis	:	string	:=	"enable";
		l1_exit_latency_diffclock	:	bit_vector	:=	B"000";
		l1_exit_latency_sameclock	:	bit_vector	:=	B"000";
		l2_async_logic	:	string	:=	"enable";
		lane_mask	:	string	:=	"ln_mask_x4";
		lane_rate	:	string	:=	"gen1";
		link_width	:	string	:=	"x1";
		lmi_hold_off_cfg_timer_en	:	string	:=	"disable";
		low_priority_vc	:	string	:=	"single_vc_low_pr";
		ltr_mechanism	:	string	:=	"false";
		ltssm_1ms_timeout	:	string	:=	"disable";
		ltssm_freqlocked_check	:	string	:=	"disable";
		malformed_tlp_truncate_en	:	string	:=	"disable";
		max_link_width	:	string	:=	"x4_link_width";
		max_payload_size	:	string	:=	"payload_512";
		maximum_current	:	bit_vector	:=	B"000";
		millisecond_cycle_count	:	bit_vector	:=	B"00000000000000000000";
		msi_64bit_addressing_capable	:	string	:=	"true";
		msi_masking_capable	:	string	:=	"false";
		msi_multi_message_capable	:	string	:=	"count_4";
		msi_support	:	string	:=	"true";
		msix_pba_bir	:	bit_vector	:=	B"000";
		msix_pba_offset	:	bit_vector	:=	B"00000000000000000000000000000";
		msix_table_bir	:	bit_vector	:=	B"000";
		msix_table_offset	:	bit_vector	:=	B"00000000000000000000000000000";
		msix_table_size	:	bit_vector	:=	B"00000000000";
		national_inst_thru_enhance	:	string	:=	"true";
		no_command_completed	:	string	:=	"true";
		no_soft_reset	:	string	:=	"false";
		not_use_k_gbl_bits	:	string	:=	"not_used_k_gbl";
		operating_voltage	:	string	:=	"standard";
		pcie_base_spec	:	string	:=	"pcie_2p1";
		pcie_mode	:	string	:=	"shared_mode";
		pcie_spec_1p0_compliance	:	string	:=	"spec_1p1";
		pcie_spec_version	:	string	:=	"v2";
		pclk_out_sel	:	string	:=	"pclk";
		pld_in_use_reg	:	string	:=	"false";
		pm_latency_patch_dis	:	string	:=	"enable";
		pm_txdl_patch_dis	:	string	:=	"enable";
		pme_clock	:	string	:=	"false";
		port_link_number	:	bit_vector	:=	B"00000001";
		port_type	:	string	:=	"native_ep";
		powerdown_mode	:	string	:=	"powerup";
		prefetchable_mem_window_addr_width	:	string	:=	"prefetch_32";
		r2c_mask_easy	:	string	:=	"false";
		r2c_mask_enable	:	string	:=	"false";
		rec_frqlk_mon_en	:	string	:=	"disable";
		register_pipe_signals	:	string	:=	"true";
		retry_buffer_last_active_address	:	bit_vector	:=	B"1111111111";
		retry_buffer_memory_settings	:	string	:=	"000000000000000000000000000000000000";
		retry_ecc_corr_mask_dis	:	string	:=	"enable";
		revision_id	:	bit_vector	:=	B"00000001";
		role_based_error_reporting	:	string	:=	"false";
		rp_bug_fix_pri_sec_stat_reg	:	bit_vector	:=	B"1111111";
		rpltim_base	:	bit_vector	:=	B"00000000000000";
		rpltim_set	:	string	:=	"false";
		rstctl_ltssm_dis	:	string	:=	"false";
		rstctrl_1ms_count_fref_clk	:	bit_vector	:=	B"00001111010000100100";
		rstctrl_1us_count_fref_clk	:	bit_vector	:=	B"00000000000000111111";
		rstctrl_altpe3_crst_n_inv	:	string	:=	"false";
		rstctrl_altpe3_rst_n_inv	:	string	:=	"false";
		rstctrl_altpe3_srst_n_inv	:	string	:=	"false";
		rstctrl_chnl_cal_done_select	:	string	:=	"not_active_chnl_cal_done";
		rstctrl_debug_en	:	string	:=	"false";
		rstctrl_force_inactive_rst	:	string	:=	"false";
		rstctrl_fref_clk_select	:	string	:=	"ch0_sel";
		rstctrl_hard_block_enable	:	string	:=	"hard_rst_ctl";
		rstctrl_hip_ep	:	string	:=	"hip_ep";
		rstctrl_mask_tx_pll_lock_select	:	string	:=	"not_active_mask_tx_pll_lock";
		rstctrl_perst_enable	:	string	:=	"level";
		rstctrl_perstn_select	:	string	:=	"perstn_pin";
		rstctrl_pld_clr	:	string	:=	"false";
		rstctrl_pll_cal_done_select	:	string	:=	"not_active_pll_cal_done";
		rstctrl_rx_pcs_rst_n_inv	:	string	:=	"false";
		rstctrl_rx_pcs_rst_n_select	:	string	:=	"not_active_rx_pcs_rst";
		rstctrl_rx_pll_freq_lock_select	:	string	:=	"not_active_rx_pll_f_lock";
		rstctrl_rx_pll_lock_select	:	string	:=	"not_active_rx_pll_lock";
		rstctrl_rx_pma_rstb_inv	:	string	:=	"false";
		rstctrl_rx_pma_rstb_select	:	string	:=	"not_active_rx_pma_rstb";
		rstctrl_timer_a	:	bit_vector	:=	B"00001010";
		rstctrl_timer_a_type	:	string	:=	"a_timer_milli_secs";
		rstctrl_timer_b	:	bit_vector	:=	B"00001010";
		rstctrl_timer_b_type	:	string	:=	"b_timer_milli_secs";
		rstctrl_timer_c	:	bit_vector	:=	B"00001010";
		rstctrl_timer_c_type	:	string	:=	"c_timer_milli_secs";
		rstctrl_timer_d	:	bit_vector	:=	B"00010100";
		rstctrl_timer_d_type	:	string	:=	"d_timer_milli_secs";
		rstctrl_timer_e	:	bit_vector	:=	B"00000001";
		rstctrl_timer_e_type	:	string	:=	"e_timer_milli_secs";
		rstctrl_timer_f	:	bit_vector	:=	B"00001010";
		rstctrl_timer_f_type	:	string	:=	"f_timer_milli_secs";
		rstctrl_timer_g	:	bit_vector	:=	B"00001010";
		rstctrl_timer_g_type	:	string	:=	"g_timer_milli_secs";
		rstctrl_timer_h	:	bit_vector	:=	B"00000100";
		rstctrl_timer_h_type	:	string	:=	"h_timer_milli_secs";
		rstctrl_timer_i	:	bit_vector	:=	B"00010100";
		rstctrl_timer_i_type	:	string	:=	"i_timer_milli_secs";
		rstctrl_timer_j	:	bit_vector	:=	B"00010100";
		rstctrl_timer_j_type	:	string	:=	"j_timer_milli_secs";
		rstctrl_tx_lcff_pll_lock_select	:	string	:=	"not_active_lcff_pll_lock";
		rstctrl_tx_lcff_pll_rstb_select	:	string	:=	"not_active_lcff_pll_rstb";
		rstctrl_tx_pcs_rst_n_inv	:	string	:=	"false";
		rstctrl_tx_pcs_rst_n_select	:	string	:=	"not_active_tx_pcs_rst";
		rstctrl_tx_pma_rstb_inv	:	string	:=	"false";
		rstctrl_tx_pma_syncp_inv	:	string	:=	"false";
		rstctrl_tx_pma_syncp_select	:	string	:=	"not_active_tx_pma_syncp";
		rx_ast_parity	:	string	:=	"disable";
		rx_buffer_credit_alloc	:	string	:=	"balance";
		rx_buffer_fc_protect	:	bit_vector	:=	B"00000000000001000100";
		rx_buffer_protect	:	bit_vector	:=	B"00001000100";
		rx_cdc_almost_empty	:	bit_vector	:=	B"0011";
		rx_cdc_almost_full	:	bit_vector	:=	B"1100";
		rx_cred_ctl_param	:	string	:=	"disable";
		rx_ei_l0s	:	string	:=	"disable";
		rx_l0s_count_idl	:	bit_vector	:=	B"00000000";
		rx_ptr0_nonposted_dpram_max	:	bit_vector	:=	B"00000000000";
		rx_ptr0_nonposted_dpram_min	:	bit_vector	:=	B"00000000000";
		rx_ptr0_posted_dpram_max	:	bit_vector	:=	B"00000000000";
		rx_ptr0_posted_dpram_min	:	bit_vector	:=	B"00000000000";
		rx_runt_patch_dis	:	string	:=	"enable";
		rx_sop_ctrl	:	string	:=	"rx_sop_boundary_64";
		rx_trunc_patch_dis	:	string	:=	"enable";
		rx_use_prst	:	string	:=	"false";
		rx_use_prst_ep	:	string	:=	"true";
		rxbuf_ecc_corr_mask_dis	:	string	:=	"enable";
		rxdl_bad_sop_eop_filter_dis	:	string	:=	"rxdlbug1_enable_both";
		rxdl_bad_tlp_patch_dis	:	string	:=	"rxdlbug2_enable_both";
		rxdl_lcrc_patch_dis	:	string	:=	"rxdlbug3_enable_both";
		sameclock_nfts_count	:	bit_vector	:=	B"00000000";
		sel_enable_pcs_rx_fifo_err	:	string	:=	"disable_sel";
		silicon_rev	:	string	:=	"20nm5es";
		sim_mode	:	string	:=	"disable";
		simple_ro_fifo_control_en	:	string	:=	"disable";
		single_rx_detect	:	string	:=	"detect_all_lanes";
		skp_os_gen3_count	:	bit_vector	:=	B"00000000000";
		skp_os_schedule_count	:	bit_vector	:=	B"00000000000";
		slot_number	:	bit_vector	:=	B"0000000000000";
		slot_power_limit	:	bit_vector	:=	B"00000000";
		slot_power_scale	:	bit_vector	:=	B"00";
		slotclk_cfg	:	string	:=	"static_slotclkcfgon";
		ssid	:	bit_vector	:=	B"0000000000000000";
		ssvid	:	bit_vector	:=	B"0000000000000000";
		subsystem_device_id	:	bit_vector	:=	B"1110000000000001";
		subsystem_vendor_id	:	bit_vector	:=	B"0001000101110010";
		sup_mode	:	string	:=	"user_mode";
		surprise_down_error_support	:	string	:=	"false";
		tl_cfg_div	:	string	:=	"cfg_clk_div_7";
		tl_tx_check_parity_msg	:	string	:=	"disable";
		tph_completer	:	string	:=	"false";
		tx_ast_parity	:	string	:=	"disable";
		tx_cdc_almost_empty	:	bit_vector	:=	B"0101";
		tx_cdc_almost_full	:	bit_vector	:=	B"1100";
		tx_sop_ctrl	:	string	:=	"boundary_64";
		tx_swing	:	bit_vector	:=	B"00000000";
		txdl_fair_arbiter_counter	:	bit_vector	:=	B"0000";
		txdl_fair_arbiter_en	:	string	:=	"enable";
		txrate_adv	:	string	:=	"capability";
		uc_calibration_en	:	string	:=	"uc_calibration_dis";
		use_aer	:	string	:=	"false";
		use_crc_forwarding	:	string	:=	"false";
		user_id	:	bit_vector	:=	B"0000000000000000";
		vc0_clk_enable	:	string	:=	"true";
		vc0_rx_buffer_memory_settings	:	string	:=	"000000000000000000000000000000000000";
		vc0_rx_flow_ctrl_compl_data	:	bit_vector	:=	B"000111000000";
		vc0_rx_flow_ctrl_compl_header	:	bit_vector	:=	B"01110000";
		vc0_rx_flow_ctrl_nonposted_data	:	bit_vector	:=	B"00000000";
		vc0_rx_flow_ctrl_nonposted_header	:	bit_vector	:=	B"00110110";
		vc0_rx_flow_ctrl_posted_data	:	bit_vector	:=	B"000101101000";
		vc0_rx_flow_ctrl_posted_header	:	bit_vector	:=	B"00110010";
		vc1_clk_enable	:	string	:=	"false";
		vc_arbitration	:	string	:=	"single_vc_arb";
		vc_enable	:	string	:=	"single_vc";
		vendor_id	:	bit_vector	:=	B"0001000101110010";
		vsec_cap	:	bit_vector	:=	B"0000";
		vsec_id	:	bit_vector	:=	B"0001000101110010";
		wrong_device_id	:	string	:=	"disable"
	);
	port (
		-- Entity ports
		aer_msi_num	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		app_int_err	:	in	std_logic_vector(1 downto 0)	:=	"00";
		app_inta_sts	:	in	std_logic	:=	'0';
		app_msi_num	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		app_msi_req	:	in	std_logic	:=	'0';
		app_msi_tc	:	in	std_logic_vector(2 downto 0)	:=	"000";
		atpg_los_en_n	:	in	std_logic	:=	'0';
		avmm_address	:	in	std_logic_vector(9 downto 0)	:=	"0000000000";
		avmm_byte_en	:	in	std_logic_vector(1 downto 0)	:=	"00";
		avmm_clk	:	in	std_logic	:=	'0';
		avmm_read	:	in	std_logic	:=	'0';
		avmm_rst_n	:	in	std_logic	:=	'0';
		avmm_write	:	in	std_logic	:=	'0';
		avmm_writedata	:	in	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		bist_scanen	:	in	std_logic	:=	'0';
		bist_scanin	:	in	std_logic	:=	'0';
		bisten_rcv_n	:	in	std_logic	:=	'0';
		bisten_rpl_n	:	in	std_logic	:=	'0';
		bistmode_n	:	in	std_logic	:=	'0';
		cfg_link2csr_pld	:	in	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		cfg_prmbus_pld	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		chnl_cal_done0	:	in	std_logic	:=	'0';
		chnl_cal_done1	:	in	std_logic	:=	'0';
		chnl_cal_done2	:	in	std_logic	:=	'0';
		chnl_cal_done3	:	in	std_logic	:=	'0';
		chnl_cal_done4	:	in	std_logic	:=	'0';
		chnl_cal_done5	:	in	std_logic	:=	'0';
		chnl_cal_done6	:	in	std_logic	:=	'0';
		chnl_cal_done7	:	in	std_logic	:=	'0';
		core_clk_in	:	in	std_logic	:=	'0';
		core_crst	:	in	std_logic	:=	'0';
		core_por	:	in	std_logic	:=	'0';
		core_rst	:	in	std_logic	:=	'0';
		core_srst	:	in	std_logic	:=	'0';
		cpl_err	:	in	std_logic_vector(6 downto 0)	:=	"0000000";
		cpl_pending	:	in	std_logic	:=	'0';
		cseb_rddata	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		cseb_rddata_parity	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		cseb_rdresponse	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		cseb_waitrequest	:	in	std_logic	:=	'0';
		cseb_wrresp_valid	:	in	std_logic	:=	'0';
		cseb_wrresponse	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		csr_cbdin	:	in	std_logic	:=	'0';
		csr_clk	:	in	std_logic	:=	'0';
		csr_din	:	in	std_logic	:=	'0';
		csr_en	:	in	std_logic	:=	'0';
		csr_enscan	:	in	std_logic	:=	'0';
		csr_entest	:	in	std_logic	:=	'0';
		csr_in	:	in	std_logic	:=	'0';
		csr_load_csr	:	in	std_logic	:=	'0';
		csr_pipe_in	:	in	std_logic	:=	'0';
		csr_seg	:	in	std_logic	:=	'0';
		csr_tcsrin	:	in	std_logic	:=	'0';
		csr_tverify	:	in	std_logic	:=	'0';
		cvp_config_done	:	in	std_logic	:=	'0';
		cvp_config_error	:	in	std_logic	:=	'0';
		cvp_config_ready	:	in	std_logic	:=	'0';
		cvp_en	:	in	std_logic	:=	'0';
		egress_blk_err	:	in	std_logic	:=	'0';
		entest	:	in	std_logic	:=	'0';
		flr_reset	:	in	std_logic	:=	'0';
		force_tx_eidle	:	in	std_logic	:=	'0';
		fref_clk0	:	in	std_logic	:=	'0';
		fref_clk1	:	in	std_logic	:=	'0';
		fref_clk2	:	in	std_logic	:=	'0';
		fref_clk3	:	in	std_logic	:=	'0';
		fref_clk4	:	in	std_logic	:=	'0';
		fref_clk5	:	in	std_logic	:=	'0';
		fref_clk6	:	in	std_logic	:=	'0';
		fref_clk7	:	in	std_logic	:=	'0';
		frzlogic	:	in	std_logic	:=	'0';
		frzreg	:	in	std_logic	:=	'0';
		hold_ltssm_rec	:	in	std_logic	:=	'0';
		hpg_ctrler	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		iocsrrdy_dly	:	in	std_logic	:=	'0';
		lmi_addr	:	in	std_logic_vector(11 downto 0)	:=	"000000000000";
		lmi_din	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		lmi_rden	:	in	std_logic	:=	'0';
		lmi_wren	:	in	std_logic	:=	'0';
		m10k_select	:	in	std_logic_vector(2 downto 0)	:=	"000";
		mask_tx_pll_lock0	:	in	std_logic	:=	'0';
		mask_tx_pll_lock1	:	in	std_logic	:=	'0';
		mask_tx_pll_lock2	:	in	std_logic	:=	'0';
		mask_tx_pll_lock3	:	in	std_logic	:=	'0';
		mask_tx_pll_lock4	:	in	std_logic	:=	'0';
		mask_tx_pll_lock5	:	in	std_logic	:=	'0';
		mask_tx_pll_lock6	:	in	std_logic	:=	'0';
		mask_tx_pll_lock7	:	in	std_logic	:=	'0';
		mem_hip_test_enable	:	in	std_logic	:=	'0';
		mem_regscanen_n	:	in	std_logic	:=	'0';
		mem_rscin_rcv_bot	:	in	std_logic	:=	'0';
		mem_rscin_rcv_top	:	in	std_logic	:=	'0';
		mem_rscin_rtry	:	in	std_logic	:=	'0';
		nfrzdrv	:	in	std_logic	:=	'0';
		npor	:	in	std_logic	:=	'0';
		pclk_central	:	in	std_logic	:=	'0';
		pclk_ch0	:	in	std_logic	:=	'0';
		pclk_ch1	:	in	std_logic	:=	'0';
		pex_msi_num	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		phy_rst	:	in	std_logic	:=	'0';
		phy_srst	:	in	std_logic	:=	'0';
		phystatus0	:	in	std_logic	:=	'0';
		phystatus1	:	in	std_logic	:=	'0';
		phystatus2	:	in	std_logic	:=	'0';
		phystatus3	:	in	std_logic	:=	'0';
		phystatus4	:	in	std_logic	:=	'0';
		phystatus5	:	in	std_logic	:=	'0';
		phystatus6	:	in	std_logic	:=	'0';
		phystatus7	:	in	std_logic	:=	'0';
		pin_perst_n	:	in	std_logic	:=	'0';
		pld_clk	:	in	std_logic	:=	'0';
		pld_clrhip_n	:	in	std_logic	:=	'0';
		pld_clrpcship_n	:	in	std_logic	:=	'0';
		pld_clrpmapcship_n	:	in	std_logic	:=	'0';
		pld_core_ready	:	in	std_logic	:=	'0';
		pld_gp_status	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		pld_perst_n	:	in	std_logic	:=	'0';
		pll_cal_done0	:	in	std_logic	:=	'0';
		pll_cal_done1	:	in	std_logic	:=	'0';
		pll_cal_done2	:	in	std_logic	:=	'0';
		pll_cal_done3	:	in	std_logic	:=	'0';
		pll_cal_done4	:	in	std_logic	:=	'0';
		pll_cal_done5	:	in	std_logic	:=	'0';
		pll_cal_done6	:	in	std_logic	:=	'0';
		pll_cal_done7	:	in	std_logic	:=	'0';
		pll_fixed_clk_central	:	in	std_logic	:=	'0';
		pll_fixed_clk_ch0	:	in	std_logic	:=	'0';
		pll_fixed_clk_ch1	:	in	std_logic	:=	'0';
		plniotri	:	in	std_logic	:=	'0';
		pm_auxpwr	:	in	std_logic	:=	'0';
		pm_data	:	in	std_logic_vector(9 downto 0)	:=	"0000000000";
		pm_event	:	in	std_logic	:=	'0';
		pm_exit_d0_ack	:	in	std_logic	:=	'0';
		pme_to_cr	:	in	std_logic	:=	'0';
		reserved_clk_in	:	in	std_logic	:=	'0';
		reserved_in	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		rx_cred_ctl	:	in	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		rx_pll_freq_lock0	:	in	std_logic	:=	'0';
		rx_pll_freq_lock1	:	in	std_logic	:=	'0';
		rx_pll_freq_lock2	:	in	std_logic	:=	'0';
		rx_pll_freq_lock3	:	in	std_logic	:=	'0';
		rx_pll_freq_lock4	:	in	std_logic	:=	'0';
		rx_pll_freq_lock5	:	in	std_logic	:=	'0';
		rx_pll_freq_lock6	:	in	std_logic	:=	'0';
		rx_pll_freq_lock7	:	in	std_logic	:=	'0';
		rx_pll_phase_lock0	:	in	std_logic	:=	'0';
		rx_pll_phase_lock1	:	in	std_logic	:=	'0';
		rx_pll_phase_lock2	:	in	std_logic	:=	'0';
		rx_pll_phase_lock3	:	in	std_logic	:=	'0';
		rx_pll_phase_lock4	:	in	std_logic	:=	'0';
		rx_pll_phase_lock5	:	in	std_logic	:=	'0';
		rx_pll_phase_lock6	:	in	std_logic	:=	'0';
		rx_pll_phase_lock7	:	in	std_logic	:=	'0';
		rx_st_mask	:	in	std_logic	:=	'0';
		rx_st_ready	:	in	std_logic	:=	'0';
		rxblkst0	:	in	std_logic	:=	'0';
		rxblkst1	:	in	std_logic	:=	'0';
		rxblkst2	:	in	std_logic	:=	'0';
		rxblkst3	:	in	std_logic	:=	'0';
		rxblkst4	:	in	std_logic	:=	'0';
		rxblkst5	:	in	std_logic	:=	'0';
		rxblkst6	:	in	std_logic	:=	'0';
		rxblkst7	:	in	std_logic	:=	'0';
		rxdata0	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata1	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata2	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata3	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata4	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata5	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata6	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata7	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdatak0	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak1	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak2	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak3	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak4	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak5	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak6	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak7	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdataskip0	:	in	std_logic	:=	'0';
		rxdataskip1	:	in	std_logic	:=	'0';
		rxdataskip2	:	in	std_logic	:=	'0';
		rxdataskip3	:	in	std_logic	:=	'0';
		rxdataskip4	:	in	std_logic	:=	'0';
		rxdataskip5	:	in	std_logic	:=	'0';
		rxdataskip6	:	in	std_logic	:=	'0';
		rxdataskip7	:	in	std_logic	:=	'0';
		rxelecidle0	:	in	std_logic	:=	'0';
		rxelecidle1	:	in	std_logic	:=	'0';
		rxelecidle2	:	in	std_logic	:=	'0';
		rxelecidle3	:	in	std_logic	:=	'0';
		rxelecidle4	:	in	std_logic	:=	'0';
		rxelecidle5	:	in	std_logic	:=	'0';
		rxelecidle6	:	in	std_logic	:=	'0';
		rxelecidle7	:	in	std_logic	:=	'0';
		rxfreqlocked0	:	in	std_logic	:=	'0';
		rxfreqlocked1	:	in	std_logic	:=	'0';
		rxfreqlocked2	:	in	std_logic	:=	'0';
		rxfreqlocked3	:	in	std_logic	:=	'0';
		rxfreqlocked4	:	in	std_logic	:=	'0';
		rxfreqlocked5	:	in	std_logic	:=	'0';
		rxfreqlocked6	:	in	std_logic	:=	'0';
		rxfreqlocked7	:	in	std_logic	:=	'0';
		rxstatus0	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus1	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus2	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus3	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus4	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus5	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus6	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus7	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxsynchd0	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd1	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd2	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd3	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd4	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd5	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd6	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd7	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxvalid0	:	in	std_logic	:=	'0';
		rxvalid1	:	in	std_logic	:=	'0';
		rxvalid2	:	in	std_logic	:=	'0';
		rxvalid3	:	in	std_logic	:=	'0';
		rxvalid4	:	in	std_logic	:=	'0';
		rxvalid5	:	in	std_logic	:=	'0';
		rxvalid6	:	in	std_logic	:=	'0';
		rxvalid7	:	in	std_logic	:=	'0';
		scan_mode_n	:	in	std_logic	:=	'0';
		scan_shift_n	:	in	std_logic	:=	'0';
		sw_ctmod	:	in	std_logic_vector(1 downto 0)	:=	"00";
		swdn_in	:	in	std_logic_vector(2 downto 0)	:=	"000";
		swup_in	:	in	std_logic_vector(6 downto 0)	:=	"0000000";
		test_in_1_hip	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		test_in_hip	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		test_pl_dbg_eqin	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		tx_cred_cons_select	:	in	std_logic	:=	'0';
		tx_cred_fc_sel	:	in	std_logic_vector(1 downto 0)	:=	"00";
		tx_lcff_pll_lock0	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock1	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock2	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock3	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock4	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock5	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock6	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock7	:	in	std_logic	:=	'0';
		tx_st_data	:	in	std_logic_vector(255 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		tx_st_empty	:	in	std_logic_vector(1 downto 0)	:=	"00";
		tx_st_eop	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		tx_st_err	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		tx_st_parity	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		tx_st_sop	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		tx_st_valid	:	in	std_logic	:=	'0';
		user_mode	:	in	std_logic	:=	'0';
		sta_hd_altpe3_hip_core_top_hd_altpe3_hip_core_u_clkmux_core_clk_cnt_reg_0_0_Q	:	out	std_logic	:=	'0';
		sta_hd_altpe3_hip_core_top_hd_altpe3_hip_core_u_clkmux_core_clk_cnt_reg_1_0_Q	:	out	std_logic	:=	'0';
		sta_hd_altpe3_hip_core_top_hd_altpe3_hip_core_u_clkmux_core_clk_cnt_reg_2_0_Q	:	out	std_logic	:=	'0';
		app_inta_ack	:	out	std_logic	:=	'0';
		app_msi_ack	:	out	std_logic	:=	'0';
		avmm_readdata	:	out	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		cfg_par_err	:	out	std_logic	:=	'0';
		core_clk_out	:	out	std_logic	:=	'0';
		cseb_addr	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		cseb_addr_parity	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		cseb_be	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		cseb_is_shadow	:	out	std_logic	:=	'0';
		cseb_rden	:	out	std_logic	:=	'0';
		cseb_wrdata	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		cseb_wrdata_parity	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		cseb_wren	:	out	std_logic	:=	'0';
		cseb_wrresp_req	:	out	std_logic	:=	'0';
		csr_dout	:	out	std_logic	:=	'0';
		csr_out	:	out	std_logic	:=	'0';
		csr_pipe_out	:	out	std_logic	:=	'0';
		current_coeff0	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff1	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff2	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff3	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff4	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff5	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff6	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff7	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_rxpreset0	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset1	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset2	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset3	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset4	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset5	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset6	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset7	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_speed	:	out	std_logic_vector(1 downto 0)	:=	"00";
		cvp_clk	:	out	std_logic	:=	'0';
		cvp_config	:	out	std_logic	:=	'0';
		cvp_data	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		cvp_full_config	:	out	std_logic	:=	'0';
		cvp_start_xfer	:	out	std_logic	:=	'0';
		dl_up	:	out	std_logic	:=	'0';
		dlup_exit	:	out	std_logic	:=	'0';
		eidle_infer_sel0	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel1	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel2	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel3	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel4	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel5	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel6	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel7	:	out	std_logic_vector(2 downto 0)	:=	"000";
		ev_128ns	:	out	std_logic	:=	'0';
		ev_1us	:	out	std_logic	:=	'0';
		flr_sts	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n0	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n1	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n2	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n3	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n4	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n5	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n6	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n7	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n0	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n1	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n2	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n3	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n4	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n5	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n6	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n7	:	out	std_logic	:=	'0';
		hotrst_exit	:	out	std_logic	:=	'0';
		int_status	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		k_hip_pcs_chnl_en	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		k_hrc_chnl_en	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		k_hrc_chnl_txpll_master_cgb_rst_en	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		k_hrc_chnl_txpll_rst_en	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		l2_exit	:	out	std_logic	:=	'0';
		lane_act	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		lmi_ack	:	out	std_logic	:=	'0';
		lmi_dout	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		ltssm_state	:	out	std_logic_vector(4 downto 0)	:=	"00000";
		mem_rscout_rcv_bot	:	out	std_logic	:=	'0';
		mem_rscout_rcv_top	:	out	std_logic	:=	'0';
		mem_rscout_rtry	:	out	std_logic	:=	'0';
		pld_clk_in_use	:	out	std_logic	:=	'0';
		pld_gp_ctrl	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		pm_exit_d0_req	:	out	std_logic	:=	'0';
		pme_to_sr	:	out	std_logic	:=	'0';
		powerdown0	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown1	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown2	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown3	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown4	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown5	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown6	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown7	:	out	std_logic_vector(1 downto 0)	:=	"00";
		r2c_unc_ecc	:	out	std_logic	:=	'0';
		rate0	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate1	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate2	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate3	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate4	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate5	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate6	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate7	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate_ctrl	:	out	std_logic_vector(1 downto 0)	:=	"00";
		reserved_clk_out	:	out	std_logic	:=	'0';
		reserved_out	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		reset_status	:	out	std_logic	:=	'0';
		retry_corr_ecc	:	out	std_logic	:=	'0';
		retry_unc_ecc	:	out	std_logic	:=	'0';
		rx_corr_ecc	:	out	std_logic	:=	'0';
		rx_cred_status	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		rx_par_err	:	out	std_logic	:=	'0';
		rx_pcs_rst_n0	:	out	std_logic	:=	'0';
		rx_pcs_rst_n1	:	out	std_logic	:=	'0';
		rx_pcs_rst_n2	:	out	std_logic	:=	'0';
		rx_pcs_rst_n3	:	out	std_logic	:=	'0';
		rx_pcs_rst_n4	:	out	std_logic	:=	'0';
		rx_pcs_rst_n5	:	out	std_logic	:=	'0';
		rx_pcs_rst_n6	:	out	std_logic	:=	'0';
		rx_pcs_rst_n7	:	out	std_logic	:=	'0';
		rx_pma_rstb0	:	out	std_logic	:=	'0';
		rx_pma_rstb1	:	out	std_logic	:=	'0';
		rx_pma_rstb2	:	out	std_logic	:=	'0';
		rx_pma_rstb3	:	out	std_logic	:=	'0';
		rx_pma_rstb4	:	out	std_logic	:=	'0';
		rx_pma_rstb5	:	out	std_logic	:=	'0';
		rx_pma_rstb6	:	out	std_logic	:=	'0';
		rx_pma_rstb7	:	out	std_logic	:=	'0';
		rx_st_bardec1	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		rx_st_bardec2	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		rx_st_be	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rx_st_data	:	out	std_logic_vector(255 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		rx_st_empty	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rx_st_eop	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		rx_st_err	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		rx_st_parity	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rx_st_sop	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		rx_st_valid	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		rxfc_cplbuf_ovf	:	out	std_logic	:=	'0';
		rxfc_cplovf_tag	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		rxpolarity0	:	out	std_logic	:=	'0';
		rxpolarity1	:	out	std_logic	:=	'0';
		rxpolarity2	:	out	std_logic	:=	'0';
		rxpolarity3	:	out	std_logic	:=	'0';
		rxpolarity4	:	out	std_logic	:=	'0';
		rxpolarity5	:	out	std_logic	:=	'0';
		rxpolarity6	:	out	std_logic	:=	'0';
		rxpolarity7	:	out	std_logic	:=	'0';
		serr_out	:	out	std_logic	:=	'0';
		swdn_out	:	out	std_logic_vector(6 downto 0)	:=	"0000000";
		swup_out	:	out	std_logic_vector(2 downto 0)	:=	"000";
		test_fref_clk	:	out	std_logic	:=	'0';
		test_out_1_hip	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		test_out_hip	:	out	std_logic_vector(255 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		tl_cfg_add	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		tl_cfg_ctl	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		tl_cfg_sts	:	out	std_logic_vector(52 downto 0)	:=	"00000000000000000000000000000000000000000000000000000";
		tl_cfg_sts_wr	:	out	std_logic	:=	'0';
		tx_cred_data_fc	:	out	std_logic_vector(11 downto 0)	:=	"000000000000";
		tx_cred_fc_hip_cons	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		tx_cred_fc_infinite	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		tx_cred_hdr_fc	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		tx_deemph0	:	out	std_logic	:=	'0';
		tx_deemph1	:	out	std_logic	:=	'0';
		tx_deemph2	:	out	std_logic	:=	'0';
		tx_deemph3	:	out	std_logic	:=	'0';
		tx_deemph4	:	out	std_logic	:=	'0';
		tx_deemph5	:	out	std_logic	:=	'0';
		tx_deemph6	:	out	std_logic	:=	'0';
		tx_deemph7	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb0	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb1	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb2	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb3	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb4	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb5	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb6	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb7	:	out	std_logic	:=	'0';
		tx_margin0	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin1	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin2	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin3	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin4	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin5	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin6	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin7	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_par_err	:	out	std_logic_vector(1 downto 0)	:=	"00";
		tx_pcs_rst_n0	:	out	std_logic	:=	'0';
		tx_pcs_rst_n1	:	out	std_logic	:=	'0';
		tx_pcs_rst_n2	:	out	std_logic	:=	'0';
		tx_pcs_rst_n3	:	out	std_logic	:=	'0';
		tx_pcs_rst_n4	:	out	std_logic	:=	'0';
		tx_pcs_rst_n5	:	out	std_logic	:=	'0';
		tx_pcs_rst_n6	:	out	std_logic	:=	'0';
		tx_pcs_rst_n7	:	out	std_logic	:=	'0';
		tx_pma_syncp0	:	out	std_logic	:=	'0';
		tx_pma_syncp1	:	out	std_logic	:=	'0';
		tx_pma_syncp2	:	out	std_logic	:=	'0';
		tx_pma_syncp3	:	out	std_logic	:=	'0';
		tx_pma_syncp4	:	out	std_logic	:=	'0';
		tx_pma_syncp5	:	out	std_logic	:=	'0';
		tx_pma_syncp6	:	out	std_logic	:=	'0';
		tx_pma_syncp7	:	out	std_logic	:=	'0';
		tx_st_ready	:	out	std_logic	:=	'0';
		txblkst0	:	out	std_logic	:=	'0';
		txblkst1	:	out	std_logic	:=	'0';
		txblkst2	:	out	std_logic	:=	'0';
		txblkst3	:	out	std_logic	:=	'0';
		txblkst4	:	out	std_logic	:=	'0';
		txblkst5	:	out	std_logic	:=	'0';
		txblkst6	:	out	std_logic	:=	'0';
		txblkst7	:	out	std_logic	:=	'0';
		txcompl0	:	out	std_logic	:=	'0';
		txcompl1	:	out	std_logic	:=	'0';
		txcompl2	:	out	std_logic	:=	'0';
		txcompl3	:	out	std_logic	:=	'0';
		txcompl4	:	out	std_logic	:=	'0';
		txcompl5	:	out	std_logic	:=	'0';
		txcompl6	:	out	std_logic	:=	'0';
		txcompl7	:	out	std_logic	:=	'0';
		txdata0	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata1	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata2	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata3	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata4	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata5	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata6	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata7	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdatak0	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak1	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak2	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak3	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak4	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak5	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak6	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak7	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdataskip0	:	out	std_logic	:=	'0';
		txdataskip1	:	out	std_logic	:=	'0';
		txdataskip2	:	out	std_logic	:=	'0';
		txdataskip3	:	out	std_logic	:=	'0';
		txdataskip4	:	out	std_logic	:=	'0';
		txdataskip5	:	out	std_logic	:=	'0';
		txdataskip6	:	out	std_logic	:=	'0';
		txdataskip7	:	out	std_logic	:=	'0';
		txdetectrx0	:	out	std_logic	:=	'0';
		txdetectrx1	:	out	std_logic	:=	'0';
		txdetectrx2	:	out	std_logic	:=	'0';
		txdetectrx3	:	out	std_logic	:=	'0';
		txdetectrx4	:	out	std_logic	:=	'0';
		txdetectrx5	:	out	std_logic	:=	'0';
		txdetectrx6	:	out	std_logic	:=	'0';
		txdetectrx7	:	out	std_logic	:=	'0';
		txelecidle0	:	out	std_logic	:=	'0';
		txelecidle1	:	out	std_logic	:=	'0';
		txelecidle2	:	out	std_logic	:=	'0';
		txelecidle3	:	out	std_logic	:=	'0';
		txelecidle4	:	out	std_logic	:=	'0';
		txelecidle5	:	out	std_logic	:=	'0';
		txelecidle6	:	out	std_logic	:=	'0';
		txelecidle7	:	out	std_logic	:=	'0';
		txst_prot_err	:	out	std_logic	:=	'0';
		txswing0	:	out	std_logic	:=	'0';
		txswing1	:	out	std_logic	:=	'0';
		txswing2	:	out	std_logic	:=	'0';
		txswing3	:	out	std_logic	:=	'0';
		txswing4	:	out	std_logic	:=	'0';
		txswing5	:	out	std_logic	:=	'0';
		txswing6	:	out	std_logic	:=	'0';
		txswing7	:	out	std_logic	:=	'0';
		txsynchd0	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd1	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd2	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd3	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd4	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd5	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd6	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd7	:	out	std_logic_vector(1 downto 0)	:=	"00";
		wake_oen	:	out	std_logic	:=	'0'
	);
end twentynm_hssi_gen3_x8_pcie_hip;

architecture behavior of twentynm_hssi_gen3_x8_pcie_hip	is

constant acknack_base_int	:	integer	:=	bin2int(acknack_base);
constant arb_upfc_30us_counter_int	:	integer	:=	bin2int(arb_upfc_30us_counter);
constant bar0_size_mask_int	:	integer	:=	bin2int(bar0_size_mask);
constant bar1_size_mask_int	:	integer	:=	bin2int(bar1_size_mask);
constant bar2_size_mask_int	:	integer	:=	bin2int(bar2_size_mask);
constant bar3_size_mask_int	:	integer	:=	bin2int(bar3_size_mask);
constant bar4_size_mask_int	:	integer	:=	bin2int(bar4_size_mask);
constant bar5_size_mask_int	:	integer	:=	bin2int(bar5_size_mask);
constant cdc_dummy_insert_limit_int	:	integer	:=	bin2int(cdc_dummy_insert_limit);
constant class_code_int	:	integer	:=	bin2int(class_code);
constant device_id_int	:	integer	:=	bin2int(device_id);
constant device_number_int	:	integer	:=	bin2int(device_number);
constant diffclock_nfts_count_int	:	integer	:=	bin2int(diffclock_nfts_count);
constant ei_delay_powerdown_count_int	:	integer	:=	bin2int(ei_delay_powerdown_count);
constant eie_before_nfts_count_int	:	integer	:=	bin2int(eie_before_nfts_count);
constant endpoint_l0_latency_int	:	integer	:=	bin2int(endpoint_l0_latency);
constant endpoint_l1_latency_int	:	integer	:=	bin2int(endpoint_l1_latency);
constant eql_rq_int_en_number_int	:	integer	:=	bin2int(eql_rq_int_en_number);
constant fc_init_timer_int	:	integer	:=	bin2int(fc_init_timer);
constant flow_control_timeout_count_int	:	integer	:=	bin2int(flow_control_timeout_count);
constant flow_control_update_count_int	:	integer	:=	bin2int(flow_control_update_count);
constant g3_dn_rx_hint_eqlz_0_int	:	integer	:=	bin2int(g3_dn_rx_hint_eqlz_0);
constant g3_dn_rx_hint_eqlz_1_int	:	integer	:=	bin2int(g3_dn_rx_hint_eqlz_1);
constant g3_dn_rx_hint_eqlz_2_int	:	integer	:=	bin2int(g3_dn_rx_hint_eqlz_2);
constant g3_dn_rx_hint_eqlz_3_int	:	integer	:=	bin2int(g3_dn_rx_hint_eqlz_3);
constant g3_dn_rx_hint_eqlz_4_int	:	integer	:=	bin2int(g3_dn_rx_hint_eqlz_4);
constant g3_dn_rx_hint_eqlz_5_int	:	integer	:=	bin2int(g3_dn_rx_hint_eqlz_5);
constant g3_dn_rx_hint_eqlz_6_int	:	integer	:=	bin2int(g3_dn_rx_hint_eqlz_6);
constant g3_dn_rx_hint_eqlz_7_int	:	integer	:=	bin2int(g3_dn_rx_hint_eqlz_7);
constant g3_dn_tx_preset_eqlz_0_int	:	integer	:=	bin2int(g3_dn_tx_preset_eqlz_0);
constant g3_dn_tx_preset_eqlz_1_int	:	integer	:=	bin2int(g3_dn_tx_preset_eqlz_1);
constant g3_dn_tx_preset_eqlz_2_int	:	integer	:=	bin2int(g3_dn_tx_preset_eqlz_2);
constant g3_dn_tx_preset_eqlz_3_int	:	integer	:=	bin2int(g3_dn_tx_preset_eqlz_3);
constant g3_dn_tx_preset_eqlz_4_int	:	integer	:=	bin2int(g3_dn_tx_preset_eqlz_4);
constant g3_dn_tx_preset_eqlz_5_int	:	integer	:=	bin2int(g3_dn_tx_preset_eqlz_5);
constant g3_dn_tx_preset_eqlz_6_int	:	integer	:=	bin2int(g3_dn_tx_preset_eqlz_6);
constant g3_dn_tx_preset_eqlz_7_int	:	integer	:=	bin2int(g3_dn_tx_preset_eqlz_7);
constant g3_up_rx_hint_eqlz_0_int	:	integer	:=	bin2int(g3_up_rx_hint_eqlz_0);
constant g3_up_rx_hint_eqlz_1_int	:	integer	:=	bin2int(g3_up_rx_hint_eqlz_1);
constant g3_up_rx_hint_eqlz_2_int	:	integer	:=	bin2int(g3_up_rx_hint_eqlz_2);
constant g3_up_rx_hint_eqlz_3_int	:	integer	:=	bin2int(g3_up_rx_hint_eqlz_3);
constant g3_up_rx_hint_eqlz_4_int	:	integer	:=	bin2int(g3_up_rx_hint_eqlz_4);
constant g3_up_rx_hint_eqlz_5_int	:	integer	:=	bin2int(g3_up_rx_hint_eqlz_5);
constant g3_up_rx_hint_eqlz_6_int	:	integer	:=	bin2int(g3_up_rx_hint_eqlz_6);
constant g3_up_rx_hint_eqlz_7_int	:	integer	:=	bin2int(g3_up_rx_hint_eqlz_7);
constant g3_up_tx_preset_eqlz_0_int	:	integer	:=	bin2int(g3_up_tx_preset_eqlz_0);
constant g3_up_tx_preset_eqlz_1_int	:	integer	:=	bin2int(g3_up_tx_preset_eqlz_1);
constant g3_up_tx_preset_eqlz_2_int	:	integer	:=	bin2int(g3_up_tx_preset_eqlz_2);
constant g3_up_tx_preset_eqlz_3_int	:	integer	:=	bin2int(g3_up_tx_preset_eqlz_3);
constant g3_up_tx_preset_eqlz_4_int	:	integer	:=	bin2int(g3_up_tx_preset_eqlz_4);
constant g3_up_tx_preset_eqlz_5_int	:	integer	:=	bin2int(g3_up_tx_preset_eqlz_5);
constant g3_up_tx_preset_eqlz_6_int	:	integer	:=	bin2int(g3_up_tx_preset_eqlz_6);
constant g3_up_tx_preset_eqlz_7_int	:	integer	:=	bin2int(g3_up_tx_preset_eqlz_7);
constant gen2_diffclock_nfts_count_int	:	integer	:=	bin2int(gen2_diffclock_nfts_count);
constant gen2_sameclock_nfts_count_int	:	integer	:=	bin2int(gen2_sameclock_nfts_count);
constant gen3_coeff_1_int	:	integer	:=	bin2int(gen3_coeff_1);
constant gen3_coeff_10_int	:	integer	:=	bin2int(gen3_coeff_10);
constant gen3_coeff_10_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_10_ber_meas);
constant gen3_coeff_10_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_10_nxtber_less);
constant gen3_coeff_10_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_10_nxtber_more);
constant gen3_coeff_10_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_10_preset_hint);
constant gen3_coeff_10_reqber_int	:	integer	:=	bin2int(gen3_coeff_10_reqber);
constant gen3_coeff_11_int	:	integer	:=	bin2int(gen3_coeff_11);
constant gen3_coeff_11_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_11_ber_meas);
constant gen3_coeff_11_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_11_nxtber_less);
constant gen3_coeff_11_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_11_nxtber_more);
constant gen3_coeff_11_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_11_preset_hint);
constant gen3_coeff_11_reqber_int	:	integer	:=	bin2int(gen3_coeff_11_reqber);
constant gen3_coeff_12_int	:	integer	:=	bin2int(gen3_coeff_12);
constant gen3_coeff_12_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_12_ber_meas);
constant gen3_coeff_12_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_12_nxtber_less);
constant gen3_coeff_12_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_12_nxtber_more);
constant gen3_coeff_12_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_12_preset_hint);
constant gen3_coeff_12_reqber_int	:	integer	:=	bin2int(gen3_coeff_12_reqber);
constant gen3_coeff_13_int	:	integer	:=	bin2int(gen3_coeff_13);
constant gen3_coeff_13_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_13_ber_meas);
constant gen3_coeff_13_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_13_nxtber_less);
constant gen3_coeff_13_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_13_nxtber_more);
constant gen3_coeff_13_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_13_preset_hint);
constant gen3_coeff_13_reqber_int	:	integer	:=	bin2int(gen3_coeff_13_reqber);
constant gen3_coeff_14_int	:	integer	:=	bin2int(gen3_coeff_14);
constant gen3_coeff_14_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_14_ber_meas);
constant gen3_coeff_14_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_14_nxtber_less);
constant gen3_coeff_14_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_14_nxtber_more);
constant gen3_coeff_14_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_14_preset_hint);
constant gen3_coeff_14_reqber_int	:	integer	:=	bin2int(gen3_coeff_14_reqber);
constant gen3_coeff_15_int	:	integer	:=	bin2int(gen3_coeff_15);
constant gen3_coeff_15_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_15_ber_meas);
constant gen3_coeff_15_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_15_nxtber_less);
constant gen3_coeff_15_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_15_nxtber_more);
constant gen3_coeff_15_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_15_preset_hint);
constant gen3_coeff_15_reqber_int	:	integer	:=	bin2int(gen3_coeff_15_reqber);
constant gen3_coeff_16_int	:	integer	:=	bin2int(gen3_coeff_16);
constant gen3_coeff_16_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_16_ber_meas);
constant gen3_coeff_16_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_16_nxtber_less);
constant gen3_coeff_16_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_16_nxtber_more);
constant gen3_coeff_16_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_16_preset_hint);
constant gen3_coeff_16_reqber_int	:	integer	:=	bin2int(gen3_coeff_16_reqber);
constant gen3_coeff_17_int	:	integer	:=	bin2int(gen3_coeff_17);
constant gen3_coeff_17_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_17_ber_meas);
constant gen3_coeff_17_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_17_nxtber_less);
constant gen3_coeff_17_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_17_nxtber_more);
constant gen3_coeff_17_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_17_preset_hint);
constant gen3_coeff_17_reqber_int	:	integer	:=	bin2int(gen3_coeff_17_reqber);
constant gen3_coeff_18_int	:	integer	:=	bin2int(gen3_coeff_18);
constant gen3_coeff_18_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_18_ber_meas);
constant gen3_coeff_18_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_18_nxtber_less);
constant gen3_coeff_18_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_18_nxtber_more);
constant gen3_coeff_18_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_18_preset_hint);
constant gen3_coeff_18_reqber_int	:	integer	:=	bin2int(gen3_coeff_18_reqber);
constant gen3_coeff_19_int	:	integer	:=	bin2int(gen3_coeff_19);
constant gen3_coeff_19_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_19_ber_meas);
constant gen3_coeff_19_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_19_nxtber_less);
constant gen3_coeff_19_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_19_nxtber_more);
constant gen3_coeff_19_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_19_preset_hint);
constant gen3_coeff_19_reqber_int	:	integer	:=	bin2int(gen3_coeff_19_reqber);
constant gen3_coeff_1_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_1_ber_meas);
constant gen3_coeff_1_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_1_nxtber_less);
constant gen3_coeff_1_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_1_nxtber_more);
constant gen3_coeff_1_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_1_preset_hint);
constant gen3_coeff_1_reqber_int	:	integer	:=	bin2int(gen3_coeff_1_reqber);
constant gen3_coeff_2_int	:	integer	:=	bin2int(gen3_coeff_2);
constant gen3_coeff_20_int	:	integer	:=	bin2int(gen3_coeff_20);
constant gen3_coeff_20_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_20_ber_meas);
constant gen3_coeff_20_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_20_nxtber_less);
constant gen3_coeff_20_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_20_nxtber_more);
constant gen3_coeff_20_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_20_preset_hint);
constant gen3_coeff_20_reqber_int	:	integer	:=	bin2int(gen3_coeff_20_reqber);
constant gen3_coeff_21_int	:	integer	:=	bin2int(gen3_coeff_21);
constant gen3_coeff_21_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_21_ber_meas);
constant gen3_coeff_21_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_21_nxtber_less);
constant gen3_coeff_21_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_21_nxtber_more);
constant gen3_coeff_21_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_21_preset_hint);
constant gen3_coeff_21_reqber_int	:	integer	:=	bin2int(gen3_coeff_21_reqber);
constant gen3_coeff_22_int	:	integer	:=	bin2int(gen3_coeff_22);
constant gen3_coeff_22_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_22_ber_meas);
constant gen3_coeff_22_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_22_nxtber_less);
constant gen3_coeff_22_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_22_nxtber_more);
constant gen3_coeff_22_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_22_preset_hint);
constant gen3_coeff_22_reqber_int	:	integer	:=	bin2int(gen3_coeff_22_reqber);
constant gen3_coeff_23_int	:	integer	:=	bin2int(gen3_coeff_23);
constant gen3_coeff_23_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_23_ber_meas);
constant gen3_coeff_23_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_23_nxtber_less);
constant gen3_coeff_23_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_23_nxtber_more);
constant gen3_coeff_23_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_23_preset_hint);
constant gen3_coeff_23_reqber_int	:	integer	:=	bin2int(gen3_coeff_23_reqber);
constant gen3_coeff_24_int	:	integer	:=	bin2int(gen3_coeff_24);
constant gen3_coeff_24_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_24_ber_meas);
constant gen3_coeff_24_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_24_nxtber_less);
constant gen3_coeff_24_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_24_nxtber_more);
constant gen3_coeff_24_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_24_preset_hint);
constant gen3_coeff_24_reqber_int	:	integer	:=	bin2int(gen3_coeff_24_reqber);
constant gen3_coeff_2_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_2_ber_meas);
constant gen3_coeff_2_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_2_nxtber_less);
constant gen3_coeff_2_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_2_nxtber_more);
constant gen3_coeff_2_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_2_preset_hint);
constant gen3_coeff_2_reqber_int	:	integer	:=	bin2int(gen3_coeff_2_reqber);
constant gen3_coeff_3_int	:	integer	:=	bin2int(gen3_coeff_3);
constant gen3_coeff_3_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_3_ber_meas);
constant gen3_coeff_3_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_3_nxtber_less);
constant gen3_coeff_3_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_3_nxtber_more);
constant gen3_coeff_3_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_3_preset_hint);
constant gen3_coeff_3_reqber_int	:	integer	:=	bin2int(gen3_coeff_3_reqber);
constant gen3_coeff_4_int	:	integer	:=	bin2int(gen3_coeff_4);
constant gen3_coeff_4_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_4_ber_meas);
constant gen3_coeff_4_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_4_nxtber_less);
constant gen3_coeff_4_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_4_nxtber_more);
constant gen3_coeff_4_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_4_preset_hint);
constant gen3_coeff_4_reqber_int	:	integer	:=	bin2int(gen3_coeff_4_reqber);
constant gen3_coeff_5_int	:	integer	:=	bin2int(gen3_coeff_5);
constant gen3_coeff_5_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_5_ber_meas);
constant gen3_coeff_5_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_5_nxtber_less);
constant gen3_coeff_5_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_5_nxtber_more);
constant gen3_coeff_5_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_5_preset_hint);
constant gen3_coeff_5_reqber_int	:	integer	:=	bin2int(gen3_coeff_5_reqber);
constant gen3_coeff_6_int	:	integer	:=	bin2int(gen3_coeff_6);
constant gen3_coeff_6_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_6_ber_meas);
constant gen3_coeff_6_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_6_nxtber_less);
constant gen3_coeff_6_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_6_nxtber_more);
constant gen3_coeff_6_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_6_preset_hint);
constant gen3_coeff_6_reqber_int	:	integer	:=	bin2int(gen3_coeff_6_reqber);
constant gen3_coeff_7_int	:	integer	:=	bin2int(gen3_coeff_7);
constant gen3_coeff_7_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_7_ber_meas);
constant gen3_coeff_7_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_7_nxtber_less);
constant gen3_coeff_7_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_7_nxtber_more);
constant gen3_coeff_7_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_7_preset_hint);
constant gen3_coeff_7_reqber_int	:	integer	:=	bin2int(gen3_coeff_7_reqber);
constant gen3_coeff_8_int	:	integer	:=	bin2int(gen3_coeff_8);
constant gen3_coeff_8_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_8_ber_meas);
constant gen3_coeff_8_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_8_nxtber_less);
constant gen3_coeff_8_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_8_nxtber_more);
constant gen3_coeff_8_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_8_preset_hint);
constant gen3_coeff_8_reqber_int	:	integer	:=	bin2int(gen3_coeff_8_reqber);
constant gen3_coeff_9_int	:	integer	:=	bin2int(gen3_coeff_9);
constant gen3_coeff_9_ber_meas_int	:	integer	:=	bin2int(gen3_coeff_9_ber_meas);
constant gen3_coeff_9_nxtber_less_int	:	integer	:=	bin2int(gen3_coeff_9_nxtber_less);
constant gen3_coeff_9_nxtber_more_int	:	integer	:=	bin2int(gen3_coeff_9_nxtber_more);
constant gen3_coeff_9_preset_hint_int	:	integer	:=	bin2int(gen3_coeff_9_preset_hint);
constant gen3_coeff_9_reqber_int	:	integer	:=	bin2int(gen3_coeff_9_reqber);
constant gen3_coeff_delay_count_int	:	integer	:=	bin2int(gen3_coeff_delay_count);
constant gen3_diffclock_nfts_count_int	:	integer	:=	bin2int(gen3_diffclock_nfts_count);
constant gen3_full_swing_int	:	integer	:=	bin2int(gen3_full_swing);
constant gen3_low_freq_int	:	integer	:=	bin2int(gen3_low_freq);
constant gen3_preset_coeff_1_int	:	integer	:=	bin2int(gen3_preset_coeff_1);
constant gen3_preset_coeff_10_int	:	integer	:=	bin2int(gen3_preset_coeff_10);
constant gen3_preset_coeff_11_int	:	integer	:=	bin2int(gen3_preset_coeff_11);
constant gen3_preset_coeff_2_int	:	integer	:=	bin2int(gen3_preset_coeff_2);
constant gen3_preset_coeff_3_int	:	integer	:=	bin2int(gen3_preset_coeff_3);
constant gen3_preset_coeff_4_int	:	integer	:=	bin2int(gen3_preset_coeff_4);
constant gen3_preset_coeff_5_int	:	integer	:=	bin2int(gen3_preset_coeff_5);
constant gen3_preset_coeff_6_int	:	integer	:=	bin2int(gen3_preset_coeff_6);
constant gen3_preset_coeff_7_int	:	integer	:=	bin2int(gen3_preset_coeff_7);
constant gen3_preset_coeff_8_int	:	integer	:=	bin2int(gen3_preset_coeff_8);
constant gen3_preset_coeff_9_int	:	integer	:=	bin2int(gen3_preset_coeff_9);
constant gen3_rxfreqlock_counter_int	:	integer	:=	bin2int(gen3_rxfreqlock_counter);
constant gen3_sameclock_nfts_count_int	:	integer	:=	bin2int(gen3_sameclock_nfts_count);
constant hip_ac_pwr_clk_freq_in_hz_int	:	integer	:=	bin2int(hip_ac_pwr_clk_freq_in_hz);
constant hip_ac_pwr_uw_per_mhz_int	:	integer	:=	bin2int(hip_ac_pwr_uw_per_mhz);
constant hip_base_address_int	:	integer	:=	bin2int(hip_base_address);
constant hot_plug_support_int	:	integer	:=	bin2int(hot_plug_support);
constant indicator_int	:	integer	:=	bin2int(indicator);
constant ko_compl_data_int	:	integer	:=	bin2int(ko_compl_data);
constant ko_compl_header_int	:	integer	:=	bin2int(ko_compl_header);
constant l01_entry_latency_int	:	integer	:=	bin2int(l01_entry_latency);
constant l0_exit_latency_diffclock_int	:	integer	:=	bin2int(l0_exit_latency_diffclock);
constant l0_exit_latency_sameclock_int	:	integer	:=	bin2int(l0_exit_latency_sameclock);
constant l1_exit_latency_diffclock_int	:	integer	:=	bin2int(l1_exit_latency_diffclock);
constant l1_exit_latency_sameclock_int	:	integer	:=	bin2int(l1_exit_latency_sameclock);
constant maximum_current_int	:	integer	:=	bin2int(maximum_current);
constant millisecond_cycle_count_int	:	integer	:=	bin2int(millisecond_cycle_count);
constant msix_pba_bir_int	:	integer	:=	bin2int(msix_pba_bir);
constant msix_pba_offset_int	:	integer	:=	bin2int(msix_pba_offset);
constant msix_table_bir_int	:	integer	:=	bin2int(msix_table_bir);
constant msix_table_offset_int	:	integer	:=	bin2int(msix_table_offset);
constant msix_table_size_int	:	integer	:=	bin2int(msix_table_size);
constant port_link_number_int	:	integer	:=	bin2int(port_link_number);
constant retry_buffer_last_active_address_int	:	integer	:=	bin2int(retry_buffer_last_active_address);
constant revision_id_int	:	integer	:=	bin2int(revision_id);
constant rp_bug_fix_pri_sec_stat_reg_int	:	integer	:=	bin2int(rp_bug_fix_pri_sec_stat_reg);
constant rpltim_base_int	:	integer	:=	bin2int(rpltim_base);
constant rstctrl_1ms_count_fref_clk_int	:	integer	:=	bin2int(rstctrl_1ms_count_fref_clk);
constant rstctrl_1us_count_fref_clk_int	:	integer	:=	bin2int(rstctrl_1us_count_fref_clk);
constant rstctrl_timer_a_int	:	integer	:=	bin2int(rstctrl_timer_a);
constant rstctrl_timer_b_int	:	integer	:=	bin2int(rstctrl_timer_b);
constant rstctrl_timer_c_int	:	integer	:=	bin2int(rstctrl_timer_c);
constant rstctrl_timer_d_int	:	integer	:=	bin2int(rstctrl_timer_d);
constant rstctrl_timer_e_int	:	integer	:=	bin2int(rstctrl_timer_e);
constant rstctrl_timer_f_int	:	integer	:=	bin2int(rstctrl_timer_f);
constant rstctrl_timer_g_int	:	integer	:=	bin2int(rstctrl_timer_g);
constant rstctrl_timer_h_int	:	integer	:=	bin2int(rstctrl_timer_h);
constant rstctrl_timer_i_int	:	integer	:=	bin2int(rstctrl_timer_i);
constant rstctrl_timer_j_int	:	integer	:=	bin2int(rstctrl_timer_j);
constant rx_buffer_fc_protect_int	:	integer	:=	bin2int(rx_buffer_fc_protect);
constant rx_buffer_protect_int	:	integer	:=	bin2int(rx_buffer_protect);
constant rx_cdc_almost_empty_int	:	integer	:=	bin2int(rx_cdc_almost_empty);
constant rx_cdc_almost_full_int	:	integer	:=	bin2int(rx_cdc_almost_full);
constant rx_l0s_count_idl_int	:	integer	:=	bin2int(rx_l0s_count_idl);
constant rx_ptr0_nonposted_dpram_max_int	:	integer	:=	bin2int(rx_ptr0_nonposted_dpram_max);
constant rx_ptr0_nonposted_dpram_min_int	:	integer	:=	bin2int(rx_ptr0_nonposted_dpram_min);
constant rx_ptr0_posted_dpram_max_int	:	integer	:=	bin2int(rx_ptr0_posted_dpram_max);
constant rx_ptr0_posted_dpram_min_int	:	integer	:=	bin2int(rx_ptr0_posted_dpram_min);
constant sameclock_nfts_count_int	:	integer	:=	bin2int(sameclock_nfts_count);
constant skp_os_gen3_count_int	:	integer	:=	bin2int(skp_os_gen3_count);
constant skp_os_schedule_count_int	:	integer	:=	bin2int(skp_os_schedule_count);
constant slot_number_int	:	integer	:=	bin2int(slot_number);
constant slot_power_limit_int	:	integer	:=	bin2int(slot_power_limit);
constant slot_power_scale_int	:	integer	:=	bin2int(slot_power_scale);
constant ssid_int	:	integer	:=	bin2int(ssid);
constant ssvid_int	:	integer	:=	bin2int(ssvid);
constant subsystem_device_id_int	:	integer	:=	bin2int(subsystem_device_id);
constant subsystem_vendor_id_int	:	integer	:=	bin2int(subsystem_vendor_id);
constant tx_cdc_almost_empty_int	:	integer	:=	bin2int(tx_cdc_almost_empty);
constant tx_cdc_almost_full_int	:	integer	:=	bin2int(tx_cdc_almost_full);
constant tx_swing_int	:	integer	:=	bin2int(tx_swing);
constant txdl_fair_arbiter_counter_int	:	integer	:=	bin2int(txdl_fair_arbiter_counter);
constant user_id_int	:	integer	:=	bin2int(user_id);
constant vc0_rx_flow_ctrl_compl_data_int	:	integer	:=	bin2int(vc0_rx_flow_ctrl_compl_data);
constant vc0_rx_flow_ctrl_compl_header_int	:	integer	:=	bin2int(vc0_rx_flow_ctrl_compl_header);
constant vc0_rx_flow_ctrl_nonposted_data_int	:	integer	:=	bin2int(vc0_rx_flow_ctrl_nonposted_data);
constant vc0_rx_flow_ctrl_nonposted_header_int	:	integer	:=	bin2int(vc0_rx_flow_ctrl_nonposted_header);
constant vc0_rx_flow_ctrl_posted_data_int	:	integer	:=	bin2int(vc0_rx_flow_ctrl_posted_data);
constant vc0_rx_flow_ctrl_posted_header_int	:	integer	:=	bin2int(vc0_rx_flow_ctrl_posted_header);
constant vendor_id_int	:	integer	:=	bin2int(vendor_id);
constant vsec_cap_int	:	integer	:=	bin2int(vsec_cap);
constant vsec_id_int	:	integer	:=	bin2int(vsec_id);



component	twentynm_hssi_gen3_x8_pcie_hip_encrypted
	generic (
		-- Architecture parameters
		acknack_base	:	integer	:=	0;
		acknack_set	:	string	:=	"false";
		advance_error_reporting	:	string	:=	"disable";
		app_interface_width	:	string	:=	"avst_64bit";
		arb_upfc_30us_counter	:	integer	:=	0;
		arb_upfc_30us_en	:	string	:=	"enable";
		aspm_config_management	:	string	:=	"true";
		aspm_patch_disable	:	string	:=	"enable_both";
		ast_width_rx	:	string	:=	"rx_64";
		ast_width_tx	:	string	:=	"tx_64";
		atomic_malformed	:	string	:=	"false";
		atomic_op_completer_32bit	:	string	:=	"false";
		atomic_op_completer_64bit	:	string	:=	"false";
		atomic_op_routing	:	string	:=	"false";
		auto_msg_drop_enable	:	string	:=	"false";
		avmm_cvp_inter_sel_csr_ctrl	:	string	:=	"disable";
		avmm_dprio_broadcast_en_csr_ctrl	:	string	:=	"disable";
		avmm_force_inter_sel_csr_ctrl	:	string	:=	"disable";
		avmm_power_iso_en_csr_ctrl	:	string	:=	"disable";
		bar0_size_mask	:	integer	:=	268435455;
		bar0_type	:	string	:=	"bar0_64bit_prefetch_mem";
		bar1_size_mask	:	integer	:=	0;
		bar1_type	:	string	:=	"bar1_disable";
		bar2_size_mask	:	integer	:=	0;
		bar2_type	:	string	:=	"bar2_disable";
		bar3_size_mask	:	integer	:=	0;
		bar3_type	:	string	:=	"bar3_disable";
		bar4_size_mask	:	integer	:=	0;
		bar4_type	:	string	:=	"bar4_disable";
		bar5_size_mask	:	integer	:=	0;
		bar5_type	:	string	:=	"bar5_disable";
		base_counter_sel	:	string	:=	"count_clk_62p5";
		bist_memory_settings	:	string	:=	"000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		bridge_port_ssid_support	:	string	:=	"false";
		bridge_port_vga_enable	:	string	:=	"false";
		bypass_cdc	:	string	:=	"false";
		bypass_clk_switch	:	string	:=	"false";
		bypass_tl	:	string	:=	"false";
		capab_rate_rxcfg_en	:	string	:=	"disable";
		cas_completer_128bit	:	string	:=	"false";
		cdc_clk_relation	:	string	:=	"plesiochronous";
		cdc_dummy_insert_limit	:	integer	:=	11;
		cfg_parchk_ena	:	string	:=	"disable";
		cfgbp_req_recov_disable	:	string	:=	"false";
		class_code	:	integer	:=	16711680;
		clock_pwr_management	:	string	:=	"false";
		completion_timeout	:	string	:=	"abcd";
		core_clk_divider	:	string	:=	"div_1";
		core_clk_freq_mhz	:	string	:=	"core_clk_250mhz";
		core_clk_out_sel	:	string	:=	"core_clk_out_div_1";
		core_clk_sel	:	string	:=	"pld_clk";
		core_clk_source	:	string	:=	"pll_fixed_clk";
		cseb_bar_match_checking	:	string	:=	"enable";
		cseb_config_bypass	:	string	:=	"disable";
		cseb_cpl_status_during_cvp	:	string	:=	"completer_abort";
		cseb_cpl_tag_checking	:	string	:=	"enable";
		cseb_disable_auto_crs	:	string	:=	"false";
		cseb_extend_pci	:	string	:=	"false";
		cseb_extend_pcie	:	string	:=	"false";
		cseb_min_error_checking	:	string	:=	"false";
		cseb_route_to_avl_rx_st	:	string	:=	"cseb";
		cseb_temp_busy_crs	:	string	:=	"completer_abort_tmp_busy";
		cvp_clk_reset	:	string	:=	"false";
		cvp_data_compressed	:	string	:=	"false";
		cvp_data_encrypted	:	string	:=	"false";
		cvp_enable	:	string	:=	"cvp_dis";
		cvp_mode_reset	:	string	:=	"false";
		cvp_rate_sel	:	string	:=	"full_rate";
		d0_pme	:	string	:=	"false";
		d1_pme	:	string	:=	"false";
		d1_support	:	string	:=	"false";
		d2_pme	:	string	:=	"false";
		d2_support	:	string	:=	"false";
		d3_cold_pme	:	string	:=	"false";
		d3_hot_pme	:	string	:=	"false";
		data_pack_rx	:	string	:=	"disable";
		deemphasis_enable	:	string	:=	"false";
		deskew_comma	:	string	:=	"skp_eieos_deskw";
		device_id	:	integer	:=	57345;
		device_number	:	integer	:=	0;
		device_specific_init	:	string	:=	"false";
		dft_clock_obsrv_en	:	string	:=	"disable";
		dft_clock_obsrv_sel	:	string	:=	"dft_pclk";
		diffclock_nfts_count	:	integer	:=	0;
		dis_cplovf	:	string	:=	"disable";
		dis_paritychk	:	string	:=	"enable";
		disable_link_x2_support	:	string	:=	"false";
		disable_snoop_packet	:	string	:=	"false";
		dl_tx_check_parity_edb	:	string	:=	"disable";
		dll_active_report_support	:	string	:=	"false";
		early_dl_up	:	string	:=	"true";
		eco_fb332688_dis	:	string	:=	"true";
		ecrc_check_capable	:	string	:=	"true";
		ecrc_gen_capable	:	string	:=	"true";
		egress_block_err_report_ena	:	string	:=	"false";
		ei_delay_powerdown_count	:	integer	:=	10;
		eie_before_nfts_count	:	integer	:=	4;
		electromech_interlock	:	string	:=	"false";
		en_ieiupdatefc	:	string	:=	"false";
		en_lane_errchk	:	string	:=	"false";
		en_phystatus_dly	:	string	:=	"false";
		ena_ido_cpl	:	string	:=	"false";
		ena_ido_req	:	string	:=	"false";
		enable_adapter_half_rate_mode	:	string	:=	"false";
		enable_ch01_pclk_out	:	string	:=	"pclk_ch0";
		enable_ch0_pclk_out	:	string	:=	"pclk_ch01";
		enable_completion_timeout_disable	:	string	:=	"true";
		enable_directed_spd_chng	:	string	:=	"false";
		enable_function_msix_support	:	string	:=	"true";
		enable_l0s_aspm	:	string	:=	"false";
		enable_l1_aspm	:	string	:=	"false";
		enable_rx_buffer_checking	:	string	:=	"false";
		enable_rx_reordering	:	string	:=	"true";
		enable_slot_register	:	string	:=	"false";
		endpoint_l0_latency	:	integer	:=	0;
		endpoint_l1_latency	:	integer	:=	0;
		eql_rq_int_en_number	:	integer	:=	0;
		errmgt_fcpe_patch_dis	:	string	:=	"enable";
		errmgt_fep_patch_dis	:	string	:=	"enable";
		expansion_base_address_register	:	string	:=	"00000000000000000000000000000000";
		extend_tag_field	:	string	:=	"false";
		extended_format_field	:	string	:=	"true";
		extended_tag_reset	:	string	:=	"false";
		fc_init_timer	:	integer	:=	1024;
		flow_control_timeout_count	:	integer	:=	200;
		flow_control_update_count	:	integer	:=	30;
		flr_capability	:	string	:=	"true";
		force_dis_to_det	:	string	:=	"false";
		force_gen1_dis	:	string	:=	"false";
		force_tx_coeff_preset_lpbk	:	string	:=	"false";
		frame_err_patch_dis	:	string	:=	"enable";
		func_mode	:	string	:=	"disable";
		g3_bypass_equlz	:	string	:=	"false";
		g3_coeff_done_tmout	:	string	:=	"enable";
		g3_deskew_char	:	string	:=	"default_sdsos";
		g3_dis_be_frm_err	:	string	:=	"false";
		g3_dn_rx_hint_eqlz_0	:	integer	:=	0;
		g3_dn_rx_hint_eqlz_1	:	integer	:=	0;
		g3_dn_rx_hint_eqlz_2	:	integer	:=	0;
		g3_dn_rx_hint_eqlz_3	:	integer	:=	0;
		g3_dn_rx_hint_eqlz_4	:	integer	:=	0;
		g3_dn_rx_hint_eqlz_5	:	integer	:=	0;
		g3_dn_rx_hint_eqlz_6	:	integer	:=	0;
		g3_dn_rx_hint_eqlz_7	:	integer	:=	0;
		g3_dn_tx_preset_eqlz_0	:	integer	:=	0;
		g3_dn_tx_preset_eqlz_1	:	integer	:=	0;
		g3_dn_tx_preset_eqlz_2	:	integer	:=	0;
		g3_dn_tx_preset_eqlz_3	:	integer	:=	0;
		g3_dn_tx_preset_eqlz_4	:	integer	:=	0;
		g3_dn_tx_preset_eqlz_5	:	integer	:=	0;
		g3_dn_tx_preset_eqlz_6	:	integer	:=	0;
		g3_dn_tx_preset_eqlz_7	:	integer	:=	0;
		g3_force_ber_max	:	string	:=	"false";
		g3_force_ber_min	:	string	:=	"false";
		g3_lnk_trn_rx_ts	:	string	:=	"false";
		g3_ltssm_eq_dbg	:	string	:=	"false";
		g3_ltssm_rec_dbg	:	string	:=	"false";
		g3_pause_ltssm_rec_en	:	string	:=	"disable";
		g3_quiesce_guarant	:	string	:=	"false";
		g3_redo_equlz_dis	:	string	:=	"false";
		g3_redo_equlz_en	:	string	:=	"false";
		g3_up_rx_hint_eqlz_0	:	integer	:=	0;
		g3_up_rx_hint_eqlz_1	:	integer	:=	0;
		g3_up_rx_hint_eqlz_2	:	integer	:=	0;
		g3_up_rx_hint_eqlz_3	:	integer	:=	0;
		g3_up_rx_hint_eqlz_4	:	integer	:=	0;
		g3_up_rx_hint_eqlz_5	:	integer	:=	0;
		g3_up_rx_hint_eqlz_6	:	integer	:=	0;
		g3_up_rx_hint_eqlz_7	:	integer	:=	0;
		g3_up_tx_preset_eqlz_0	:	integer	:=	0;
		g3_up_tx_preset_eqlz_1	:	integer	:=	0;
		g3_up_tx_preset_eqlz_2	:	integer	:=	0;
		g3_up_tx_preset_eqlz_3	:	integer	:=	0;
		g3_up_tx_preset_eqlz_4	:	integer	:=	0;
		g3_up_tx_preset_eqlz_5	:	integer	:=	0;
		g3_up_tx_preset_eqlz_6	:	integer	:=	0;
		g3_up_tx_preset_eqlz_7	:	integer	:=	0;
		gen123_lane_rate_mode	:	string	:=	"gen1_rate";
		gen2_diffclock_nfts_count	:	integer	:=	255;
		gen2_pma_pll_usage	:	string	:=	"not_applicaple";
		gen2_sameclock_nfts_count	:	integer	:=	255;
		gen3_coeff_1	:	integer	:=	4;
		gen3_coeff_10	:	integer	:=	7;
		gen3_coeff_10_ber_meas	:	integer	:=	2;
		gen3_coeff_10_nxtber_less	:	integer	:=	15;
		gen3_coeff_10_nxtber_more	:	integer	:=	10;
		gen3_coeff_10_preset_hint	:	integer	:=	3;
		gen3_coeff_10_reqber	:	integer	:=	8;
		gen3_coeff_10_sel	:	string	:=	"preset_10";
		gen3_coeff_11	:	integer	:=	7;
		gen3_coeff_11_ber_meas	:	integer	:=	2;
		gen3_coeff_11_nxtber_less	:	integer	:=	15;
		gen3_coeff_11_nxtber_more	:	integer	:=	15;
		gen3_coeff_11_preset_hint	:	integer	:=	4;
		gen3_coeff_11_reqber	:	integer	:=	8;
		gen3_coeff_11_sel	:	string	:=	"preset_11";
		gen3_coeff_12	:	integer	:=	7;
		gen3_coeff_12_ber_meas	:	integer	:=	2;
		gen3_coeff_12_nxtber_less	:	integer	:=	15;
		gen3_coeff_12_nxtber_more	:	integer	:=	15;
		gen3_coeff_12_preset_hint	:	integer	:=	2;
		gen3_coeff_12_reqber	:	integer	:=	8;
		gen3_coeff_12_sel	:	string	:=	"preset_12";
		gen3_coeff_13	:	integer	:=	4;
		gen3_coeff_13_ber_meas	:	integer	:=	2;
		gen3_coeff_13_nxtber_less	:	integer	:=	13;
		gen3_coeff_13_nxtber_more	:	integer	:=	1;
		gen3_coeff_13_preset_hint	:	integer	:=	4;
		gen3_coeff_13_reqber	:	integer	:=	8;
		gen3_coeff_13_sel	:	string	:=	"preset_13";
		gen3_coeff_14	:	integer	:=	4;
		gen3_coeff_14_ber_meas	:	integer	:=	2;
		gen3_coeff_14_nxtber_less	:	integer	:=	15;
		gen3_coeff_14_nxtber_more	:	integer	:=	2;
		gen3_coeff_14_preset_hint	:	integer	:=	0;
		gen3_coeff_14_reqber	:	integer	:=	8;
		gen3_coeff_14_sel	:	string	:=	"preset_14";
		gen3_coeff_15	:	integer	:=	0;
		gen3_coeff_15_ber_meas	:	integer	:=	2;
		gen3_coeff_15_nxtber_less	:	integer	:=	0;
		gen3_coeff_15_nxtber_more	:	integer	:=	0;
		gen3_coeff_15_preset_hint	:	integer	:=	0;
		gen3_coeff_15_reqber	:	integer	:=	0;
		gen3_coeff_15_sel	:	string	:=	"coeff_15";
		gen3_coeff_16	:	integer	:=	0;
		gen3_coeff_16_ber_meas	:	integer	:=	0;
		gen3_coeff_16_nxtber_less	:	integer	:=	0;
		gen3_coeff_16_nxtber_more	:	integer	:=	0;
		gen3_coeff_16_preset_hint	:	integer	:=	0;
		gen3_coeff_16_reqber	:	integer	:=	0;
		gen3_coeff_16_sel	:	string	:=	"coeff_16";
		gen3_coeff_17	:	integer	:=	0;
		gen3_coeff_17_ber_meas	:	integer	:=	0;
		gen3_coeff_17_nxtber_less	:	integer	:=	0;
		gen3_coeff_17_nxtber_more	:	integer	:=	0;
		gen3_coeff_17_preset_hint	:	integer	:=	0;
		gen3_coeff_17_reqber	:	integer	:=	0;
		gen3_coeff_17_sel	:	string	:=	"coeff_17";
		gen3_coeff_18	:	integer	:=	0;
		gen3_coeff_18_ber_meas	:	integer	:=	0;
		gen3_coeff_18_nxtber_less	:	integer	:=	0;
		gen3_coeff_18_nxtber_more	:	integer	:=	0;
		gen3_coeff_18_preset_hint	:	integer	:=	0;
		gen3_coeff_18_reqber	:	integer	:=	0;
		gen3_coeff_18_sel	:	string	:=	"coeff_18";
		gen3_coeff_19	:	integer	:=	0;
		gen3_coeff_19_ber_meas	:	integer	:=	0;
		gen3_coeff_19_nxtber_less	:	integer	:=	0;
		gen3_coeff_19_nxtber_more	:	integer	:=	0;
		gen3_coeff_19_preset_hint	:	integer	:=	0;
		gen3_coeff_19_reqber	:	integer	:=	0;
		gen3_coeff_19_sel	:	string	:=	"coeff_19";
		gen3_coeff_1_ber_meas	:	integer	:=	2;
		gen3_coeff_1_nxtber_less	:	integer	:=	12;
		gen3_coeff_1_nxtber_more	:	integer	:=	6;
		gen3_coeff_1_preset_hint	:	integer	:=	2;
		gen3_coeff_1_reqber	:	integer	:=	8;
		gen3_coeff_1_sel	:	string	:=	"preset_1";
		gen3_coeff_2	:	integer	:=	1;
		gen3_coeff_20	:	integer	:=	0;
		gen3_coeff_20_ber_meas	:	integer	:=	0;
		gen3_coeff_20_nxtber_less	:	integer	:=	0;
		gen3_coeff_20_nxtber_more	:	integer	:=	0;
		gen3_coeff_20_preset_hint	:	integer	:=	0;
		gen3_coeff_20_reqber	:	integer	:=	0;
		gen3_coeff_20_sel	:	string	:=	"coeff_20";
		gen3_coeff_21	:	integer	:=	0;
		gen3_coeff_21_ber_meas	:	integer	:=	0;
		gen3_coeff_21_nxtber_less	:	integer	:=	0;
		gen3_coeff_21_nxtber_more	:	integer	:=	0;
		gen3_coeff_21_preset_hint	:	integer	:=	0;
		gen3_coeff_21_reqber	:	integer	:=	0;
		gen3_coeff_21_sel	:	string	:=	"coeff_21";
		gen3_coeff_22	:	integer	:=	0;
		gen3_coeff_22_ber_meas	:	integer	:=	0;
		gen3_coeff_22_nxtber_less	:	integer	:=	0;
		gen3_coeff_22_nxtber_more	:	integer	:=	0;
		gen3_coeff_22_preset_hint	:	integer	:=	0;
		gen3_coeff_22_reqber	:	integer	:=	0;
		gen3_coeff_22_sel	:	string	:=	"coeff_22";
		gen3_coeff_23	:	integer	:=	0;
		gen3_coeff_23_ber_meas	:	integer	:=	0;
		gen3_coeff_23_nxtber_less	:	integer	:=	0;
		gen3_coeff_23_nxtber_more	:	integer	:=	0;
		gen3_coeff_23_preset_hint	:	integer	:=	0;
		gen3_coeff_23_reqber	:	integer	:=	0;
		gen3_coeff_23_sel	:	string	:=	"coeff_23";
		gen3_coeff_24	:	integer	:=	0;
		gen3_coeff_24_ber_meas	:	integer	:=	0;
		gen3_coeff_24_nxtber_less	:	integer	:=	0;
		gen3_coeff_24_nxtber_more	:	integer	:=	0;
		gen3_coeff_24_preset_hint	:	integer	:=	0;
		gen3_coeff_24_reqber	:	integer	:=	0;
		gen3_coeff_24_sel	:	string	:=	"coeff_24";
		gen3_coeff_2_ber_meas	:	integer	:=	2;
		gen3_coeff_2_nxtber_less	:	integer	:=	2;
		gen3_coeff_2_nxtber_more	:	integer	:=	4;
		gen3_coeff_2_preset_hint	:	integer	:=	4;
		gen3_coeff_2_reqber	:	integer	:=	8;
		gen3_coeff_2_sel	:	string	:=	"preset_2";
		gen3_coeff_3	:	integer	:=	1;
		gen3_coeff_3_ber_meas	:	integer	:=	2;
		gen3_coeff_3_nxtber_less	:	integer	:=	15;
		gen3_coeff_3_nxtber_more	:	integer	:=	3;
		gen3_coeff_3_preset_hint	:	integer	:=	0;
		gen3_coeff_3_reqber	:	integer	:=	8;
		gen3_coeff_3_sel	:	string	:=	"preset_3";
		gen3_coeff_4	:	integer	:=	0;
		gen3_coeff_4_ber_meas	:	integer	:=	2;
		gen3_coeff_4_nxtber_less	:	integer	:=	15;
		gen3_coeff_4_nxtber_more	:	integer	:=	4;
		gen3_coeff_4_preset_hint	:	integer	:=	0;
		gen3_coeff_4_reqber	:	integer	:=	8;
		gen3_coeff_4_sel	:	string	:=	"preset_4";
		gen3_coeff_5	:	integer	:=	0;
		gen3_coeff_5_ber_meas	:	integer	:=	2;
		gen3_coeff_5_nxtber_less	:	integer	:=	15;
		gen3_coeff_5_nxtber_more	:	integer	:=	5;
		gen3_coeff_5_preset_hint	:	integer	:=	4;
		gen3_coeff_5_reqber	:	integer	:=	8;
		gen3_coeff_5_sel	:	string	:=	"preset_5";
		gen3_coeff_6	:	integer	:=	7;
		gen3_coeff_6_ber_meas	:	integer	:=	2;
		gen3_coeff_6_nxtber_less	:	integer	:=	15;
		gen3_coeff_6_nxtber_more	:	integer	:=	15;
		gen3_coeff_6_preset_hint	:	integer	:=	4;
		gen3_coeff_6_reqber	:	integer	:=	8;
		gen3_coeff_6_sel	:	string	:=	"preset_6";
		gen3_coeff_7	:	integer	:=	1;
		gen3_coeff_7_ber_meas	:	integer	:=	2;
		gen3_coeff_7_nxtber_less	:	integer	:=	1;
		gen3_coeff_7_nxtber_more	:	integer	:=	7;
		gen3_coeff_7_preset_hint	:	integer	:=	2;
		gen3_coeff_7_reqber	:	integer	:=	8;
		gen3_coeff_7_sel	:	string	:=	"preset_7";
		gen3_coeff_8	:	integer	:=	0;
		gen3_coeff_8_ber_meas	:	integer	:=	2;
		gen3_coeff_8_nxtber_less	:	integer	:=	4;
		gen3_coeff_8_nxtber_more	:	integer	:=	8;
		gen3_coeff_8_preset_hint	:	integer	:=	2;
		gen3_coeff_8_reqber	:	integer	:=	8;
		gen3_coeff_8_sel	:	string	:=	"preset_8";
		gen3_coeff_9	:	integer	:=	0;
		gen3_coeff_9_ber_meas	:	integer	:=	2;
		gen3_coeff_9_nxtber_less	:	integer	:=	11;
		gen3_coeff_9_nxtber_more	:	integer	:=	9;
		gen3_coeff_9_preset_hint	:	integer	:=	3;
		gen3_coeff_9_reqber	:	integer	:=	8;
		gen3_coeff_9_sel	:	string	:=	"preset_9";
		gen3_coeff_delay_count	:	integer	:=	125;
		gen3_coeff_errchk	:	string	:=	"enable";
		gen3_dcbal_en	:	string	:=	"true";
		gen3_diffclock_nfts_count	:	integer	:=	128;
		gen3_force_local_coeff	:	string	:=	"false";
		gen3_full_swing	:	integer	:=	63;
		gen3_half_swing	:	string	:=	"false";
		gen3_low_freq	:	integer	:=	1;
		gen3_paritychk	:	string	:=	"enable";
		gen3_pl_framing_err_dis	:	string	:=	"enable";
		gen3_preset_coeff_1	:	integer	:=	3402;
		gen3_preset_coeff_10	:	integer	:=	48384;
		gen3_preset_coeff_11	:	integer	:=	124992;
		gen3_preset_coeff_2	:	integer	:=	3339;
		gen3_preset_coeff_3	:	integer	:=	3213;
		gen3_preset_coeff_4	:	integer	:=	3528;
		gen3_preset_coeff_5	:	integer	:=	4032;
		gen3_preset_coeff_6	:	integer	:=	28224;
		gen3_preset_coeff_7	:	integer	:=	36288;
		gen3_preset_coeff_8	:	integer	:=	27405;
		gen3_preset_coeff_9	:	integer	:=	35784;
		gen3_reset_eieos_cnt_bit	:	string	:=	"false";
		gen3_rxfreqlock_counter	:	integer	:=	0;
		gen3_sameclock_nfts_count	:	integer	:=	128;
		gen3_scrdscr_bypass	:	string	:=	"false";
		gen3_skip_ph2_ph3	:	string	:=	"false";
		hard_reset_bypass	:	string	:=	"false";
		hard_rst_sig_chnl_en	:	string	:=	"disable_hrc_sig";
		hard_rst_tx_pll_rst_chnl_en	:	string	:=	"disable_hrc_txpll_rst";
		hip_ac_pwr_clk_freq_in_hz	:	integer	:=	0;
		hip_ac_pwr_uw_per_mhz	:	integer	:=	0;
		hip_base_address	:	integer	:=	0;
		hip_clock_dis	:	string	:=	"enable_hip_clk";
		hip_hard_reset	:	string	:=	"enable";
		hip_pcs_sig_chnl_en	:	string	:=	"disable_hip_pcs_sig";
		hot_plug_support	:	integer	:=	0;
		hrc_chnl_txpll_master_cgb_rst_select	:	string	:=	"disable_master_cgb_sel";
		hrdrstctrl_en	:	string	:=	"hrdrstctrl_dis";
		iei_enable_settings	:	string	:=	"gen3gen2_infei_infsd_gen1_infei_sd";
		indicator	:	integer	:=	7;
		intel_id_access	:	string	:=	"false";
		interrupt_pin	:	string	:=	"inta";
		io_window_addr_width	:	string	:=	"window_32_bit";
		jtag_id	:	string	:=	"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		ko_compl_data	:	integer	:=	0;
		ko_compl_header	:	integer	:=	0;
		l01_entry_latency	:	integer	:=	31;
		l0_exit_latency_diffclock	:	integer	:=	6;
		l0_exit_latency_sameclock	:	integer	:=	6;
		l0s_adj_rply_timer_dis	:	string	:=	"enable";
		l1_exit_latency_diffclock	:	integer	:=	0;
		l1_exit_latency_sameclock	:	integer	:=	0;
		l2_async_logic	:	string	:=	"enable";
		lane_mask	:	string	:=	"ln_mask_x4";
		lane_rate	:	string	:=	"gen1";
		link_width	:	string	:=	"x1";
		lmi_hold_off_cfg_timer_en	:	string	:=	"disable";
		low_priority_vc	:	string	:=	"single_vc_low_pr";
		ltr_mechanism	:	string	:=	"false";
		ltssm_1ms_timeout	:	string	:=	"disable";
		ltssm_freqlocked_check	:	string	:=	"disable";
		malformed_tlp_truncate_en	:	string	:=	"disable";
		max_link_width	:	string	:=	"x4_link_width";
		max_payload_size	:	string	:=	"payload_512";
		maximum_current	:	integer	:=	0;
		millisecond_cycle_count	:	integer	:=	0;
		msi_64bit_addressing_capable	:	string	:=	"true";
		msi_masking_capable	:	string	:=	"false";
		msi_multi_message_capable	:	string	:=	"count_4";
		msi_support	:	string	:=	"true";
		msix_pba_bir	:	integer	:=	0;
		msix_pba_offset	:	integer	:=	0;
		msix_table_bir	:	integer	:=	0;
		msix_table_offset	:	integer	:=	0;
		msix_table_size	:	integer	:=	0;
		national_inst_thru_enhance	:	string	:=	"true";
		no_command_completed	:	string	:=	"true";
		no_soft_reset	:	string	:=	"false";
		not_use_k_gbl_bits	:	string	:=	"not_used_k_gbl";
		operating_voltage	:	string	:=	"standard";
		pcie_base_spec	:	string	:=	"pcie_2p1";
		pcie_mode	:	string	:=	"shared_mode";
		pcie_spec_1p0_compliance	:	string	:=	"spec_1p1";
		pcie_spec_version	:	string	:=	"v2";
		pclk_out_sel	:	string	:=	"pclk";
		pld_in_use_reg	:	string	:=	"false";
		pm_latency_patch_dis	:	string	:=	"enable";
		pm_txdl_patch_dis	:	string	:=	"enable";
		pme_clock	:	string	:=	"false";
		port_link_number	:	integer	:=	1;
		port_type	:	string	:=	"native_ep";
		powerdown_mode	:	string	:=	"powerup";
		prefetchable_mem_window_addr_width	:	string	:=	"prefetch_32";
		r2c_mask_easy	:	string	:=	"false";
		r2c_mask_enable	:	string	:=	"false";
		rec_frqlk_mon_en	:	string	:=	"disable";
		register_pipe_signals	:	string	:=	"true";
		retry_buffer_last_active_address	:	integer	:=	1023;
		retry_buffer_memory_settings	:	string	:=	"000000000000000000000000000000000000";
		retry_ecc_corr_mask_dis	:	string	:=	"enable";
		revision_id	:	integer	:=	1;
		role_based_error_reporting	:	string	:=	"false";
		rp_bug_fix_pri_sec_stat_reg	:	integer	:=	127;
		rpltim_base	:	integer	:=	0;
		rpltim_set	:	string	:=	"false";
		rstctl_ltssm_dis	:	string	:=	"false";
		rstctrl_1ms_count_fref_clk	:	integer	:=	62500;
		rstctrl_1us_count_fref_clk	:	integer	:=	63;
		rstctrl_altpe3_crst_n_inv	:	string	:=	"false";
		rstctrl_altpe3_rst_n_inv	:	string	:=	"false";
		rstctrl_altpe3_srst_n_inv	:	string	:=	"false";
		rstctrl_chnl_cal_done_select	:	string	:=	"not_active_chnl_cal_done";
		rstctrl_debug_en	:	string	:=	"false";
		rstctrl_force_inactive_rst	:	string	:=	"false";
		rstctrl_fref_clk_select	:	string	:=	"ch0_sel";
		rstctrl_hard_block_enable	:	string	:=	"hard_rst_ctl";
		rstctrl_hip_ep	:	string	:=	"hip_ep";
		rstctrl_mask_tx_pll_lock_select	:	string	:=	"not_active_mask_tx_pll_lock";
		rstctrl_perst_enable	:	string	:=	"level";
		rstctrl_perstn_select	:	string	:=	"perstn_pin";
		rstctrl_pld_clr	:	string	:=	"false";
		rstctrl_pll_cal_done_select	:	string	:=	"not_active_pll_cal_done";
		rstctrl_rx_pcs_rst_n_inv	:	string	:=	"false";
		rstctrl_rx_pcs_rst_n_select	:	string	:=	"not_active_rx_pcs_rst";
		rstctrl_rx_pll_freq_lock_select	:	string	:=	"not_active_rx_pll_f_lock";
		rstctrl_rx_pll_lock_select	:	string	:=	"not_active_rx_pll_lock";
		rstctrl_rx_pma_rstb_inv	:	string	:=	"false";
		rstctrl_rx_pma_rstb_select	:	string	:=	"not_active_rx_pma_rstb";
		rstctrl_timer_a	:	integer	:=	10;
		rstctrl_timer_a_type	:	string	:=	"a_timer_milli_secs";
		rstctrl_timer_b	:	integer	:=	10;
		rstctrl_timer_b_type	:	string	:=	"b_timer_milli_secs";
		rstctrl_timer_c	:	integer	:=	10;
		rstctrl_timer_c_type	:	string	:=	"c_timer_milli_secs";
		rstctrl_timer_d	:	integer	:=	20;
		rstctrl_timer_d_type	:	string	:=	"d_timer_milli_secs";
		rstctrl_timer_e	:	integer	:=	1;
		rstctrl_timer_e_type	:	string	:=	"e_timer_milli_secs";
		rstctrl_timer_f	:	integer	:=	10;
		rstctrl_timer_f_type	:	string	:=	"f_timer_milli_secs";
		rstctrl_timer_g	:	integer	:=	10;
		rstctrl_timer_g_type	:	string	:=	"g_timer_milli_secs";
		rstctrl_timer_h	:	integer	:=	4;
		rstctrl_timer_h_type	:	string	:=	"h_timer_milli_secs";
		rstctrl_timer_i	:	integer	:=	20;
		rstctrl_timer_i_type	:	string	:=	"i_timer_milli_secs";
		rstctrl_timer_j	:	integer	:=	20;
		rstctrl_timer_j_type	:	string	:=	"j_timer_milli_secs";
		rstctrl_tx_lcff_pll_lock_select	:	string	:=	"not_active_lcff_pll_lock";
		rstctrl_tx_lcff_pll_rstb_select	:	string	:=	"not_active_lcff_pll_rstb";
		rstctrl_tx_pcs_rst_n_inv	:	string	:=	"false";
		rstctrl_tx_pcs_rst_n_select	:	string	:=	"not_active_tx_pcs_rst";
		rstctrl_tx_pma_rstb_inv	:	string	:=	"false";
		rstctrl_tx_pma_syncp_inv	:	string	:=	"false";
		rstctrl_tx_pma_syncp_select	:	string	:=	"not_active_tx_pma_syncp";
		rx_ast_parity	:	string	:=	"disable";
		rx_buffer_credit_alloc	:	string	:=	"balance";
		rx_buffer_fc_protect	:	integer	:=	68;
		rx_buffer_protect	:	integer	:=	68;
		rx_cdc_almost_empty	:	integer	:=	3;
		rx_cdc_almost_full	:	integer	:=	12;
		rx_cred_ctl_param	:	string	:=	"disable";
		rx_ei_l0s	:	string	:=	"disable";
		rx_l0s_count_idl	:	integer	:=	0;
		rx_ptr0_nonposted_dpram_max	:	integer	:=	0;
		rx_ptr0_nonposted_dpram_min	:	integer	:=	0;
		rx_ptr0_posted_dpram_max	:	integer	:=	0;
		rx_ptr0_posted_dpram_min	:	integer	:=	0;
		rx_runt_patch_dis	:	string	:=	"enable";
		rx_sop_ctrl	:	string	:=	"rx_sop_boundary_64";
		rx_trunc_patch_dis	:	string	:=	"enable";
		rx_use_prst	:	string	:=	"false";
		rx_use_prst_ep	:	string	:=	"true";
		rxbuf_ecc_corr_mask_dis	:	string	:=	"enable";
		rxdl_bad_sop_eop_filter_dis	:	string	:=	"rxdlbug1_enable_both";
		rxdl_bad_tlp_patch_dis	:	string	:=	"rxdlbug2_enable_both";
		rxdl_lcrc_patch_dis	:	string	:=	"rxdlbug3_enable_both";
		sameclock_nfts_count	:	integer	:=	0;
		sel_enable_pcs_rx_fifo_err	:	string	:=	"disable_sel";
		silicon_rev	:	string	:=	"20nm5es";
		sim_mode	:	string	:=	"disable";
		simple_ro_fifo_control_en	:	string	:=	"disable";
		single_rx_detect	:	string	:=	"detect_all_lanes";
		skp_os_gen3_count	:	integer	:=	0;
		skp_os_schedule_count	:	integer	:=	0;
		slot_number	:	integer	:=	0;
		slot_power_limit	:	integer	:=	0;
		slot_power_scale	:	integer	:=	0;
		slotclk_cfg	:	string	:=	"static_slotclkcfgon";
		ssid	:	integer	:=	0;
		ssvid	:	integer	:=	0;
		subsystem_device_id	:	integer	:=	57345;
		subsystem_vendor_id	:	integer	:=	4466;
		sup_mode	:	string	:=	"user_mode";
		surprise_down_error_support	:	string	:=	"false";
		tl_cfg_div	:	string	:=	"cfg_clk_div_7";
		tl_tx_check_parity_msg	:	string	:=	"disable";
		tph_completer	:	string	:=	"false";
		tx_ast_parity	:	string	:=	"disable";
		tx_cdc_almost_empty	:	integer	:=	5;
		tx_cdc_almost_full	:	integer	:=	12;
		tx_sop_ctrl	:	string	:=	"boundary_64";
		tx_swing	:	integer	:=	0;
		txdl_fair_arbiter_counter	:	integer	:=	0;
		txdl_fair_arbiter_en	:	string	:=	"enable";
		txrate_adv	:	string	:=	"capability";
		uc_calibration_en	:	string	:=	"uc_calibration_dis";
		use_aer	:	string	:=	"false";
		use_crc_forwarding	:	string	:=	"false";
		user_id	:	integer	:=	0;
		vc0_clk_enable	:	string	:=	"true";
		vc0_rx_buffer_memory_settings	:	string	:=	"000000000000000000000000000000000000";
		vc0_rx_flow_ctrl_compl_data	:	integer	:=	448;
		vc0_rx_flow_ctrl_compl_header	:	integer	:=	112;
		vc0_rx_flow_ctrl_nonposted_data	:	integer	:=	0;
		vc0_rx_flow_ctrl_nonposted_header	:	integer	:=	54;
		vc0_rx_flow_ctrl_posted_data	:	integer	:=	360;
		vc0_rx_flow_ctrl_posted_header	:	integer	:=	50;
		vc1_clk_enable	:	string	:=	"false";
		vc_arbitration	:	string	:=	"single_vc_arb";
		vc_enable	:	string	:=	"single_vc";
		vendor_id	:	integer	:=	4466;
		vsec_cap	:	integer	:=	0;
		vsec_id	:	integer	:=	4466;
		wrong_device_id	:	string	:=	"disable"
	);
	port (
		-- Architecture ports
		aer_msi_num	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		app_int_err	:	in	std_logic_vector(1 downto 0)	:=	"00";
		app_inta_sts	:	in	std_logic	:=	'0';
		app_msi_num	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		app_msi_req	:	in	std_logic	:=	'0';
		app_msi_tc	:	in	std_logic_vector(2 downto 0)	:=	"000";
		atpg_los_en_n	:	in	std_logic	:=	'0';
		avmm_address	:	in	std_logic_vector(9 downto 0)	:=	"0000000000";
		avmm_byte_en	:	in	std_logic_vector(1 downto 0)	:=	"00";
		avmm_clk	:	in	std_logic	:=	'0';
		avmm_read	:	in	std_logic	:=	'0';
		avmm_rst_n	:	in	std_logic	:=	'0';
		avmm_write	:	in	std_logic	:=	'0';
		avmm_writedata	:	in	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		bist_scanen	:	in	std_logic	:=	'0';
		bist_scanin	:	in	std_logic	:=	'0';
		bisten_rcv_n	:	in	std_logic	:=	'0';
		bisten_rpl_n	:	in	std_logic	:=	'0';
		bistmode_n	:	in	std_logic	:=	'0';
		cfg_link2csr_pld	:	in	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		cfg_prmbus_pld	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		chnl_cal_done0	:	in	std_logic	:=	'0';
		chnl_cal_done1	:	in	std_logic	:=	'0';
		chnl_cal_done2	:	in	std_logic	:=	'0';
		chnl_cal_done3	:	in	std_logic	:=	'0';
		chnl_cal_done4	:	in	std_logic	:=	'0';
		chnl_cal_done5	:	in	std_logic	:=	'0';
		chnl_cal_done6	:	in	std_logic	:=	'0';
		chnl_cal_done7	:	in	std_logic	:=	'0';
		core_clk_in	:	in	std_logic	:=	'0';
		core_crst	:	in	std_logic	:=	'0';
		core_por	:	in	std_logic	:=	'0';
		core_rst	:	in	std_logic	:=	'0';
		core_srst	:	in	std_logic	:=	'0';
		cpl_err	:	in	std_logic_vector(6 downto 0)	:=	"0000000";
		cpl_pending	:	in	std_logic	:=	'0';
		cseb_rddata	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		cseb_rddata_parity	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		cseb_rdresponse	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		cseb_waitrequest	:	in	std_logic	:=	'0';
		cseb_wrresp_valid	:	in	std_logic	:=	'0';
		cseb_wrresponse	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		csr_cbdin	:	in	std_logic	:=	'0';
		csr_clk	:	in	std_logic	:=	'0';
		csr_din	:	in	std_logic	:=	'0';
		csr_en	:	in	std_logic	:=	'0';
		csr_enscan	:	in	std_logic	:=	'0';
		csr_entest	:	in	std_logic	:=	'0';
		csr_in	:	in	std_logic	:=	'0';
		csr_load_csr	:	in	std_logic	:=	'0';
		csr_pipe_in	:	in	std_logic	:=	'0';
		csr_seg	:	in	std_logic	:=	'0';
		csr_tcsrin	:	in	std_logic	:=	'0';
		csr_tverify	:	in	std_logic	:=	'0';
		cvp_config_done	:	in	std_logic	:=	'0';
		cvp_config_error	:	in	std_logic	:=	'0';
		cvp_config_ready	:	in	std_logic	:=	'0';
		cvp_en	:	in	std_logic	:=	'0';
		egress_blk_err	:	in	std_logic	:=	'0';
		entest	:	in	std_logic	:=	'0';
		flr_reset	:	in	std_logic	:=	'0';
		force_tx_eidle	:	in	std_logic	:=	'0';
		fref_clk0	:	in	std_logic	:=	'0';
		fref_clk1	:	in	std_logic	:=	'0';
		fref_clk2	:	in	std_logic	:=	'0';
		fref_clk3	:	in	std_logic	:=	'0';
		fref_clk4	:	in	std_logic	:=	'0';
		fref_clk5	:	in	std_logic	:=	'0';
		fref_clk6	:	in	std_logic	:=	'0';
		fref_clk7	:	in	std_logic	:=	'0';
		frzlogic	:	in	std_logic	:=	'0';
		frzreg	:	in	std_logic	:=	'0';
		hold_ltssm_rec	:	in	std_logic	:=	'0';
		hpg_ctrler	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		iocsrrdy_dly	:	in	std_logic	:=	'0';
		lmi_addr	:	in	std_logic_vector(11 downto 0)	:=	"000000000000";
		lmi_din	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		lmi_rden	:	in	std_logic	:=	'0';
		lmi_wren	:	in	std_logic	:=	'0';
		m10k_select	:	in	std_logic_vector(2 downto 0)	:=	"000";
		mask_tx_pll_lock0	:	in	std_logic	:=	'0';
		mask_tx_pll_lock1	:	in	std_logic	:=	'0';
		mask_tx_pll_lock2	:	in	std_logic	:=	'0';
		mask_tx_pll_lock3	:	in	std_logic	:=	'0';
		mask_tx_pll_lock4	:	in	std_logic	:=	'0';
		mask_tx_pll_lock5	:	in	std_logic	:=	'0';
		mask_tx_pll_lock6	:	in	std_logic	:=	'0';
		mask_tx_pll_lock7	:	in	std_logic	:=	'0';
		mem_hip_test_enable	:	in	std_logic	:=	'0';
		mem_regscanen_n	:	in	std_logic	:=	'0';
		mem_rscin_rcv_bot	:	in	std_logic	:=	'0';
		mem_rscin_rcv_top	:	in	std_logic	:=	'0';
		mem_rscin_rtry	:	in	std_logic	:=	'0';
		nfrzdrv	:	in	std_logic	:=	'0';
		npor	:	in	std_logic	:=	'0';
		pclk_central	:	in	std_logic	:=	'0';
		pclk_ch0	:	in	std_logic	:=	'0';
		pclk_ch1	:	in	std_logic	:=	'0';
		pex_msi_num	:	in	std_logic_vector(4 downto 0)	:=	"00000";
		phy_rst	:	in	std_logic	:=	'0';
		phy_srst	:	in	std_logic	:=	'0';
		phystatus0	:	in	std_logic	:=	'0';
		phystatus1	:	in	std_logic	:=	'0';
		phystatus2	:	in	std_logic	:=	'0';
		phystatus3	:	in	std_logic	:=	'0';
		phystatus4	:	in	std_logic	:=	'0';
		phystatus5	:	in	std_logic	:=	'0';
		phystatus6	:	in	std_logic	:=	'0';
		phystatus7	:	in	std_logic	:=	'0';
		pin_perst_n	:	in	std_logic	:=	'0';
		pld_clk	:	in	std_logic	:=	'0';
		pld_clrhip_n	:	in	std_logic	:=	'0';
		pld_clrpcship_n	:	in	std_logic	:=	'0';
		pld_clrpmapcship_n	:	in	std_logic	:=	'0';
		pld_core_ready	:	in	std_logic	:=	'0';
		pld_gp_status	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		pld_perst_n	:	in	std_logic	:=	'0';
		pll_cal_done0	:	in	std_logic	:=	'0';
		pll_cal_done1	:	in	std_logic	:=	'0';
		pll_cal_done2	:	in	std_logic	:=	'0';
		pll_cal_done3	:	in	std_logic	:=	'0';
		pll_cal_done4	:	in	std_logic	:=	'0';
		pll_cal_done5	:	in	std_logic	:=	'0';
		pll_cal_done6	:	in	std_logic	:=	'0';
		pll_cal_done7	:	in	std_logic	:=	'0';
		pll_fixed_clk_central	:	in	std_logic	:=	'0';
		pll_fixed_clk_ch0	:	in	std_logic	:=	'0';
		pll_fixed_clk_ch1	:	in	std_logic	:=	'0';
		plniotri	:	in	std_logic	:=	'0';
		pm_auxpwr	:	in	std_logic	:=	'0';
		pm_data	:	in	std_logic_vector(9 downto 0)	:=	"0000000000";
		pm_event	:	in	std_logic	:=	'0';
		pm_exit_d0_ack	:	in	std_logic	:=	'0';
		pme_to_cr	:	in	std_logic	:=	'0';
		reserved_clk_in	:	in	std_logic	:=	'0';
		reserved_in	:	in	std_logic_vector(7 downto 0)	:=	"00000000";
		rx_cred_ctl	:	in	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		rx_pll_freq_lock0	:	in	std_logic	:=	'0';
		rx_pll_freq_lock1	:	in	std_logic	:=	'0';
		rx_pll_freq_lock2	:	in	std_logic	:=	'0';
		rx_pll_freq_lock3	:	in	std_logic	:=	'0';
		rx_pll_freq_lock4	:	in	std_logic	:=	'0';
		rx_pll_freq_lock5	:	in	std_logic	:=	'0';
		rx_pll_freq_lock6	:	in	std_logic	:=	'0';
		rx_pll_freq_lock7	:	in	std_logic	:=	'0';
		rx_pll_phase_lock0	:	in	std_logic	:=	'0';
		rx_pll_phase_lock1	:	in	std_logic	:=	'0';
		rx_pll_phase_lock2	:	in	std_logic	:=	'0';
		rx_pll_phase_lock3	:	in	std_logic	:=	'0';
		rx_pll_phase_lock4	:	in	std_logic	:=	'0';
		rx_pll_phase_lock5	:	in	std_logic	:=	'0';
		rx_pll_phase_lock6	:	in	std_logic	:=	'0';
		rx_pll_phase_lock7	:	in	std_logic	:=	'0';
		rx_st_mask	:	in	std_logic	:=	'0';
		rx_st_ready	:	in	std_logic	:=	'0';
		rxblkst0	:	in	std_logic	:=	'0';
		rxblkst1	:	in	std_logic	:=	'0';
		rxblkst2	:	in	std_logic	:=	'0';
		rxblkst3	:	in	std_logic	:=	'0';
		rxblkst4	:	in	std_logic	:=	'0';
		rxblkst5	:	in	std_logic	:=	'0';
		rxblkst6	:	in	std_logic	:=	'0';
		rxblkst7	:	in	std_logic	:=	'0';
		rxdata0	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata1	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata2	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata3	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata4	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata5	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata6	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdata7	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rxdatak0	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak1	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak2	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak3	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak4	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak5	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak6	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdatak7	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		rxdataskip0	:	in	std_logic	:=	'0';
		rxdataskip1	:	in	std_logic	:=	'0';
		rxdataskip2	:	in	std_logic	:=	'0';
		rxdataskip3	:	in	std_logic	:=	'0';
		rxdataskip4	:	in	std_logic	:=	'0';
		rxdataskip5	:	in	std_logic	:=	'0';
		rxdataskip6	:	in	std_logic	:=	'0';
		rxdataskip7	:	in	std_logic	:=	'0';
		rxelecidle0	:	in	std_logic	:=	'0';
		rxelecidle1	:	in	std_logic	:=	'0';
		rxelecidle2	:	in	std_logic	:=	'0';
		rxelecidle3	:	in	std_logic	:=	'0';
		rxelecidle4	:	in	std_logic	:=	'0';
		rxelecidle5	:	in	std_logic	:=	'0';
		rxelecidle6	:	in	std_logic	:=	'0';
		rxelecidle7	:	in	std_logic	:=	'0';
		rxfreqlocked0	:	in	std_logic	:=	'0';
		rxfreqlocked1	:	in	std_logic	:=	'0';
		rxfreqlocked2	:	in	std_logic	:=	'0';
		rxfreqlocked3	:	in	std_logic	:=	'0';
		rxfreqlocked4	:	in	std_logic	:=	'0';
		rxfreqlocked5	:	in	std_logic	:=	'0';
		rxfreqlocked6	:	in	std_logic	:=	'0';
		rxfreqlocked7	:	in	std_logic	:=	'0';
		rxstatus0	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus1	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus2	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus3	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus4	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus5	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus6	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxstatus7	:	in	std_logic_vector(2 downto 0)	:=	"000";
		rxsynchd0	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd1	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd2	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd3	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd4	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd5	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd6	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxsynchd7	:	in	std_logic_vector(1 downto 0)	:=	"00";
		rxvalid0	:	in	std_logic	:=	'0';
		rxvalid1	:	in	std_logic	:=	'0';
		rxvalid2	:	in	std_logic	:=	'0';
		rxvalid3	:	in	std_logic	:=	'0';
		rxvalid4	:	in	std_logic	:=	'0';
		rxvalid5	:	in	std_logic	:=	'0';
		rxvalid6	:	in	std_logic	:=	'0';
		rxvalid7	:	in	std_logic	:=	'0';
		scan_mode_n	:	in	std_logic	:=	'0';
		scan_shift_n	:	in	std_logic	:=	'0';
		sw_ctmod	:	in	std_logic_vector(1 downto 0)	:=	"00";
		swdn_in	:	in	std_logic_vector(2 downto 0)	:=	"000";
		swup_in	:	in	std_logic_vector(6 downto 0)	:=	"0000000";
		test_in_1_hip	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		test_in_hip	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		test_pl_dbg_eqin	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		tx_cred_cons_select	:	in	std_logic	:=	'0';
		tx_cred_fc_sel	:	in	std_logic_vector(1 downto 0)	:=	"00";
		tx_lcff_pll_lock0	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock1	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock2	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock3	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock4	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock5	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock6	:	in	std_logic	:=	'0';
		tx_lcff_pll_lock7	:	in	std_logic	:=	'0';
		tx_st_data	:	in	std_logic_vector(255 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		tx_st_empty	:	in	std_logic_vector(1 downto 0)	:=	"00";
		tx_st_eop	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		tx_st_err	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		tx_st_parity	:	in	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		tx_st_sop	:	in	std_logic_vector(3 downto 0)	:=	"0000";
		tx_st_valid	:	in	std_logic	:=	'0';
		user_mode	:	in	std_logic	:=	'0';
		sta_hd_altpe3_hip_core_top_hd_altpe3_hip_core_u_clkmux_core_clk_cnt_reg_0_0_Q	:	out	std_logic	:=	'0';
		sta_hd_altpe3_hip_core_top_hd_altpe3_hip_core_u_clkmux_core_clk_cnt_reg_1_0_Q	:	out	std_logic	:=	'0';
		sta_hd_altpe3_hip_core_top_hd_altpe3_hip_core_u_clkmux_core_clk_cnt_reg_2_0_Q	:	out	std_logic	:=	'0';
		app_inta_ack	:	out	std_logic	:=	'0';
		app_msi_ack	:	out	std_logic	:=	'0';
		avmm_readdata	:	out	std_logic_vector(15 downto 0)	:=	"0000000000000000";
		cfg_par_err	:	out	std_logic	:=	'0';
		core_clk_out	:	out	std_logic	:=	'0';
		cseb_addr	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		cseb_addr_parity	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		cseb_be	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		cseb_is_shadow	:	out	std_logic	:=	'0';
		cseb_rden	:	out	std_logic	:=	'0';
		cseb_wrdata	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		cseb_wrdata_parity	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		cseb_wren	:	out	std_logic	:=	'0';
		cseb_wrresp_req	:	out	std_logic	:=	'0';
		csr_dout	:	out	std_logic	:=	'0';
		csr_out	:	out	std_logic	:=	'0';
		csr_pipe_out	:	out	std_logic	:=	'0';
		current_coeff0	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff1	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff2	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff3	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff4	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff5	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff6	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_coeff7	:	out	std_logic_vector(17 downto 0)	:=	"000000000000000000";
		current_rxpreset0	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset1	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset2	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset3	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset4	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset5	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset6	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_rxpreset7	:	out	std_logic_vector(2 downto 0)	:=	"000";
		current_speed	:	out	std_logic_vector(1 downto 0)	:=	"00";
		cvp_clk	:	out	std_logic	:=	'0';
		cvp_config	:	out	std_logic	:=	'0';
		cvp_data	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		cvp_full_config	:	out	std_logic	:=	'0';
		cvp_start_xfer	:	out	std_logic	:=	'0';
		dl_up	:	out	std_logic	:=	'0';
		dlup_exit	:	out	std_logic	:=	'0';
		eidle_infer_sel0	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel1	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel2	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel3	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel4	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel5	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel6	:	out	std_logic_vector(2 downto 0)	:=	"000";
		eidle_infer_sel7	:	out	std_logic_vector(2 downto 0)	:=	"000";
		ev_128ns	:	out	std_logic	:=	'0';
		ev_1us	:	out	std_logic	:=	'0';
		flr_sts	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n0	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n1	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n2	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n3	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n4	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n5	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n6	:	out	std_logic	:=	'0';
		g3_rx_pcs_rst_n7	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n0	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n1	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n2	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n3	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n4	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n5	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n6	:	out	std_logic	:=	'0';
		g3_tx_pcs_rst_n7	:	out	std_logic	:=	'0';
		hotrst_exit	:	out	std_logic	:=	'0';
		int_status	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		k_hip_pcs_chnl_en	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		k_hrc_chnl_en	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		k_hrc_chnl_txpll_master_cgb_rst_en	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		k_hrc_chnl_txpll_rst_en	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		l2_exit	:	out	std_logic	:=	'0';
		lane_act	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		lmi_ack	:	out	std_logic	:=	'0';
		lmi_dout	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		ltssm_state	:	out	std_logic_vector(4 downto 0)	:=	"00000";
		mem_rscout_rcv_bot	:	out	std_logic	:=	'0';
		mem_rscout_rcv_top	:	out	std_logic	:=	'0';
		mem_rscout_rtry	:	out	std_logic	:=	'0';
		pld_clk_in_use	:	out	std_logic	:=	'0';
		pld_gp_ctrl	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		pm_exit_d0_req	:	out	std_logic	:=	'0';
		pme_to_sr	:	out	std_logic	:=	'0';
		powerdown0	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown1	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown2	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown3	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown4	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown5	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown6	:	out	std_logic_vector(1 downto 0)	:=	"00";
		powerdown7	:	out	std_logic_vector(1 downto 0)	:=	"00";
		r2c_unc_ecc	:	out	std_logic	:=	'0';
		rate0	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate1	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate2	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate3	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate4	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate5	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate6	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate7	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rate_ctrl	:	out	std_logic_vector(1 downto 0)	:=	"00";
		reserved_clk_out	:	out	std_logic	:=	'0';
		reserved_out	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		reset_status	:	out	std_logic	:=	'0';
		retry_corr_ecc	:	out	std_logic	:=	'0';
		retry_unc_ecc	:	out	std_logic	:=	'0';
		rx_corr_ecc	:	out	std_logic	:=	'0';
		rx_cred_status	:	out	std_logic_vector(19 downto 0)	:=	"00000000000000000000";
		rx_par_err	:	out	std_logic	:=	'0';
		rx_pcs_rst_n0	:	out	std_logic	:=	'0';
		rx_pcs_rst_n1	:	out	std_logic	:=	'0';
		rx_pcs_rst_n2	:	out	std_logic	:=	'0';
		rx_pcs_rst_n3	:	out	std_logic	:=	'0';
		rx_pcs_rst_n4	:	out	std_logic	:=	'0';
		rx_pcs_rst_n5	:	out	std_logic	:=	'0';
		rx_pcs_rst_n6	:	out	std_logic	:=	'0';
		rx_pcs_rst_n7	:	out	std_logic	:=	'0';
		rx_pma_rstb0	:	out	std_logic	:=	'0';
		rx_pma_rstb1	:	out	std_logic	:=	'0';
		rx_pma_rstb2	:	out	std_logic	:=	'0';
		rx_pma_rstb3	:	out	std_logic	:=	'0';
		rx_pma_rstb4	:	out	std_logic	:=	'0';
		rx_pma_rstb5	:	out	std_logic	:=	'0';
		rx_pma_rstb6	:	out	std_logic	:=	'0';
		rx_pma_rstb7	:	out	std_logic	:=	'0';
		rx_st_bardec1	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		rx_st_bardec2	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		rx_st_be	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rx_st_data	:	out	std_logic_vector(255 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		rx_st_empty	:	out	std_logic_vector(1 downto 0)	:=	"00";
		rx_st_eop	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		rx_st_err	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		rx_st_parity	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		rx_st_sop	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		rx_st_valid	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		rxfc_cplbuf_ovf	:	out	std_logic	:=	'0';
		rxfc_cplovf_tag	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		rxpolarity0	:	out	std_logic	:=	'0';
		rxpolarity1	:	out	std_logic	:=	'0';
		rxpolarity2	:	out	std_logic	:=	'0';
		rxpolarity3	:	out	std_logic	:=	'0';
		rxpolarity4	:	out	std_logic	:=	'0';
		rxpolarity5	:	out	std_logic	:=	'0';
		rxpolarity6	:	out	std_logic	:=	'0';
		rxpolarity7	:	out	std_logic	:=	'0';
		serr_out	:	out	std_logic	:=	'0';
		swdn_out	:	out	std_logic_vector(6 downto 0)	:=	"0000000";
		swup_out	:	out	std_logic_vector(2 downto 0)	:=	"000";
		test_fref_clk	:	out	std_logic	:=	'0';
		test_out_1_hip	:	out	std_logic_vector(63 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000";
		test_out_hip	:	out	std_logic_vector(255 downto 0)	:=	"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		tl_cfg_add	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		tl_cfg_ctl	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		tl_cfg_sts	:	out	std_logic_vector(52 downto 0)	:=	"00000000000000000000000000000000000000000000000000000";
		tl_cfg_sts_wr	:	out	std_logic	:=	'0';
		tx_cred_data_fc	:	out	std_logic_vector(11 downto 0)	:=	"000000000000";
		tx_cred_fc_hip_cons	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		tx_cred_fc_infinite	:	out	std_logic_vector(5 downto 0)	:=	"000000";
		tx_cred_hdr_fc	:	out	std_logic_vector(7 downto 0)	:=	"00000000";
		tx_deemph0	:	out	std_logic	:=	'0';
		tx_deemph1	:	out	std_logic	:=	'0';
		tx_deemph2	:	out	std_logic	:=	'0';
		tx_deemph3	:	out	std_logic	:=	'0';
		tx_deemph4	:	out	std_logic	:=	'0';
		tx_deemph5	:	out	std_logic	:=	'0';
		tx_deemph6	:	out	std_logic	:=	'0';
		tx_deemph7	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb0	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb1	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb2	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb3	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb4	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb5	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb6	:	out	std_logic	:=	'0';
		tx_lcff_pll_rstb7	:	out	std_logic	:=	'0';
		tx_margin0	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin1	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin2	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin3	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin4	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin5	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin6	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_margin7	:	out	std_logic_vector(2 downto 0)	:=	"000";
		tx_par_err	:	out	std_logic_vector(1 downto 0)	:=	"00";
		tx_pcs_rst_n0	:	out	std_logic	:=	'0';
		tx_pcs_rst_n1	:	out	std_logic	:=	'0';
		tx_pcs_rst_n2	:	out	std_logic	:=	'0';
		tx_pcs_rst_n3	:	out	std_logic	:=	'0';
		tx_pcs_rst_n4	:	out	std_logic	:=	'0';
		tx_pcs_rst_n5	:	out	std_logic	:=	'0';
		tx_pcs_rst_n6	:	out	std_logic	:=	'0';
		tx_pcs_rst_n7	:	out	std_logic	:=	'0';
		tx_pma_syncp0	:	out	std_logic	:=	'0';
		tx_pma_syncp1	:	out	std_logic	:=	'0';
		tx_pma_syncp2	:	out	std_logic	:=	'0';
		tx_pma_syncp3	:	out	std_logic	:=	'0';
		tx_pma_syncp4	:	out	std_logic	:=	'0';
		tx_pma_syncp5	:	out	std_logic	:=	'0';
		tx_pma_syncp6	:	out	std_logic	:=	'0';
		tx_pma_syncp7	:	out	std_logic	:=	'0';
		tx_st_ready	:	out	std_logic	:=	'0';
		txblkst0	:	out	std_logic	:=	'0';
		txblkst1	:	out	std_logic	:=	'0';
		txblkst2	:	out	std_logic	:=	'0';
		txblkst3	:	out	std_logic	:=	'0';
		txblkst4	:	out	std_logic	:=	'0';
		txblkst5	:	out	std_logic	:=	'0';
		txblkst6	:	out	std_logic	:=	'0';
		txblkst7	:	out	std_logic	:=	'0';
		txcompl0	:	out	std_logic	:=	'0';
		txcompl1	:	out	std_logic	:=	'0';
		txcompl2	:	out	std_logic	:=	'0';
		txcompl3	:	out	std_logic	:=	'0';
		txcompl4	:	out	std_logic	:=	'0';
		txcompl5	:	out	std_logic	:=	'0';
		txcompl6	:	out	std_logic	:=	'0';
		txcompl7	:	out	std_logic	:=	'0';
		txdata0	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata1	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata2	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata3	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata4	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata5	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata6	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdata7	:	out	std_logic_vector(31 downto 0)	:=	"00000000000000000000000000000000";
		txdatak0	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak1	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak2	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak3	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak4	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak5	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak6	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdatak7	:	out	std_logic_vector(3 downto 0)	:=	"0000";
		txdataskip0	:	out	std_logic	:=	'0';
		txdataskip1	:	out	std_logic	:=	'0';
		txdataskip2	:	out	std_logic	:=	'0';
		txdataskip3	:	out	std_logic	:=	'0';
		txdataskip4	:	out	std_logic	:=	'0';
		txdataskip5	:	out	std_logic	:=	'0';
		txdataskip6	:	out	std_logic	:=	'0';
		txdataskip7	:	out	std_logic	:=	'0';
		txdetectrx0	:	out	std_logic	:=	'0';
		txdetectrx1	:	out	std_logic	:=	'0';
		txdetectrx2	:	out	std_logic	:=	'0';
		txdetectrx3	:	out	std_logic	:=	'0';
		txdetectrx4	:	out	std_logic	:=	'0';
		txdetectrx5	:	out	std_logic	:=	'0';
		txdetectrx6	:	out	std_logic	:=	'0';
		txdetectrx7	:	out	std_logic	:=	'0';
		txelecidle0	:	out	std_logic	:=	'0';
		txelecidle1	:	out	std_logic	:=	'0';
		txelecidle2	:	out	std_logic	:=	'0';
		txelecidle3	:	out	std_logic	:=	'0';
		txelecidle4	:	out	std_logic	:=	'0';
		txelecidle5	:	out	std_logic	:=	'0';
		txelecidle6	:	out	std_logic	:=	'0';
		txelecidle7	:	out	std_logic	:=	'0';
		txst_prot_err	:	out	std_logic	:=	'0';
		txswing0	:	out	std_logic	:=	'0';
		txswing1	:	out	std_logic	:=	'0';
		txswing2	:	out	std_logic	:=	'0';
		txswing3	:	out	std_logic	:=	'0';
		txswing4	:	out	std_logic	:=	'0';
		txswing5	:	out	std_logic	:=	'0';
		txswing6	:	out	std_logic	:=	'0';
		txswing7	:	out	std_logic	:=	'0';
		txsynchd0	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd1	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd2	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd3	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd4	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd5	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd6	:	out	std_logic_vector(1 downto 0)	:=	"00";
		txsynchd7	:	out	std_logic_vector(1 downto 0)	:=	"00";
		wake_oen	:	out	std_logic	:=	'0'
	);
end component;

begin



inst : twentynm_hssi_gen3_x8_pcie_hip_encrypted
	generic map (
		-- Instance parameters
		acknack_base	=>	acknack_base_int,
		acknack_set	=>	acknack_set,
		advance_error_reporting	=>	advance_error_reporting,
		app_interface_width	=>	app_interface_width,
		arb_upfc_30us_counter	=>	arb_upfc_30us_counter_int,
		arb_upfc_30us_en	=>	arb_upfc_30us_en,
		aspm_config_management	=>	aspm_config_management,
		aspm_patch_disable	=>	aspm_patch_disable,
		ast_width_rx	=>	ast_width_rx,
		ast_width_tx	=>	ast_width_tx,
		atomic_malformed	=>	atomic_malformed,
		atomic_op_completer_32bit	=>	atomic_op_completer_32bit,
		atomic_op_completer_64bit	=>	atomic_op_completer_64bit,
		atomic_op_routing	=>	atomic_op_routing,
		auto_msg_drop_enable	=>	auto_msg_drop_enable,
		avmm_cvp_inter_sel_csr_ctrl	=>	avmm_cvp_inter_sel_csr_ctrl,
		avmm_dprio_broadcast_en_csr_ctrl	=>	avmm_dprio_broadcast_en_csr_ctrl,
		avmm_force_inter_sel_csr_ctrl	=>	avmm_force_inter_sel_csr_ctrl,
		avmm_power_iso_en_csr_ctrl	=>	avmm_power_iso_en_csr_ctrl,
		bar0_size_mask	=>	bar0_size_mask_int,
		bar0_type	=>	bar0_type,
		bar1_size_mask	=>	bar1_size_mask_int,
		bar1_type	=>	bar1_type,
		bar2_size_mask	=>	bar2_size_mask_int,
		bar2_type	=>	bar2_type,
		bar3_size_mask	=>	bar3_size_mask_int,
		bar3_type	=>	bar3_type,
		bar4_size_mask	=>	bar4_size_mask_int,
		bar4_type	=>	bar4_type,
		bar5_size_mask	=>	bar5_size_mask_int,
		bar5_type	=>	bar5_type,
		base_counter_sel	=>	base_counter_sel,
		bist_memory_settings	=>	bist_memory_settings,
		bridge_port_ssid_support	=>	bridge_port_ssid_support,
		bridge_port_vga_enable	=>	bridge_port_vga_enable,
		bypass_cdc	=>	bypass_cdc,
		bypass_clk_switch	=>	bypass_clk_switch,
		bypass_tl	=>	bypass_tl,
		capab_rate_rxcfg_en	=>	capab_rate_rxcfg_en,
		cas_completer_128bit	=>	cas_completer_128bit,
		cdc_clk_relation	=>	cdc_clk_relation,
		cdc_dummy_insert_limit	=>	cdc_dummy_insert_limit_int,
		cfg_parchk_ena	=>	cfg_parchk_ena,
		cfgbp_req_recov_disable	=>	cfgbp_req_recov_disable,
		class_code	=>	class_code_int,
		clock_pwr_management	=>	clock_pwr_management,
		completion_timeout	=>	completion_timeout,
		core_clk_divider	=>	core_clk_divider,
		core_clk_freq_mhz	=>	core_clk_freq_mhz,
		core_clk_out_sel	=>	core_clk_out_sel,
		core_clk_sel	=>	core_clk_sel,
		core_clk_source	=>	core_clk_source,
		cseb_bar_match_checking	=>	cseb_bar_match_checking,
		cseb_config_bypass	=>	cseb_config_bypass,
		cseb_cpl_status_during_cvp	=>	cseb_cpl_status_during_cvp,
		cseb_cpl_tag_checking	=>	cseb_cpl_tag_checking,
		cseb_disable_auto_crs	=>	cseb_disable_auto_crs,
		cseb_extend_pci	=>	cseb_extend_pci,
		cseb_extend_pcie	=>	cseb_extend_pcie,
		cseb_min_error_checking	=>	cseb_min_error_checking,
		cseb_route_to_avl_rx_st	=>	cseb_route_to_avl_rx_st,
		cseb_temp_busy_crs	=>	cseb_temp_busy_crs,
		cvp_clk_reset	=>	cvp_clk_reset,
		cvp_data_compressed	=>	cvp_data_compressed,
		cvp_data_encrypted	=>	cvp_data_encrypted,
		cvp_enable	=>	cvp_enable,
		cvp_mode_reset	=>	cvp_mode_reset,
		cvp_rate_sel	=>	cvp_rate_sel,
		d0_pme	=>	d0_pme,
		d1_pme	=>	d1_pme,
		d1_support	=>	d1_support,
		d2_pme	=>	d2_pme,
		d2_support	=>	d2_support,
		d3_cold_pme	=>	d3_cold_pme,
		d3_hot_pme	=>	d3_hot_pme,
		data_pack_rx	=>	data_pack_rx,
		deemphasis_enable	=>	deemphasis_enable,
		deskew_comma	=>	deskew_comma,
		device_id	=>	device_id_int,
		device_number	=>	device_number_int,
		device_specific_init	=>	device_specific_init,
		dft_clock_obsrv_en	=>	dft_clock_obsrv_en,
		dft_clock_obsrv_sel	=>	dft_clock_obsrv_sel,
		diffclock_nfts_count	=>	diffclock_nfts_count_int,
		dis_cplovf	=>	dis_cplovf,
		dis_paritychk	=>	dis_paritychk,
		disable_link_x2_support	=>	disable_link_x2_support,
		disable_snoop_packet	=>	disable_snoop_packet,
		dl_tx_check_parity_edb	=>	dl_tx_check_parity_edb,
		dll_active_report_support	=>	dll_active_report_support,
		early_dl_up	=>	early_dl_up,
		eco_fb332688_dis	=>	eco_fb332688_dis,
		ecrc_check_capable	=>	ecrc_check_capable,
		ecrc_gen_capable	=>	ecrc_gen_capable,
		egress_block_err_report_ena	=>	egress_block_err_report_ena,
		ei_delay_powerdown_count	=>	ei_delay_powerdown_count_int,
		eie_before_nfts_count	=>	eie_before_nfts_count_int,
		electromech_interlock	=>	electromech_interlock,
		en_ieiupdatefc	=>	en_ieiupdatefc,
		en_lane_errchk	=>	en_lane_errchk,
		en_phystatus_dly	=>	en_phystatus_dly,
		ena_ido_cpl	=>	ena_ido_cpl,
		ena_ido_req	=>	ena_ido_req,
		enable_adapter_half_rate_mode	=>	enable_adapter_half_rate_mode,
		enable_ch01_pclk_out	=>	enable_ch01_pclk_out,
		enable_ch0_pclk_out	=>	enable_ch0_pclk_out,
		enable_completion_timeout_disable	=>	enable_completion_timeout_disable,
		enable_directed_spd_chng	=>	enable_directed_spd_chng,
		enable_function_msix_support	=>	enable_function_msix_support,
		enable_l0s_aspm	=>	enable_l0s_aspm,
		enable_l1_aspm	=>	enable_l1_aspm,
		enable_rx_buffer_checking	=>	enable_rx_buffer_checking,
		enable_rx_reordering	=>	enable_rx_reordering,
		enable_slot_register	=>	enable_slot_register,
		endpoint_l0_latency	=>	endpoint_l0_latency_int,
		endpoint_l1_latency	=>	endpoint_l1_latency_int,
		eql_rq_int_en_number	=>	eql_rq_int_en_number_int,
		errmgt_fcpe_patch_dis	=>	errmgt_fcpe_patch_dis,
		errmgt_fep_patch_dis	=>	errmgt_fep_patch_dis,
		expansion_base_address_register	=>	expansion_base_address_register,
		extend_tag_field	=>	extend_tag_field,
		extended_format_field	=>	extended_format_field,
		extended_tag_reset	=>	extended_tag_reset,
		fc_init_timer	=>	fc_init_timer_int,
		flow_control_timeout_count	=>	flow_control_timeout_count_int,
		flow_control_update_count	=>	flow_control_update_count_int,
		flr_capability	=>	flr_capability,
		force_dis_to_det	=>	force_dis_to_det,
		force_gen1_dis	=>	force_gen1_dis,
		force_tx_coeff_preset_lpbk	=>	force_tx_coeff_preset_lpbk,
		frame_err_patch_dis	=>	frame_err_patch_dis,
		func_mode	=>	func_mode,
		g3_bypass_equlz	=>	g3_bypass_equlz,
		g3_coeff_done_tmout	=>	g3_coeff_done_tmout,
		g3_deskew_char	=>	g3_deskew_char,
		g3_dis_be_frm_err	=>	g3_dis_be_frm_err,
		g3_dn_rx_hint_eqlz_0	=>	g3_dn_rx_hint_eqlz_0_int,
		g3_dn_rx_hint_eqlz_1	=>	g3_dn_rx_hint_eqlz_1_int,
		g3_dn_rx_hint_eqlz_2	=>	g3_dn_rx_hint_eqlz_2_int,
		g3_dn_rx_hint_eqlz_3	=>	g3_dn_rx_hint_eqlz_3_int,
		g3_dn_rx_hint_eqlz_4	=>	g3_dn_rx_hint_eqlz_4_int,
		g3_dn_rx_hint_eqlz_5	=>	g3_dn_rx_hint_eqlz_5_int,
		g3_dn_rx_hint_eqlz_6	=>	g3_dn_rx_hint_eqlz_6_int,
		g3_dn_rx_hint_eqlz_7	=>	g3_dn_rx_hint_eqlz_7_int,
		g3_dn_tx_preset_eqlz_0	=>	g3_dn_tx_preset_eqlz_0_int,
		g3_dn_tx_preset_eqlz_1	=>	g3_dn_tx_preset_eqlz_1_int,
		g3_dn_tx_preset_eqlz_2	=>	g3_dn_tx_preset_eqlz_2_int,
		g3_dn_tx_preset_eqlz_3	=>	g3_dn_tx_preset_eqlz_3_int,
		g3_dn_tx_preset_eqlz_4	=>	g3_dn_tx_preset_eqlz_4_int,
		g3_dn_tx_preset_eqlz_5	=>	g3_dn_tx_preset_eqlz_5_int,
		g3_dn_tx_preset_eqlz_6	=>	g3_dn_tx_preset_eqlz_6_int,
		g3_dn_tx_preset_eqlz_7	=>	g3_dn_tx_preset_eqlz_7_int,
		g3_force_ber_max	=>	g3_force_ber_max,
		g3_force_ber_min	=>	g3_force_ber_min,
		g3_lnk_trn_rx_ts	=>	g3_lnk_trn_rx_ts,
		g3_ltssm_eq_dbg	=>	g3_ltssm_eq_dbg,
		g3_ltssm_rec_dbg	=>	g3_ltssm_rec_dbg,
		g3_pause_ltssm_rec_en	=>	g3_pause_ltssm_rec_en,
		g3_quiesce_guarant	=>	g3_quiesce_guarant,
		g3_redo_equlz_dis	=>	g3_redo_equlz_dis,
		g3_redo_equlz_en	=>	g3_redo_equlz_en,
		g3_up_rx_hint_eqlz_0	=>	g3_up_rx_hint_eqlz_0_int,
		g3_up_rx_hint_eqlz_1	=>	g3_up_rx_hint_eqlz_1_int,
		g3_up_rx_hint_eqlz_2	=>	g3_up_rx_hint_eqlz_2_int,
		g3_up_rx_hint_eqlz_3	=>	g3_up_rx_hint_eqlz_3_int,
		g3_up_rx_hint_eqlz_4	=>	g3_up_rx_hint_eqlz_4_int,
		g3_up_rx_hint_eqlz_5	=>	g3_up_rx_hint_eqlz_5_int,
		g3_up_rx_hint_eqlz_6	=>	g3_up_rx_hint_eqlz_6_int,
		g3_up_rx_hint_eqlz_7	=>	g3_up_rx_hint_eqlz_7_int,
		g3_up_tx_preset_eqlz_0	=>	g3_up_tx_preset_eqlz_0_int,
		g3_up_tx_preset_eqlz_1	=>	g3_up_tx_preset_eqlz_1_int,
		g3_up_tx_preset_eqlz_2	=>	g3_up_tx_preset_eqlz_2_int,
		g3_up_tx_preset_eqlz_3	=>	g3_up_tx_preset_eqlz_3_int,
		g3_up_tx_preset_eqlz_4	=>	g3_up_tx_preset_eqlz_4_int,
		g3_up_tx_preset_eqlz_5	=>	g3_up_tx_preset_eqlz_5_int,
		g3_up_tx_preset_eqlz_6	=>	g3_up_tx_preset_eqlz_6_int,
		g3_up_tx_preset_eqlz_7	=>	g3_up_tx_preset_eqlz_7_int,
		gen123_lane_rate_mode	=>	gen123_lane_rate_mode,
		gen2_diffclock_nfts_count	=>	gen2_diffclock_nfts_count_int,
		gen2_pma_pll_usage	=>	gen2_pma_pll_usage,
		gen2_sameclock_nfts_count	=>	gen2_sameclock_nfts_count_int,
		gen3_coeff_1	=>	gen3_coeff_1_int,
		gen3_coeff_10	=>	gen3_coeff_10_int,
		gen3_coeff_10_ber_meas	=>	gen3_coeff_10_ber_meas_int,
		gen3_coeff_10_nxtber_less	=>	gen3_coeff_10_nxtber_less_int,
		gen3_coeff_10_nxtber_more	=>	gen3_coeff_10_nxtber_more_int,
		gen3_coeff_10_preset_hint	=>	gen3_coeff_10_preset_hint_int,
		gen3_coeff_10_reqber	=>	gen3_coeff_10_reqber_int,
		gen3_coeff_10_sel	=>	gen3_coeff_10_sel,
		gen3_coeff_11	=>	gen3_coeff_11_int,
		gen3_coeff_11_ber_meas	=>	gen3_coeff_11_ber_meas_int,
		gen3_coeff_11_nxtber_less	=>	gen3_coeff_11_nxtber_less_int,
		gen3_coeff_11_nxtber_more	=>	gen3_coeff_11_nxtber_more_int,
		gen3_coeff_11_preset_hint	=>	gen3_coeff_11_preset_hint_int,
		gen3_coeff_11_reqber	=>	gen3_coeff_11_reqber_int,
		gen3_coeff_11_sel	=>	gen3_coeff_11_sel,
		gen3_coeff_12	=>	gen3_coeff_12_int,
		gen3_coeff_12_ber_meas	=>	gen3_coeff_12_ber_meas_int,
		gen3_coeff_12_nxtber_less	=>	gen3_coeff_12_nxtber_less_int,
		gen3_coeff_12_nxtber_more	=>	gen3_coeff_12_nxtber_more_int,
		gen3_coeff_12_preset_hint	=>	gen3_coeff_12_preset_hint_int,
		gen3_coeff_12_reqber	=>	gen3_coeff_12_reqber_int,
		gen3_coeff_12_sel	=>	gen3_coeff_12_sel,
		gen3_coeff_13	=>	gen3_coeff_13_int,
		gen3_coeff_13_ber_meas	=>	gen3_coeff_13_ber_meas_int,
		gen3_coeff_13_nxtber_less	=>	gen3_coeff_13_nxtber_less_int,
		gen3_coeff_13_nxtber_more	=>	gen3_coeff_13_nxtber_more_int,
		gen3_coeff_13_preset_hint	=>	gen3_coeff_13_preset_hint_int,
		gen3_coeff_13_reqber	=>	gen3_coeff_13_reqber_int,
		gen3_coeff_13_sel	=>	gen3_coeff_13_sel,
		gen3_coeff_14	=>	gen3_coeff_14_int,
		gen3_coeff_14_ber_meas	=>	gen3_coeff_14_ber_meas_int,
		gen3_coeff_14_nxtber_less	=>	gen3_coeff_14_nxtber_less_int,
		gen3_coeff_14_nxtber_more	=>	gen3_coeff_14_nxtber_more_int,
		gen3_coeff_14_preset_hint	=>	gen3_coeff_14_preset_hint_int,
		gen3_coeff_14_reqber	=>	gen3_coeff_14_reqber_int,
		gen3_coeff_14_sel	=>	gen3_coeff_14_sel,
		gen3_coeff_15	=>	gen3_coeff_15_int,
		gen3_coeff_15_ber_meas	=>	gen3_coeff_15_ber_meas_int,
		gen3_coeff_15_nxtber_less	=>	gen3_coeff_15_nxtber_less_int,
		gen3_coeff_15_nxtber_more	=>	gen3_coeff_15_nxtber_more_int,
		gen3_coeff_15_preset_hint	=>	gen3_coeff_15_preset_hint_int,
		gen3_coeff_15_reqber	=>	gen3_coeff_15_reqber_int,
		gen3_coeff_15_sel	=>	gen3_coeff_15_sel,
		gen3_coeff_16	=>	gen3_coeff_16_int,
		gen3_coeff_16_ber_meas	=>	gen3_coeff_16_ber_meas_int,
		gen3_coeff_16_nxtber_less	=>	gen3_coeff_16_nxtber_less_int,
		gen3_coeff_16_nxtber_more	=>	gen3_coeff_16_nxtber_more_int,
		gen3_coeff_16_preset_hint	=>	gen3_coeff_16_preset_hint_int,
		gen3_coeff_16_reqber	=>	gen3_coeff_16_reqber_int,
		gen3_coeff_16_sel	=>	gen3_coeff_16_sel,
		gen3_coeff_17	=>	gen3_coeff_17_int,
		gen3_coeff_17_ber_meas	=>	gen3_coeff_17_ber_meas_int,
		gen3_coeff_17_nxtber_less	=>	gen3_coeff_17_nxtber_less_int,
		gen3_coeff_17_nxtber_more	=>	gen3_coeff_17_nxtber_more_int,
		gen3_coeff_17_preset_hint	=>	gen3_coeff_17_preset_hint_int,
		gen3_coeff_17_reqber	=>	gen3_coeff_17_reqber_int,
		gen3_coeff_17_sel	=>	gen3_coeff_17_sel,
		gen3_coeff_18	=>	gen3_coeff_18_int,
		gen3_coeff_18_ber_meas	=>	gen3_coeff_18_ber_meas_int,
		gen3_coeff_18_nxtber_less	=>	gen3_coeff_18_nxtber_less_int,
		gen3_coeff_18_nxtber_more	=>	gen3_coeff_18_nxtber_more_int,
		gen3_coeff_18_preset_hint	=>	gen3_coeff_18_preset_hint_int,
		gen3_coeff_18_reqber	=>	gen3_coeff_18_reqber_int,
		gen3_coeff_18_sel	=>	gen3_coeff_18_sel,
		gen3_coeff_19	=>	gen3_coeff_19_int,
		gen3_coeff_19_ber_meas	=>	gen3_coeff_19_ber_meas_int,
		gen3_coeff_19_nxtber_less	=>	gen3_coeff_19_nxtber_less_int,
		gen3_coeff_19_nxtber_more	=>	gen3_coeff_19_nxtber_more_int,
		gen3_coeff_19_preset_hint	=>	gen3_coeff_19_preset_hint_int,
		gen3_coeff_19_reqber	=>	gen3_coeff_19_reqber_int,
		gen3_coeff_19_sel	=>	gen3_coeff_19_sel,
		gen3_coeff_1_ber_meas	=>	gen3_coeff_1_ber_meas_int,
		gen3_coeff_1_nxtber_less	=>	gen3_coeff_1_nxtber_less_int,
		gen3_coeff_1_nxtber_more	=>	gen3_coeff_1_nxtber_more_int,
		gen3_coeff_1_preset_hint	=>	gen3_coeff_1_preset_hint_int,
		gen3_coeff_1_reqber	=>	gen3_coeff_1_reqber_int,
		gen3_coeff_1_sel	=>	gen3_coeff_1_sel,
		gen3_coeff_2	=>	gen3_coeff_2_int,
		gen3_coeff_20	=>	gen3_coeff_20_int,
		gen3_coeff_20_ber_meas	=>	gen3_coeff_20_ber_meas_int,
		gen3_coeff_20_nxtber_less	=>	gen3_coeff_20_nxtber_less_int,
		gen3_coeff_20_nxtber_more	=>	gen3_coeff_20_nxtber_more_int,
		gen3_coeff_20_preset_hint	=>	gen3_coeff_20_preset_hint_int,
		gen3_coeff_20_reqber	=>	gen3_coeff_20_reqber_int,
		gen3_coeff_20_sel	=>	gen3_coeff_20_sel,
		gen3_coeff_21	=>	gen3_coeff_21_int,
		gen3_coeff_21_ber_meas	=>	gen3_coeff_21_ber_meas_int,
		gen3_coeff_21_nxtber_less	=>	gen3_coeff_21_nxtber_less_int,
		gen3_coeff_21_nxtber_more	=>	gen3_coeff_21_nxtber_more_int,
		gen3_coeff_21_preset_hint	=>	gen3_coeff_21_preset_hint_int,
		gen3_coeff_21_reqber	=>	gen3_coeff_21_reqber_int,
		gen3_coeff_21_sel	=>	gen3_coeff_21_sel,
		gen3_coeff_22	=>	gen3_coeff_22_int,
		gen3_coeff_22_ber_meas	=>	gen3_coeff_22_ber_meas_int,
		gen3_coeff_22_nxtber_less	=>	gen3_coeff_22_nxtber_less_int,
		gen3_coeff_22_nxtber_more	=>	gen3_coeff_22_nxtber_more_int,
		gen3_coeff_22_preset_hint	=>	gen3_coeff_22_preset_hint_int,
		gen3_coeff_22_reqber	=>	gen3_coeff_22_reqber_int,
		gen3_coeff_22_sel	=>	gen3_coeff_22_sel,
		gen3_coeff_23	=>	gen3_coeff_23_int,
		gen3_coeff_23_ber_meas	=>	gen3_coeff_23_ber_meas_int,
		gen3_coeff_23_nxtber_less	=>	gen3_coeff_23_nxtber_less_int,
		gen3_coeff_23_nxtber_more	=>	gen3_coeff_23_nxtber_more_int,
		gen3_coeff_23_preset_hint	=>	gen3_coeff_23_preset_hint_int,
		gen3_coeff_23_reqber	=>	gen3_coeff_23_reqber_int,
		gen3_coeff_23_sel	=>	gen3_coeff_23_sel,
		gen3_coeff_24	=>	gen3_coeff_24_int,
		gen3_coeff_24_ber_meas	=>	gen3_coeff_24_ber_meas_int,
		gen3_coeff_24_nxtber_less	=>	gen3_coeff_24_nxtber_less_int,
		gen3_coeff_24_nxtber_more	=>	gen3_coeff_24_nxtber_more_int,
		gen3_coeff_24_preset_hint	=>	gen3_coeff_24_preset_hint_int,
		gen3_coeff_24_reqber	=>	gen3_coeff_24_reqber_int,
		gen3_coeff_24_sel	=>	gen3_coeff_24_sel,
		gen3_coeff_2_ber_meas	=>	gen3_coeff_2_ber_meas_int,
		gen3_coeff_2_nxtber_less	=>	gen3_coeff_2_nxtber_less_int,
		gen3_coeff_2_nxtber_more	=>	gen3_coeff_2_nxtber_more_int,
		gen3_coeff_2_preset_hint	=>	gen3_coeff_2_preset_hint_int,
		gen3_coeff_2_reqber	=>	gen3_coeff_2_reqber_int,
		gen3_coeff_2_sel	=>	gen3_coeff_2_sel,
		gen3_coeff_3	=>	gen3_coeff_3_int,
		gen3_coeff_3_ber_meas	=>	gen3_coeff_3_ber_meas_int,
		gen3_coeff_3_nxtber_less	=>	gen3_coeff_3_nxtber_less_int,
		gen3_coeff_3_nxtber_more	=>	gen3_coeff_3_nxtber_more_int,
		gen3_coeff_3_preset_hint	=>	gen3_coeff_3_preset_hint_int,
		gen3_coeff_3_reqber	=>	gen3_coeff_3_reqber_int,
		gen3_coeff_3_sel	=>	gen3_coeff_3_sel,
		gen3_coeff_4	=>	gen3_coeff_4_int,
		gen3_coeff_4_ber_meas	=>	gen3_coeff_4_ber_meas_int,
		gen3_coeff_4_nxtber_less	=>	gen3_coeff_4_nxtber_less_int,
		gen3_coeff_4_nxtber_more	=>	gen3_coeff_4_nxtber_more_int,
		gen3_coeff_4_preset_hint	=>	gen3_coeff_4_preset_hint_int,
		gen3_coeff_4_reqber	=>	gen3_coeff_4_reqber_int,
		gen3_coeff_4_sel	=>	gen3_coeff_4_sel,
		gen3_coeff_5	=>	gen3_coeff_5_int,
		gen3_coeff_5_ber_meas	=>	gen3_coeff_5_ber_meas_int,
		gen3_coeff_5_nxtber_less	=>	gen3_coeff_5_nxtber_less_int,
		gen3_coeff_5_nxtber_more	=>	gen3_coeff_5_nxtber_more_int,
		gen3_coeff_5_preset_hint	=>	gen3_coeff_5_preset_hint_int,
		gen3_coeff_5_reqber	=>	gen3_coeff_5_reqber_int,
		gen3_coeff_5_sel	=>	gen3_coeff_5_sel,
		gen3_coeff_6	=>	gen3_coeff_6_int,
		gen3_coeff_6_ber_meas	=>	gen3_coeff_6_ber_meas_int,
		gen3_coeff_6_nxtber_less	=>	gen3_coeff_6_nxtber_less_int,
		gen3_coeff_6_nxtber_more	=>	gen3_coeff_6_nxtber_more_int,
		gen3_coeff_6_preset_hint	=>	gen3_coeff_6_preset_hint_int,
		gen3_coeff_6_reqber	=>	gen3_coeff_6_reqber_int,
		gen3_coeff_6_sel	=>	gen3_coeff_6_sel,
		gen3_coeff_7	=>	gen3_coeff_7_int,
		gen3_coeff_7_ber_meas	=>	gen3_coeff_7_ber_meas_int,
		gen3_coeff_7_nxtber_less	=>	gen3_coeff_7_nxtber_less_int,
		gen3_coeff_7_nxtber_more	=>	gen3_coeff_7_nxtber_more_int,
		gen3_coeff_7_preset_hint	=>	gen3_coeff_7_preset_hint_int,
		gen3_coeff_7_reqber	=>	gen3_coeff_7_reqber_int,
		gen3_coeff_7_sel	=>	gen3_coeff_7_sel,
		gen3_coeff_8	=>	gen3_coeff_8_int,
		gen3_coeff_8_ber_meas	=>	gen3_coeff_8_ber_meas_int,
		gen3_coeff_8_nxtber_less	=>	gen3_coeff_8_nxtber_less_int,
		gen3_coeff_8_nxtber_more	=>	gen3_coeff_8_nxtber_more_int,
		gen3_coeff_8_preset_hint	=>	gen3_coeff_8_preset_hint_int,
		gen3_coeff_8_reqber	=>	gen3_coeff_8_reqber_int,
		gen3_coeff_8_sel	=>	gen3_coeff_8_sel,
		gen3_coeff_9	=>	gen3_coeff_9_int,
		gen3_coeff_9_ber_meas	=>	gen3_coeff_9_ber_meas_int,
		gen3_coeff_9_nxtber_less	=>	gen3_coeff_9_nxtber_less_int,
		gen3_coeff_9_nxtber_more	=>	gen3_coeff_9_nxtber_more_int,
		gen3_coeff_9_preset_hint	=>	gen3_coeff_9_preset_hint_int,
		gen3_coeff_9_reqber	=>	gen3_coeff_9_reqber_int,
		gen3_coeff_9_sel	=>	gen3_coeff_9_sel,
		gen3_coeff_delay_count	=>	gen3_coeff_delay_count_int,
		gen3_coeff_errchk	=>	gen3_coeff_errchk,
		gen3_dcbal_en	=>	gen3_dcbal_en,
		gen3_diffclock_nfts_count	=>	gen3_diffclock_nfts_count_int,
		gen3_force_local_coeff	=>	gen3_force_local_coeff,
		gen3_full_swing	=>	gen3_full_swing_int,
		gen3_half_swing	=>	gen3_half_swing,
		gen3_low_freq	=>	gen3_low_freq_int,
		gen3_paritychk	=>	gen3_paritychk,
		gen3_pl_framing_err_dis	=>	gen3_pl_framing_err_dis,
		gen3_preset_coeff_1	=>	gen3_preset_coeff_1_int,
		gen3_preset_coeff_10	=>	gen3_preset_coeff_10_int,
		gen3_preset_coeff_11	=>	gen3_preset_coeff_11_int,
		gen3_preset_coeff_2	=>	gen3_preset_coeff_2_int,
		gen3_preset_coeff_3	=>	gen3_preset_coeff_3_int,
		gen3_preset_coeff_4	=>	gen3_preset_coeff_4_int,
		gen3_preset_coeff_5	=>	gen3_preset_coeff_5_int,
		gen3_preset_coeff_6	=>	gen3_preset_coeff_6_int,
		gen3_preset_coeff_7	=>	gen3_preset_coeff_7_int,
		gen3_preset_coeff_8	=>	gen3_preset_coeff_8_int,
		gen3_preset_coeff_9	=>	gen3_preset_coeff_9_int,
		gen3_reset_eieos_cnt_bit	=>	gen3_reset_eieos_cnt_bit,
		gen3_rxfreqlock_counter	=>	gen3_rxfreqlock_counter_int,
		gen3_sameclock_nfts_count	=>	gen3_sameclock_nfts_count_int,
		gen3_scrdscr_bypass	=>	gen3_scrdscr_bypass,
		gen3_skip_ph2_ph3	=>	gen3_skip_ph2_ph3,
		hard_reset_bypass	=>	hard_reset_bypass,
		hard_rst_sig_chnl_en	=>	hard_rst_sig_chnl_en,
		hard_rst_tx_pll_rst_chnl_en	=>	hard_rst_tx_pll_rst_chnl_en,
		hip_ac_pwr_clk_freq_in_hz	=>	hip_ac_pwr_clk_freq_in_hz_int,
		hip_ac_pwr_uw_per_mhz	=>	hip_ac_pwr_uw_per_mhz_int,
		hip_base_address	=>	hip_base_address_int,
		hip_clock_dis	=>	hip_clock_dis,
		hip_hard_reset	=>	hip_hard_reset,
		hip_pcs_sig_chnl_en	=>	hip_pcs_sig_chnl_en,
		hot_plug_support	=>	hot_plug_support_int,
		hrc_chnl_txpll_master_cgb_rst_select	=>	hrc_chnl_txpll_master_cgb_rst_select,
		hrdrstctrl_en	=>	hrdrstctrl_en,
		iei_enable_settings	=>	iei_enable_settings,
		indicator	=>	indicator_int,
		intel_id_access	=>	intel_id_access,
		interrupt_pin	=>	interrupt_pin,
		io_window_addr_width	=>	io_window_addr_width,
		jtag_id	=>	jtag_id,
		ko_compl_data	=>	ko_compl_data_int,
		ko_compl_header	=>	ko_compl_header_int,
		l01_entry_latency	=>	l01_entry_latency_int,
		l0_exit_latency_diffclock	=>	l0_exit_latency_diffclock_int,
		l0_exit_latency_sameclock	=>	l0_exit_latency_sameclock_int,
		l0s_adj_rply_timer_dis	=>	l0s_adj_rply_timer_dis,
		l1_exit_latency_diffclock	=>	l1_exit_latency_diffclock_int,
		l1_exit_latency_sameclock	=>	l1_exit_latency_sameclock_int,
		l2_async_logic	=>	l2_async_logic,
		lane_mask	=>	lane_mask,
		lane_rate	=>	lane_rate,
		link_width	=>	link_width,
		lmi_hold_off_cfg_timer_en	=>	lmi_hold_off_cfg_timer_en,
		low_priority_vc	=>	low_priority_vc,
		ltr_mechanism	=>	ltr_mechanism,
		ltssm_1ms_timeout	=>	ltssm_1ms_timeout,
		ltssm_freqlocked_check	=>	ltssm_freqlocked_check,
		malformed_tlp_truncate_en	=>	malformed_tlp_truncate_en,
		max_link_width	=>	max_link_width,
		max_payload_size	=>	max_payload_size,
		maximum_current	=>	maximum_current_int,
		millisecond_cycle_count	=>	millisecond_cycle_count_int,
		msi_64bit_addressing_capable	=>	msi_64bit_addressing_capable,
		msi_masking_capable	=>	msi_masking_capable,
		msi_multi_message_capable	=>	msi_multi_message_capable,
		msi_support	=>	msi_support,
		msix_pba_bir	=>	msix_pba_bir_int,
		msix_pba_offset	=>	msix_pba_offset_int,
		msix_table_bir	=>	msix_table_bir_int,
		msix_table_offset	=>	msix_table_offset_int,
		msix_table_size	=>	msix_table_size_int,
		national_inst_thru_enhance	=>	national_inst_thru_enhance,
		no_command_completed	=>	no_command_completed,
		no_soft_reset	=>	no_soft_reset,
		not_use_k_gbl_bits	=>	not_use_k_gbl_bits,
		operating_voltage	=>	operating_voltage,
		pcie_base_spec	=>	pcie_base_spec,
		pcie_mode	=>	pcie_mode,
		pcie_spec_1p0_compliance	=>	pcie_spec_1p0_compliance,
		pcie_spec_version	=>	pcie_spec_version,
		pclk_out_sel	=>	pclk_out_sel,
		pld_in_use_reg	=>	pld_in_use_reg,
		pm_latency_patch_dis	=>	pm_latency_patch_dis,
		pm_txdl_patch_dis	=>	pm_txdl_patch_dis,
		pme_clock	=>	pme_clock,
		port_link_number	=>	port_link_number_int,
		port_type	=>	port_type,
		powerdown_mode	=>	powerdown_mode,
		prefetchable_mem_window_addr_width	=>	prefetchable_mem_window_addr_width,
		r2c_mask_easy	=>	r2c_mask_easy,
		r2c_mask_enable	=>	r2c_mask_enable,
		rec_frqlk_mon_en	=>	rec_frqlk_mon_en,
		register_pipe_signals	=>	register_pipe_signals,
		retry_buffer_last_active_address	=>	retry_buffer_last_active_address_int,
		retry_buffer_memory_settings	=>	retry_buffer_memory_settings,
		retry_ecc_corr_mask_dis	=>	retry_ecc_corr_mask_dis,
		revision_id	=>	revision_id_int,
		role_based_error_reporting	=>	role_based_error_reporting,
		rp_bug_fix_pri_sec_stat_reg	=>	rp_bug_fix_pri_sec_stat_reg_int,
		rpltim_base	=>	rpltim_base_int,
		rpltim_set	=>	rpltim_set,
		rstctl_ltssm_dis	=>	rstctl_ltssm_dis,
		rstctrl_1ms_count_fref_clk	=>	rstctrl_1ms_count_fref_clk_int,
		rstctrl_1us_count_fref_clk	=>	rstctrl_1us_count_fref_clk_int,
		rstctrl_altpe3_crst_n_inv	=>	rstctrl_altpe3_crst_n_inv,
		rstctrl_altpe3_rst_n_inv	=>	rstctrl_altpe3_rst_n_inv,
		rstctrl_altpe3_srst_n_inv	=>	rstctrl_altpe3_srst_n_inv,
		rstctrl_chnl_cal_done_select	=>	rstctrl_chnl_cal_done_select,
		rstctrl_debug_en	=>	rstctrl_debug_en,
		rstctrl_force_inactive_rst	=>	rstctrl_force_inactive_rst,
		rstctrl_fref_clk_select	=>	rstctrl_fref_clk_select,
		rstctrl_hard_block_enable	=>	rstctrl_hard_block_enable,
		rstctrl_hip_ep	=>	rstctrl_hip_ep,
		rstctrl_mask_tx_pll_lock_select	=>	rstctrl_mask_tx_pll_lock_select,
		rstctrl_perst_enable	=>	rstctrl_perst_enable,
		rstctrl_perstn_select	=>	rstctrl_perstn_select,
		rstctrl_pld_clr	=>	rstctrl_pld_clr,
		rstctrl_pll_cal_done_select	=>	rstctrl_pll_cal_done_select,
		rstctrl_rx_pcs_rst_n_inv	=>	rstctrl_rx_pcs_rst_n_inv,
		rstctrl_rx_pcs_rst_n_select	=>	rstctrl_rx_pcs_rst_n_select,
		rstctrl_rx_pll_freq_lock_select	=>	rstctrl_rx_pll_freq_lock_select,
		rstctrl_rx_pll_lock_select	=>	rstctrl_rx_pll_lock_select,
		rstctrl_rx_pma_rstb_inv	=>	rstctrl_rx_pma_rstb_inv,
		rstctrl_rx_pma_rstb_select	=>	rstctrl_rx_pma_rstb_select,
		rstctrl_timer_a	=>	rstctrl_timer_a_int,
		rstctrl_timer_a_type	=>	rstctrl_timer_a_type,
		rstctrl_timer_b	=>	rstctrl_timer_b_int,
		rstctrl_timer_b_type	=>	rstctrl_timer_b_type,
		rstctrl_timer_c	=>	rstctrl_timer_c_int,
		rstctrl_timer_c_type	=>	rstctrl_timer_c_type,
		rstctrl_timer_d	=>	rstctrl_timer_d_int,
		rstctrl_timer_d_type	=>	rstctrl_timer_d_type,
		rstctrl_timer_e	=>	rstctrl_timer_e_int,
		rstctrl_timer_e_type	=>	rstctrl_timer_e_type,
		rstctrl_timer_f	=>	rstctrl_timer_f_int,
		rstctrl_timer_f_type	=>	rstctrl_timer_f_type,
		rstctrl_timer_g	=>	rstctrl_timer_g_int,
		rstctrl_timer_g_type	=>	rstctrl_timer_g_type,
		rstctrl_timer_h	=>	rstctrl_timer_h_int,
		rstctrl_timer_h_type	=>	rstctrl_timer_h_type,
		rstctrl_timer_i	=>	rstctrl_timer_i_int,
		rstctrl_timer_i_type	=>	rstctrl_timer_i_type,
		rstctrl_timer_j	=>	rstctrl_timer_j_int,
		rstctrl_timer_j_type	=>	rstctrl_timer_j_type,
		rstctrl_tx_lcff_pll_lock_select	=>	rstctrl_tx_lcff_pll_lock_select,
		rstctrl_tx_lcff_pll_rstb_select	=>	rstctrl_tx_lcff_pll_rstb_select,
		rstctrl_tx_pcs_rst_n_inv	=>	rstctrl_tx_pcs_rst_n_inv,
		rstctrl_tx_pcs_rst_n_select	=>	rstctrl_tx_pcs_rst_n_select,
		rstctrl_tx_pma_rstb_inv	=>	rstctrl_tx_pma_rstb_inv,
		rstctrl_tx_pma_syncp_inv	=>	rstctrl_tx_pma_syncp_inv,
		rstctrl_tx_pma_syncp_select	=>	rstctrl_tx_pma_syncp_select,
		rx_ast_parity	=>	rx_ast_parity,
		rx_buffer_credit_alloc	=>	rx_buffer_credit_alloc,
		rx_buffer_fc_protect	=>	rx_buffer_fc_protect_int,
		rx_buffer_protect	=>	rx_buffer_protect_int,
		rx_cdc_almost_empty	=>	rx_cdc_almost_empty_int,
		rx_cdc_almost_full	=>	rx_cdc_almost_full_int,
		rx_cred_ctl_param	=>	rx_cred_ctl_param,
		rx_ei_l0s	=>	rx_ei_l0s,
		rx_l0s_count_idl	=>	rx_l0s_count_idl_int,
		rx_ptr0_nonposted_dpram_max	=>	rx_ptr0_nonposted_dpram_max_int,
		rx_ptr0_nonposted_dpram_min	=>	rx_ptr0_nonposted_dpram_min_int,
		rx_ptr0_posted_dpram_max	=>	rx_ptr0_posted_dpram_max_int,
		rx_ptr0_posted_dpram_min	=>	rx_ptr0_posted_dpram_min_int,
		rx_runt_patch_dis	=>	rx_runt_patch_dis,
		rx_sop_ctrl	=>	rx_sop_ctrl,
		rx_trunc_patch_dis	=>	rx_trunc_patch_dis,
		rx_use_prst	=>	rx_use_prst,
		rx_use_prst_ep	=>	rx_use_prst_ep,
		rxbuf_ecc_corr_mask_dis	=>	rxbuf_ecc_corr_mask_dis,
		rxdl_bad_sop_eop_filter_dis	=>	rxdl_bad_sop_eop_filter_dis,
		rxdl_bad_tlp_patch_dis	=>	rxdl_bad_tlp_patch_dis,
		rxdl_lcrc_patch_dis	=>	rxdl_lcrc_patch_dis,
		sameclock_nfts_count	=>	sameclock_nfts_count_int,
		sel_enable_pcs_rx_fifo_err	=>	sel_enable_pcs_rx_fifo_err,
		silicon_rev	=>	silicon_rev,
		sim_mode	=>	sim_mode,
		simple_ro_fifo_control_en	=>	simple_ro_fifo_control_en,
		single_rx_detect	=>	single_rx_detect,
		skp_os_gen3_count	=>	skp_os_gen3_count_int,
		skp_os_schedule_count	=>	skp_os_schedule_count_int,
		slot_number	=>	slot_number_int,
		slot_power_limit	=>	slot_power_limit_int,
		slot_power_scale	=>	slot_power_scale_int,
		slotclk_cfg	=>	slotclk_cfg,
		ssid	=>	ssid_int,
		ssvid	=>	ssvid_int,
		subsystem_device_id	=>	subsystem_device_id_int,
		subsystem_vendor_id	=>	subsystem_vendor_id_int,
		sup_mode	=>	sup_mode,
		surprise_down_error_support	=>	surprise_down_error_support,
		tl_cfg_div	=>	tl_cfg_div,
		tl_tx_check_parity_msg	=>	tl_tx_check_parity_msg,
		tph_completer	=>	tph_completer,
		tx_ast_parity	=>	tx_ast_parity,
		tx_cdc_almost_empty	=>	tx_cdc_almost_empty_int,
		tx_cdc_almost_full	=>	tx_cdc_almost_full_int,
		tx_sop_ctrl	=>	tx_sop_ctrl,
		tx_swing	=>	tx_swing_int,
		txdl_fair_arbiter_counter	=>	txdl_fair_arbiter_counter_int,
		txdl_fair_arbiter_en	=>	txdl_fair_arbiter_en,
		txrate_adv	=>	txrate_adv,
		uc_calibration_en	=>	uc_calibration_en,
		use_aer	=>	use_aer,
		use_crc_forwarding	=>	use_crc_forwarding,
		user_id	=>	user_id_int,
		vc0_clk_enable	=>	vc0_clk_enable,
		vc0_rx_buffer_memory_settings	=>	vc0_rx_buffer_memory_settings,
		vc0_rx_flow_ctrl_compl_data	=>	vc0_rx_flow_ctrl_compl_data_int,
		vc0_rx_flow_ctrl_compl_header	=>	vc0_rx_flow_ctrl_compl_header_int,
		vc0_rx_flow_ctrl_nonposted_data	=>	vc0_rx_flow_ctrl_nonposted_data_int,
		vc0_rx_flow_ctrl_nonposted_header	=>	vc0_rx_flow_ctrl_nonposted_header_int,
		vc0_rx_flow_ctrl_posted_data	=>	vc0_rx_flow_ctrl_posted_data_int,
		vc0_rx_flow_ctrl_posted_header	=>	vc0_rx_flow_ctrl_posted_header_int,
		vc1_clk_enable	=>	vc1_clk_enable,
		vc_arbitration	=>	vc_arbitration,
		vc_enable	=>	vc_enable,
		vendor_id	=>	vendor_id_int,
		vsec_cap	=>	vsec_cap_int,
		vsec_id	=>	vsec_id_int,
		wrong_device_id	=>	wrong_device_id
	)
	port map (
		-- Instance ports
		aer_msi_num	=>	aer_msi_num,
		app_int_err	=>	app_int_err,
		app_inta_sts	=>	app_inta_sts,
		app_msi_num	=>	app_msi_num,
		app_msi_req	=>	app_msi_req,
		app_msi_tc	=>	app_msi_tc,
		atpg_los_en_n	=>	atpg_los_en_n,
		avmm_address	=>	avmm_address,
		avmm_byte_en	=>	avmm_byte_en,
		avmm_clk	=>	avmm_clk,
		avmm_read	=>	avmm_read,
		avmm_rst_n	=>	avmm_rst_n,
		avmm_write	=>	avmm_write,
		avmm_writedata	=>	avmm_writedata,
		bist_scanen	=>	bist_scanen,
		bist_scanin	=>	bist_scanin,
		bisten_rcv_n	=>	bisten_rcv_n,
		bisten_rpl_n	=>	bisten_rpl_n,
		bistmode_n	=>	bistmode_n,
		cfg_link2csr_pld	=>	cfg_link2csr_pld,
		cfg_prmbus_pld	=>	cfg_prmbus_pld,
		chnl_cal_done0	=>	chnl_cal_done0,
		chnl_cal_done1	=>	chnl_cal_done1,
		chnl_cal_done2	=>	chnl_cal_done2,
		chnl_cal_done3	=>	chnl_cal_done3,
		chnl_cal_done4	=>	chnl_cal_done4,
		chnl_cal_done5	=>	chnl_cal_done5,
		chnl_cal_done6	=>	chnl_cal_done6,
		chnl_cal_done7	=>	chnl_cal_done7,
		core_clk_in	=>	core_clk_in,
		core_crst	=>	core_crst,
		core_por	=>	core_por,
		core_rst	=>	core_rst,
		core_srst	=>	core_srst,
		cpl_err	=>	cpl_err,
		cpl_pending	=>	cpl_pending,
		cseb_rddata	=>	cseb_rddata,
		cseb_rddata_parity	=>	cseb_rddata_parity,
		cseb_rdresponse	=>	cseb_rdresponse,
		cseb_waitrequest	=>	cseb_waitrequest,
		cseb_wrresp_valid	=>	cseb_wrresp_valid,
		cseb_wrresponse	=>	cseb_wrresponse,
		csr_cbdin	=>	csr_cbdin,
		csr_clk	=>	csr_clk,
		csr_din	=>	csr_din,
		csr_en	=>	csr_en,
		csr_enscan	=>	csr_enscan,
		csr_entest	=>	csr_entest,
		csr_in	=>	csr_in,
		csr_load_csr	=>	csr_load_csr,
		csr_pipe_in	=>	csr_pipe_in,
		csr_seg	=>	csr_seg,
		csr_tcsrin	=>	csr_tcsrin,
		csr_tverify	=>	csr_tverify,
		cvp_config_done	=>	cvp_config_done,
		cvp_config_error	=>	cvp_config_error,
		cvp_config_ready	=>	cvp_config_ready,
		cvp_en	=>	cvp_en,
		egress_blk_err	=>	egress_blk_err,
		entest	=>	entest,
		flr_reset	=>	flr_reset,
		force_tx_eidle	=>	force_tx_eidle,
		fref_clk0	=>	fref_clk0,
		fref_clk1	=>	fref_clk1,
		fref_clk2	=>	fref_clk2,
		fref_clk3	=>	fref_clk3,
		fref_clk4	=>	fref_clk4,
		fref_clk5	=>	fref_clk5,
		fref_clk6	=>	fref_clk6,
		fref_clk7	=>	fref_clk7,
		frzlogic	=>	frzlogic,
		frzreg	=>	frzreg,
		hold_ltssm_rec	=>	hold_ltssm_rec,
		hpg_ctrler	=>	hpg_ctrler,
		iocsrrdy_dly	=>	iocsrrdy_dly,
		lmi_addr	=>	lmi_addr,
		lmi_din	=>	lmi_din,
		lmi_rden	=>	lmi_rden,
		lmi_wren	=>	lmi_wren,
		m10k_select	=>	m10k_select,
		mask_tx_pll_lock0	=>	mask_tx_pll_lock0,
		mask_tx_pll_lock1	=>	mask_tx_pll_lock1,
		mask_tx_pll_lock2	=>	mask_tx_pll_lock2,
		mask_tx_pll_lock3	=>	mask_tx_pll_lock3,
		mask_tx_pll_lock4	=>	mask_tx_pll_lock4,
		mask_tx_pll_lock5	=>	mask_tx_pll_lock5,
		mask_tx_pll_lock6	=>	mask_tx_pll_lock6,
		mask_tx_pll_lock7	=>	mask_tx_pll_lock7,
		mem_hip_test_enable	=>	mem_hip_test_enable,
		mem_regscanen_n	=>	mem_regscanen_n,
		mem_rscin_rcv_bot	=>	mem_rscin_rcv_bot,
		mem_rscin_rcv_top	=>	mem_rscin_rcv_top,
		mem_rscin_rtry	=>	mem_rscin_rtry,
		nfrzdrv	=>	nfrzdrv,
		npor	=>	npor,
		pclk_central	=>	pclk_central,
		pclk_ch0	=>	pclk_ch0,
		pclk_ch1	=>	pclk_ch1,
		pex_msi_num	=>	pex_msi_num,
		phy_rst	=>	phy_rst,
		phy_srst	=>	phy_srst,
		phystatus0	=>	phystatus0,
		phystatus1	=>	phystatus1,
		phystatus2	=>	phystatus2,
		phystatus3	=>	phystatus3,
		phystatus4	=>	phystatus4,
		phystatus5	=>	phystatus5,
		phystatus6	=>	phystatus6,
		phystatus7	=>	phystatus7,
		pin_perst_n	=>	pin_perst_n,
		pld_clk	=>	pld_clk,
		pld_clrhip_n	=>	pld_clrhip_n,
		pld_clrpcship_n	=>	pld_clrpcship_n,
		pld_clrpmapcship_n	=>	pld_clrpmapcship_n,
		pld_core_ready	=>	pld_core_ready,
		pld_gp_status	=>	pld_gp_status,
		pld_perst_n	=>	pld_perst_n,
		pll_cal_done0	=>	pll_cal_done0,
		pll_cal_done1	=>	pll_cal_done1,
		pll_cal_done2	=>	pll_cal_done2,
		pll_cal_done3	=>	pll_cal_done3,
		pll_cal_done4	=>	pll_cal_done4,
		pll_cal_done5	=>	pll_cal_done5,
		pll_cal_done6	=>	pll_cal_done6,
		pll_cal_done7	=>	pll_cal_done7,
		pll_fixed_clk_central	=>	pll_fixed_clk_central,
		pll_fixed_clk_ch0	=>	pll_fixed_clk_ch0,
		pll_fixed_clk_ch1	=>	pll_fixed_clk_ch1,
		plniotri	=>	plniotri,
		pm_auxpwr	=>	pm_auxpwr,
		pm_data	=>	pm_data,
		pm_event	=>	pm_event,
		pm_exit_d0_ack	=>	pm_exit_d0_ack,
		pme_to_cr	=>	pme_to_cr,
		reserved_clk_in	=>	reserved_clk_in,
		reserved_in	=>	reserved_in,
		rx_cred_ctl	=>	rx_cred_ctl,
		rx_pll_freq_lock0	=>	rx_pll_freq_lock0,
		rx_pll_freq_lock1	=>	rx_pll_freq_lock1,
		rx_pll_freq_lock2	=>	rx_pll_freq_lock2,
		rx_pll_freq_lock3	=>	rx_pll_freq_lock3,
		rx_pll_freq_lock4	=>	rx_pll_freq_lock4,
		rx_pll_freq_lock5	=>	rx_pll_freq_lock5,
		rx_pll_freq_lock6	=>	rx_pll_freq_lock6,
		rx_pll_freq_lock7	=>	rx_pll_freq_lock7,
		rx_pll_phase_lock0	=>	rx_pll_phase_lock0,
		rx_pll_phase_lock1	=>	rx_pll_phase_lock1,
		rx_pll_phase_lock2	=>	rx_pll_phase_lock2,
		rx_pll_phase_lock3	=>	rx_pll_phase_lock3,
		rx_pll_phase_lock4	=>	rx_pll_phase_lock4,
		rx_pll_phase_lock5	=>	rx_pll_phase_lock5,
		rx_pll_phase_lock6	=>	rx_pll_phase_lock6,
		rx_pll_phase_lock7	=>	rx_pll_phase_lock7,
		rx_st_mask	=>	rx_st_mask,
		rx_st_ready	=>	rx_st_ready,
		rxblkst0	=>	rxblkst0,
		rxblkst1	=>	rxblkst1,
		rxblkst2	=>	rxblkst2,
		rxblkst3	=>	rxblkst3,
		rxblkst4	=>	rxblkst4,
		rxblkst5	=>	rxblkst5,
		rxblkst6	=>	rxblkst6,
		rxblkst7	=>	rxblkst7,
		rxdata0	=>	rxdata0,
		rxdata1	=>	rxdata1,
		rxdata2	=>	rxdata2,
		rxdata3	=>	rxdata3,
		rxdata4	=>	rxdata4,
		rxdata5	=>	rxdata5,
		rxdata6	=>	rxdata6,
		rxdata7	=>	rxdata7,
		rxdatak0	=>	rxdatak0,
		rxdatak1	=>	rxdatak1,
		rxdatak2	=>	rxdatak2,
		rxdatak3	=>	rxdatak3,
		rxdatak4	=>	rxdatak4,
		rxdatak5	=>	rxdatak5,
		rxdatak6	=>	rxdatak6,
		rxdatak7	=>	rxdatak7,
		rxdataskip0	=>	rxdataskip0,
		rxdataskip1	=>	rxdataskip1,
		rxdataskip2	=>	rxdataskip2,
		rxdataskip3	=>	rxdataskip3,
		rxdataskip4	=>	rxdataskip4,
		rxdataskip5	=>	rxdataskip5,
		rxdataskip6	=>	rxdataskip6,
		rxdataskip7	=>	rxdataskip7,
		rxelecidle0	=>	rxelecidle0,
		rxelecidle1	=>	rxelecidle1,
		rxelecidle2	=>	rxelecidle2,
		rxelecidle3	=>	rxelecidle3,
		rxelecidle4	=>	rxelecidle4,
		rxelecidle5	=>	rxelecidle5,
		rxelecidle6	=>	rxelecidle6,
		rxelecidle7	=>	rxelecidle7,
		rxfreqlocked0	=>	rxfreqlocked0,
		rxfreqlocked1	=>	rxfreqlocked1,
		rxfreqlocked2	=>	rxfreqlocked2,
		rxfreqlocked3	=>	rxfreqlocked3,
		rxfreqlocked4	=>	rxfreqlocked4,
		rxfreqlocked5	=>	rxfreqlocked5,
		rxfreqlocked6	=>	rxfreqlocked6,
		rxfreqlocked7	=>	rxfreqlocked7,
		rxstatus0	=>	rxstatus0,
		rxstatus1	=>	rxstatus1,
		rxstatus2	=>	rxstatus2,
		rxstatus3	=>	rxstatus3,
		rxstatus4	=>	rxstatus4,
		rxstatus5	=>	rxstatus5,
		rxstatus6	=>	rxstatus6,
		rxstatus7	=>	rxstatus7,
		rxsynchd0	=>	rxsynchd0,
		rxsynchd1	=>	rxsynchd1,
		rxsynchd2	=>	rxsynchd2,
		rxsynchd3	=>	rxsynchd3,
		rxsynchd4	=>	rxsynchd4,
		rxsynchd5	=>	rxsynchd5,
		rxsynchd6	=>	rxsynchd6,
		rxsynchd7	=>	rxsynchd7,
		rxvalid0	=>	rxvalid0,
		rxvalid1	=>	rxvalid1,
		rxvalid2	=>	rxvalid2,
		rxvalid3	=>	rxvalid3,
		rxvalid4	=>	rxvalid4,
		rxvalid5	=>	rxvalid5,
		rxvalid6	=>	rxvalid6,
		rxvalid7	=>	rxvalid7,
		scan_mode_n	=>	scan_mode_n,
		scan_shift_n	=>	scan_shift_n,
		sw_ctmod	=>	sw_ctmod,
		swdn_in	=>	swdn_in,
		swup_in	=>	swup_in,
		test_in_1_hip	=>	test_in_1_hip,
		test_in_hip	=>	test_in_hip,
		test_pl_dbg_eqin	=>	test_pl_dbg_eqin,
		tx_cred_cons_select	=>	tx_cred_cons_select,
		tx_cred_fc_sel	=>	tx_cred_fc_sel,
		tx_lcff_pll_lock0	=>	tx_lcff_pll_lock0,
		tx_lcff_pll_lock1	=>	tx_lcff_pll_lock1,
		tx_lcff_pll_lock2	=>	tx_lcff_pll_lock2,
		tx_lcff_pll_lock3	=>	tx_lcff_pll_lock3,
		tx_lcff_pll_lock4	=>	tx_lcff_pll_lock4,
		tx_lcff_pll_lock5	=>	tx_lcff_pll_lock5,
		tx_lcff_pll_lock6	=>	tx_lcff_pll_lock6,
		tx_lcff_pll_lock7	=>	tx_lcff_pll_lock7,
		tx_st_data	=>	tx_st_data,
		tx_st_empty	=>	tx_st_empty,
		tx_st_eop	=>	tx_st_eop,
		tx_st_err	=>	tx_st_err,
		tx_st_parity	=>	tx_st_parity,
		tx_st_sop	=>	tx_st_sop,
		tx_st_valid	=>	tx_st_valid,
		user_mode	=>	user_mode,
		sta_hd_altpe3_hip_core_top_hd_altpe3_hip_core_u_clkmux_core_clk_cnt_reg_0_0_Q	=>	sta_hd_altpe3_hip_core_top_hd_altpe3_hip_core_u_clkmux_core_clk_cnt_reg_0_0_Q,
		sta_hd_altpe3_hip_core_top_hd_altpe3_hip_core_u_clkmux_core_clk_cnt_reg_1_0_Q	=>	sta_hd_altpe3_hip_core_top_hd_altpe3_hip_core_u_clkmux_core_clk_cnt_reg_1_0_Q,
		sta_hd_altpe3_hip_core_top_hd_altpe3_hip_core_u_clkmux_core_clk_cnt_reg_2_0_Q	=>	sta_hd_altpe3_hip_core_top_hd_altpe3_hip_core_u_clkmux_core_clk_cnt_reg_2_0_Q,
		app_inta_ack	=>	app_inta_ack,
		app_msi_ack	=>	app_msi_ack,
		avmm_readdata	=>	avmm_readdata,
		cfg_par_err	=>	cfg_par_err,
		core_clk_out	=>	core_clk_out,
		cseb_addr	=>	cseb_addr,
		cseb_addr_parity	=>	cseb_addr_parity,
		cseb_be	=>	cseb_be,
		cseb_is_shadow	=>	cseb_is_shadow,
		cseb_rden	=>	cseb_rden,
		cseb_wrdata	=>	cseb_wrdata,
		cseb_wrdata_parity	=>	cseb_wrdata_parity,
		cseb_wren	=>	cseb_wren,
		cseb_wrresp_req	=>	cseb_wrresp_req,
		csr_dout	=>	csr_dout,
		csr_out	=>	csr_out,
		csr_pipe_out	=>	csr_pipe_out,
		current_coeff0	=>	current_coeff0,
		current_coeff1	=>	current_coeff1,
		current_coeff2	=>	current_coeff2,
		current_coeff3	=>	current_coeff3,
		current_coeff4	=>	current_coeff4,
		current_coeff5	=>	current_coeff5,
		current_coeff6	=>	current_coeff6,
		current_coeff7	=>	current_coeff7,
		current_rxpreset0	=>	current_rxpreset0,
		current_rxpreset1	=>	current_rxpreset1,
		current_rxpreset2	=>	current_rxpreset2,
		current_rxpreset3	=>	current_rxpreset3,
		current_rxpreset4	=>	current_rxpreset4,
		current_rxpreset5	=>	current_rxpreset5,
		current_rxpreset6	=>	current_rxpreset6,
		current_rxpreset7	=>	current_rxpreset7,
		current_speed	=>	current_speed,
		cvp_clk	=>	cvp_clk,
		cvp_config	=>	cvp_config,
		cvp_data	=>	cvp_data,
		cvp_full_config	=>	cvp_full_config,
		cvp_start_xfer	=>	cvp_start_xfer,
		dl_up	=>	dl_up,
		dlup_exit	=>	dlup_exit,
		eidle_infer_sel0	=>	eidle_infer_sel0,
		eidle_infer_sel1	=>	eidle_infer_sel1,
		eidle_infer_sel2	=>	eidle_infer_sel2,
		eidle_infer_sel3	=>	eidle_infer_sel3,
		eidle_infer_sel4	=>	eidle_infer_sel4,
		eidle_infer_sel5	=>	eidle_infer_sel5,
		eidle_infer_sel6	=>	eidle_infer_sel6,
		eidle_infer_sel7	=>	eidle_infer_sel7,
		ev_128ns	=>	ev_128ns,
		ev_1us	=>	ev_1us,
		flr_sts	=>	flr_sts,
		g3_rx_pcs_rst_n0	=>	g3_rx_pcs_rst_n0,
		g3_rx_pcs_rst_n1	=>	g3_rx_pcs_rst_n1,
		g3_rx_pcs_rst_n2	=>	g3_rx_pcs_rst_n2,
		g3_rx_pcs_rst_n3	=>	g3_rx_pcs_rst_n3,
		g3_rx_pcs_rst_n4	=>	g3_rx_pcs_rst_n4,
		g3_rx_pcs_rst_n5	=>	g3_rx_pcs_rst_n5,
		g3_rx_pcs_rst_n6	=>	g3_rx_pcs_rst_n6,
		g3_rx_pcs_rst_n7	=>	g3_rx_pcs_rst_n7,
		g3_tx_pcs_rst_n0	=>	g3_tx_pcs_rst_n0,
		g3_tx_pcs_rst_n1	=>	g3_tx_pcs_rst_n1,
		g3_tx_pcs_rst_n2	=>	g3_tx_pcs_rst_n2,
		g3_tx_pcs_rst_n3	=>	g3_tx_pcs_rst_n3,
		g3_tx_pcs_rst_n4	=>	g3_tx_pcs_rst_n4,
		g3_tx_pcs_rst_n5	=>	g3_tx_pcs_rst_n5,
		g3_tx_pcs_rst_n6	=>	g3_tx_pcs_rst_n6,
		g3_tx_pcs_rst_n7	=>	g3_tx_pcs_rst_n7,
		hotrst_exit	=>	hotrst_exit,
		int_status	=>	int_status,
		k_hip_pcs_chnl_en	=>	k_hip_pcs_chnl_en,
		k_hrc_chnl_en	=>	k_hrc_chnl_en,
		k_hrc_chnl_txpll_master_cgb_rst_en	=>	k_hrc_chnl_txpll_master_cgb_rst_en,
		k_hrc_chnl_txpll_rst_en	=>	k_hrc_chnl_txpll_rst_en,
		l2_exit	=>	l2_exit,
		lane_act	=>	lane_act,
		lmi_ack	=>	lmi_ack,
		lmi_dout	=>	lmi_dout,
		ltssm_state	=>	ltssm_state,
		mem_rscout_rcv_bot	=>	mem_rscout_rcv_bot,
		mem_rscout_rcv_top	=>	mem_rscout_rcv_top,
		mem_rscout_rtry	=>	mem_rscout_rtry,
		pld_clk_in_use	=>	pld_clk_in_use,
		pld_gp_ctrl	=>	pld_gp_ctrl,
		pm_exit_d0_req	=>	pm_exit_d0_req,
		pme_to_sr	=>	pme_to_sr,
		powerdown0	=>	powerdown0,
		powerdown1	=>	powerdown1,
		powerdown2	=>	powerdown2,
		powerdown3	=>	powerdown3,
		powerdown4	=>	powerdown4,
		powerdown5	=>	powerdown5,
		powerdown6	=>	powerdown6,
		powerdown7	=>	powerdown7,
		r2c_unc_ecc	=>	r2c_unc_ecc,
		rate0	=>	rate0,
		rate1	=>	rate1,
		rate2	=>	rate2,
		rate3	=>	rate3,
		rate4	=>	rate4,
		rate5	=>	rate5,
		rate6	=>	rate6,
		rate7	=>	rate7,
		rate_ctrl	=>	rate_ctrl,
		reserved_clk_out	=>	reserved_clk_out,
		reserved_out	=>	reserved_out,
		reset_status	=>	reset_status,
		retry_corr_ecc	=>	retry_corr_ecc,
		retry_unc_ecc	=>	retry_unc_ecc,
		rx_corr_ecc	=>	rx_corr_ecc,
		rx_cred_status	=>	rx_cred_status,
		rx_par_err	=>	rx_par_err,
		rx_pcs_rst_n0	=>	rx_pcs_rst_n0,
		rx_pcs_rst_n1	=>	rx_pcs_rst_n1,
		rx_pcs_rst_n2	=>	rx_pcs_rst_n2,
		rx_pcs_rst_n3	=>	rx_pcs_rst_n3,
		rx_pcs_rst_n4	=>	rx_pcs_rst_n4,
		rx_pcs_rst_n5	=>	rx_pcs_rst_n5,
		rx_pcs_rst_n6	=>	rx_pcs_rst_n6,
		rx_pcs_rst_n7	=>	rx_pcs_rst_n7,
		rx_pma_rstb0	=>	rx_pma_rstb0,
		rx_pma_rstb1	=>	rx_pma_rstb1,
		rx_pma_rstb2	=>	rx_pma_rstb2,
		rx_pma_rstb3	=>	rx_pma_rstb3,
		rx_pma_rstb4	=>	rx_pma_rstb4,
		rx_pma_rstb5	=>	rx_pma_rstb5,
		rx_pma_rstb6	=>	rx_pma_rstb6,
		rx_pma_rstb7	=>	rx_pma_rstb7,
		rx_st_bardec1	=>	rx_st_bardec1,
		rx_st_bardec2	=>	rx_st_bardec2,
		rx_st_be	=>	rx_st_be,
		rx_st_data	=>	rx_st_data,
		rx_st_empty	=>	rx_st_empty,
		rx_st_eop	=>	rx_st_eop,
		rx_st_err	=>	rx_st_err,
		rx_st_parity	=>	rx_st_parity,
		rx_st_sop	=>	rx_st_sop,
		rx_st_valid	=>	rx_st_valid,
		rxfc_cplbuf_ovf	=>	rxfc_cplbuf_ovf,
		rxfc_cplovf_tag	=>	rxfc_cplovf_tag,
		rxpolarity0	=>	rxpolarity0,
		rxpolarity1	=>	rxpolarity1,
		rxpolarity2	=>	rxpolarity2,
		rxpolarity3	=>	rxpolarity3,
		rxpolarity4	=>	rxpolarity4,
		rxpolarity5	=>	rxpolarity5,
		rxpolarity6	=>	rxpolarity6,
		rxpolarity7	=>	rxpolarity7,
		serr_out	=>	serr_out,
		swdn_out	=>	swdn_out,
		swup_out	=>	swup_out,
		test_fref_clk	=>	test_fref_clk,
		test_out_1_hip	=>	test_out_1_hip,
		test_out_hip	=>	test_out_hip,
		tl_cfg_add	=>	tl_cfg_add,
		tl_cfg_ctl	=>	tl_cfg_ctl,
		tl_cfg_sts	=>	tl_cfg_sts,
		tl_cfg_sts_wr	=>	tl_cfg_sts_wr,
		tx_cred_data_fc	=>	tx_cred_data_fc,
		tx_cred_fc_hip_cons	=>	tx_cred_fc_hip_cons,
		tx_cred_fc_infinite	=>	tx_cred_fc_infinite,
		tx_cred_hdr_fc	=>	tx_cred_hdr_fc,
		tx_deemph0	=>	tx_deemph0,
		tx_deemph1	=>	tx_deemph1,
		tx_deemph2	=>	tx_deemph2,
		tx_deemph3	=>	tx_deemph3,
		tx_deemph4	=>	tx_deemph4,
		tx_deemph5	=>	tx_deemph5,
		tx_deemph6	=>	tx_deemph6,
		tx_deemph7	=>	tx_deemph7,
		tx_lcff_pll_rstb0	=>	tx_lcff_pll_rstb0,
		tx_lcff_pll_rstb1	=>	tx_lcff_pll_rstb1,
		tx_lcff_pll_rstb2	=>	tx_lcff_pll_rstb2,
		tx_lcff_pll_rstb3	=>	tx_lcff_pll_rstb3,
		tx_lcff_pll_rstb4	=>	tx_lcff_pll_rstb4,
		tx_lcff_pll_rstb5	=>	tx_lcff_pll_rstb5,
		tx_lcff_pll_rstb6	=>	tx_lcff_pll_rstb6,
		tx_lcff_pll_rstb7	=>	tx_lcff_pll_rstb7,
		tx_margin0	=>	tx_margin0,
		tx_margin1	=>	tx_margin1,
		tx_margin2	=>	tx_margin2,
		tx_margin3	=>	tx_margin3,
		tx_margin4	=>	tx_margin4,
		tx_margin5	=>	tx_margin5,
		tx_margin6	=>	tx_margin6,
		tx_margin7	=>	tx_margin7,
		tx_par_err	=>	tx_par_err,
		tx_pcs_rst_n0	=>	tx_pcs_rst_n0,
		tx_pcs_rst_n1	=>	tx_pcs_rst_n1,
		tx_pcs_rst_n2	=>	tx_pcs_rst_n2,
		tx_pcs_rst_n3	=>	tx_pcs_rst_n3,
		tx_pcs_rst_n4	=>	tx_pcs_rst_n4,
		tx_pcs_rst_n5	=>	tx_pcs_rst_n5,
		tx_pcs_rst_n6	=>	tx_pcs_rst_n6,
		tx_pcs_rst_n7	=>	tx_pcs_rst_n7,
		tx_pma_syncp0	=>	tx_pma_syncp0,
		tx_pma_syncp1	=>	tx_pma_syncp1,
		tx_pma_syncp2	=>	tx_pma_syncp2,
		tx_pma_syncp3	=>	tx_pma_syncp3,
		tx_pma_syncp4	=>	tx_pma_syncp4,
		tx_pma_syncp5	=>	tx_pma_syncp5,
		tx_pma_syncp6	=>	tx_pma_syncp6,
		tx_pma_syncp7	=>	tx_pma_syncp7,
		tx_st_ready	=>	tx_st_ready,
		txblkst0	=>	txblkst0,
		txblkst1	=>	txblkst1,
		txblkst2	=>	txblkst2,
		txblkst3	=>	txblkst3,
		txblkst4	=>	txblkst4,
		txblkst5	=>	txblkst5,
		txblkst6	=>	txblkst6,
		txblkst7	=>	txblkst7,
		txcompl0	=>	txcompl0,
		txcompl1	=>	txcompl1,
		txcompl2	=>	txcompl2,
		txcompl3	=>	txcompl3,
		txcompl4	=>	txcompl4,
		txcompl5	=>	txcompl5,
		txcompl6	=>	txcompl6,
		txcompl7	=>	txcompl7,
		txdata0	=>	txdata0,
		txdata1	=>	txdata1,
		txdata2	=>	txdata2,
		txdata3	=>	txdata3,
		txdata4	=>	txdata4,
		txdata5	=>	txdata5,
		txdata6	=>	txdata6,
		txdata7	=>	txdata7,
		txdatak0	=>	txdatak0,
		txdatak1	=>	txdatak1,
		txdatak2	=>	txdatak2,
		txdatak3	=>	txdatak3,
		txdatak4	=>	txdatak4,
		txdatak5	=>	txdatak5,
		txdatak6	=>	txdatak6,
		txdatak7	=>	txdatak7,
		txdataskip0	=>	txdataskip0,
		txdataskip1	=>	txdataskip1,
		txdataskip2	=>	txdataskip2,
		txdataskip3	=>	txdataskip3,
		txdataskip4	=>	txdataskip4,
		txdataskip5	=>	txdataskip5,
		txdataskip6	=>	txdataskip6,
		txdataskip7	=>	txdataskip7,
		txdetectrx0	=>	txdetectrx0,
		txdetectrx1	=>	txdetectrx1,
		txdetectrx2	=>	txdetectrx2,
		txdetectrx3	=>	txdetectrx3,
		txdetectrx4	=>	txdetectrx4,
		txdetectrx5	=>	txdetectrx5,
		txdetectrx6	=>	txdetectrx6,
		txdetectrx7	=>	txdetectrx7,
		txelecidle0	=>	txelecidle0,
		txelecidle1	=>	txelecidle1,
		txelecidle2	=>	txelecidle2,
		txelecidle3	=>	txelecidle3,
		txelecidle4	=>	txelecidle4,
		txelecidle5	=>	txelecidle5,
		txelecidle6	=>	txelecidle6,
		txelecidle7	=>	txelecidle7,
		txst_prot_err	=>	txst_prot_err,
		txswing0	=>	txswing0,
		txswing1	=>	txswing1,
		txswing2	=>	txswing2,
		txswing3	=>	txswing3,
		txswing4	=>	txswing4,
		txswing5	=>	txswing5,
		txswing6	=>	txswing6,
		txswing7	=>	txswing7,
		txsynchd0	=>	txsynchd0,
		txsynchd1	=>	txsynchd1,
		txsynchd2	=>	txsynchd2,
		txsynchd3	=>	txsynchd3,
		txsynchd4	=>	txsynchd4,
		txsynchd5	=>	txsynchd5,
		txsynchd6	=>	txsynchd6,
		txsynchd7	=>	txsynchd7,
		wake_oen	=>	wake_oen
	);

end behavior;
